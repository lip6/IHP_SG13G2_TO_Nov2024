* Extracted by KLayout with SG13G2 LVS runset on : 12/11/2024 03:13

.SUBCKT AC3E_USM_TDBUCK 25|VSS 8 9 10 11 12 13|A|VINR 14|A|VINS 7 15 6 16 5
+ 17|VCN|Y 19|VDD A|Y A|Y$1 A|X A|X$1 A|X$2 A|X$3 A|Y$2 A|B|Y A|X$4 A|X$5
+ A|B|Y$1 A|X$6 A|Y$3 B|X A|Y$4 A|X$7 A|X$8 A|X$9 A|X$10 A|Y$5 A|X$11 X A|Y$6 4
+ A|X$12 A|B|Y$2 A|Y$7 A|B|Y$3 A|X$13 A|X$14 A|X$15 A|X$16 A|Y$8 A|Y$9 A|Y$10
+ A|X$17 A|X$18 A|B|Y$4 A|B|X A|Y$11 A|X$19 A|Y$12 A|Y$13 A|Y$14 22 27 28
+ 18|VCP|Y 23 20 21 3 26 2 1 24
M$1 25|VSS A|Y 17|VCN|Y 25|VSS sg13_lv_nmos L=0.13u W=2.96u AS=0.6734p
+ AD=0.6734p PS=5.52u PD=5.52u
M$5 \$149 A|Y$2 25|VSS 25|VSS sg13_lv_nmos L=0.13u W=0.42u AS=0.1428p
+ AD=0.0798p PS=1.52u PD=0.8u
M$6 25|VSS \$149 \$150 25|VSS sg13_lv_nmos L=0.5u W=0.42u AS=0.0798p AD=0.1428p
+ PS=0.8u PD=1.52u
M$7 25|VSS \$150 \$151 25|VSS sg13_lv_nmos L=0.5u W=0.42u AS=0.1426p AD=0.1428p
+ PS=1.16u PD=1.52u
M$8 25|VSS \$151 A|X 25|VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.1426p AD=0.2516p
+ PS=1.16u PD=2.16u
M$9 \$153 A|X$1 25|VSS 25|VSS sg13_lv_nmos L=0.13u W=0.42u AS=0.1428p
+ AD=0.0798p PS=1.52u PD=0.8u
M$10 25|VSS \$153 \$155 25|VSS sg13_lv_nmos L=0.5u W=0.42u AS=0.0798p
+ AD=0.1428p PS=0.8u PD=1.52u
M$11 25|VSS 14|A|VINS A|Y$1 25|VSS sg13_lv_nmos L=0.13u W=1.48u AS=0.3922p
+ AD=0.3959p PS=3.28u PD=3.29u
M$13 25|VSS \$155 \$156 25|VSS sg13_lv_nmos L=0.5u W=0.42u AS=0.1426p
+ AD=0.1428p PS=1.16u PD=1.52u
M$14 25|VSS \$156 A|X$2 25|VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.1426p
+ AD=0.2516p PS=1.16u PD=2.16u
M$15 25|VSS A|Y$1 A|B|Y 25|VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.259p AD=0.259p
+ PS=2.18u PD=2.18u
M$16 25|VSS A|X$3 A|Y 25|VSS sg13_lv_nmos L=0.13u W=1.48u AS=0.3922p AD=0.3959p
+ PS=3.28u PD=3.29u
M$18 25|VSS A|B|Y A|Y$2 25|VSS sg13_lv_nmos L=0.13u W=5.92u AS=1.2395p
+ AD=1.2395p PS=10.01u PD=10.01u
M$26 \$164 \$163 25|VSS 25|VSS sg13_lv_nmos L=0.5u W=0.42u AS=0.1428p
+ AD=0.1426p PS=1.52u PD=1.16u
M$27 25|VSS \$164 A|X$1 25|VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.1426p
+ AD=0.2516p PS=1.16u PD=2.16u
M$28 25|VSS A|X$5 A|B|Y$1 25|VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.259p
+ AD=0.259p PS=2.18u PD=2.18u
M$29 \$167 A|X$7 25|VSS 25|VSS sg13_lv_nmos L=0.13u W=0.42u AS=0.1428p
+ AD=0.0798p PS=1.52u PD=0.8u
M$30 25|VSS \$167 \$168 25|VSS sg13_lv_nmos L=0.5u W=0.42u AS=0.0798p
+ AD=0.1428p PS=0.8u PD=1.52u
M$31 25|VSS \$168 \$180 25|VSS sg13_lv_nmos L=0.5u W=0.42u AS=0.1426p
+ AD=0.1428p PS=1.16u PD=1.52u
M$32 25|VSS \$180 A|X$6 25|VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.1426p
+ AD=0.2516p PS=1.16u PD=2.16u
M$33 \$170 A|X$8 25|VSS 25|VSS sg13_lv_nmos L=0.13u W=0.42u AS=0.1428p
+ AD=0.0798p PS=1.52u PD=0.8u
M$34 25|VSS \$170 \$171 25|VSS sg13_lv_nmos L=0.5u W=0.42u AS=0.0798p
+ AD=0.1428p PS=0.8u PD=1.52u
M$35 25|VSS \$171 \$182 25|VSS sg13_lv_nmos L=0.5u W=0.42u AS=0.1426p
+ AD=0.1428p PS=1.16u PD=1.52u
M$36 25|VSS \$182 A|X$3 25|VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.1426p
+ AD=0.2516p PS=1.16u PD=2.16u
M$37 \$174 A|X 25|VSS 25|VSS sg13_lv_nmos L=0.13u W=0.42u AS=0.1428p AD=0.0798p
+ PS=1.52u PD=0.8u
M$38 25|VSS \$174 \$175 25|VSS sg13_lv_nmos L=0.5u W=0.42u AS=0.0798p
+ AD=0.1428p PS=0.8u PD=1.52u
M$39 25|VSS \$175 \$184 25|VSS sg13_lv_nmos L=0.5u W=0.42u AS=0.1426p
+ AD=0.1428p PS=1.16u PD=1.52u
M$40 25|VSS \$184 A|X$4 25|VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.1426p
+ AD=0.2516p PS=1.16u PD=2.16u
M$41 \$161 A|X$4 25|VSS 25|VSS sg13_lv_nmos L=0.13u W=0.42u AS=0.1428p
+ AD=0.0798p PS=1.52u PD=0.8u
M$42 25|VSS \$161 \$163 25|VSS sg13_lv_nmos L=0.5u W=0.42u AS=0.0798p
+ AD=0.1428p PS=0.8u PD=1.52u
M$43 \$176 A|X$2 25|VSS 25|VSS sg13_lv_nmos L=0.13u W=0.42u AS=0.1428p
+ AD=0.0798p PS=1.52u PD=0.8u
M$44 25|VSS \$176 \$177 25|VSS sg13_lv_nmos L=0.5u W=0.42u AS=0.0798p
+ AD=0.1428p PS=0.8u PD=1.52u
M$45 25|VSS \$177 \$185 25|VSS sg13_lv_nmos L=0.5u W=0.42u AS=0.1426p
+ AD=0.1428p PS=1.16u PD=1.52u
M$46 25|VSS \$185 A|X$5 25|VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.1426p
+ AD=0.2516p PS=1.16u PD=2.16u
M$47 25|VSS A|B|Y$1 A|Y$3 25|VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.259p
+ AD=0.259p PS=2.18u PD=2.18u
M$48 25|VSS A|B|Y A|Y$4 25|VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.259p AD=0.259p
+ PS=2.18u PD=2.18u
M$49 \$205 \$191 25|VSS 25|VSS sg13_lv_nmos L=0.5u W=0.42u AS=0.1428p
+ AD=0.1426p PS=1.52u PD=1.16u
M$50 25|VSS \$205 A|X$9 25|VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.1426p
+ AD=0.2516p PS=1.16u PD=2.16u
M$51 \$207 \$194 25|VSS 25|VSS sg13_lv_nmos L=0.5u W=0.42u AS=0.1428p
+ AD=0.1426p PS=1.52u PD=1.16u
M$52 25|VSS \$207 A|X$10 25|VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.1426p
+ AD=0.2516p PS=1.16u PD=2.16u
M$53 \$208 \$197 25|VSS 25|VSS sg13_lv_nmos L=0.5u W=0.42u AS=0.1428p
+ AD=0.1426p PS=1.52u PD=1.16u
M$54 25|VSS \$208 A|X$8 25|VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.1426p
+ AD=0.2516p PS=1.16u PD=2.16u
M$55 25|VSS A|X$3 A|Y$5 25|VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.2516p
+ AD=0.1406p PS=2.16u PD=1.12u
M$56 A|Y$5 A|B|Y$2 25|VSS 25|VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.1406p
+ AD=0.2516p PS=1.12u PD=2.16u
M$57 \$183 A|Y$3 \$188 25|VSS sg13_lv_nmos L=0.13u W=0.64u AS=0.2176p
+ AD=0.1216p PS=1.96u PD=1.02u
M$58 25|VSS A|B|Y \$188 25|VSS sg13_lv_nmos L=0.13u W=0.64u AS=0.1331p
+ AD=0.1216p PS=1.12u PD=1.02u
M$59 25|VSS \$183 B|X 25|VSS sg13_lv_nmos L=0.13u W=1.48u AS=0.2737p AD=0.4218p
+ PS=2.24u PD=3.36u
M$61 25|VSS A|Y$7 A|B|Y$2 25|VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.2516p
+ AD=0.1406p PS=2.16u PD=1.12u
M$62 A|B|Y$2 B|X 25|VSS 25|VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.1406p
+ AD=0.2516p PS=1.12u PD=2.16u
M$63 \$199 A|Y$6 \$215 25|VSS sg13_lv_nmos L=0.13u W=0.64u AS=0.2176p
+ AD=0.1216p PS=1.96u PD=1.02u
M$64 \$215 A|B|Y$4 25|VSS 25|VSS sg13_lv_nmos L=0.13u W=0.64u AS=0.1216p
+ AD=0.1331p PS=1.02u PD=1.12u
M$65 25|VSS \$199 A|X$11 25|VSS sg13_lv_nmos L=0.13u W=1.48u AS=0.2737p
+ AD=0.4218p PS=2.24u PD=3.36u
M$67 \$201 A|Y$4 \$214 25|VSS sg13_lv_nmos L=0.13u W=0.64u AS=0.2176p
+ AD=0.1216p PS=1.96u PD=1.02u
M$68 \$214 A|B|Y$1 25|VSS 25|VSS sg13_lv_nmos L=0.13u W=0.64u AS=0.1216p
+ AD=0.1331p PS=1.02u PD=1.12u
M$69 25|VSS \$201 X 25|VSS sg13_lv_nmos L=0.13u W=1.48u AS=0.2737p AD=0.4218p
+ PS=2.24u PD=3.36u
M$71 25|VSS A|B|Y$3 A|Y$6 25|VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.259p
+ AD=0.259p PS=2.18u PD=2.18u
M$72 \$190 A|Y$5 25|VSS 25|VSS sg13_lv_nmos L=0.13u W=0.42u AS=0.1428p
+ AD=0.0798p PS=1.52u PD=0.8u
M$73 25|VSS \$190 \$191 25|VSS sg13_lv_nmos L=0.5u W=0.42u AS=0.0798p
+ AD=0.1428p PS=0.8u PD=1.52u
M$74 \$221 A|X$9 25|VSS 25|VSS sg13_lv_nmos L=0.13u W=0.42u AS=0.1428p
+ AD=0.0798p PS=1.52u PD=0.8u
M$75 25|VSS \$221 \$222 25|VSS sg13_lv_nmos L=0.5u W=0.42u AS=0.0798p
+ AD=0.1428p PS=0.8u PD=1.52u
M$76 25|VSS \$222 \$223 25|VSS sg13_lv_nmos L=0.5u W=0.42u AS=0.1426p
+ AD=0.1428p PS=1.16u PD=1.52u
M$77 25|VSS \$223 A|X$12 25|VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.1426p
+ AD=0.2516p PS=1.16u PD=2.16u
M$78 \$193 A|X$12 25|VSS 25|VSS sg13_lv_nmos L=0.13u W=0.42u AS=0.1428p
+ AD=0.0798p PS=1.52u PD=0.8u
M$79 25|VSS \$193 \$194 25|VSS sg13_lv_nmos L=0.5u W=0.42u AS=0.0798p
+ AD=0.1428p PS=0.8u PD=1.52u
M$80 \$224 A|X$10 25|VSS 25|VSS sg13_lv_nmos L=0.13u W=0.42u AS=0.1428p
+ AD=0.0798p PS=1.52u PD=0.8u
M$81 25|VSS \$224 \$225 25|VSS sg13_lv_nmos L=0.5u W=0.42u AS=0.0798p
+ AD=0.1428p PS=0.8u PD=1.52u
M$82 25|VSS \$225 \$226 25|VSS sg13_lv_nmos L=0.5u W=0.42u AS=0.1426p
+ AD=0.1428p PS=1.16u PD=1.52u
M$83 25|VSS \$226 A|X$13 25|VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.1426p
+ AD=0.2516p PS=1.16u PD=2.16u
M$84 \$196 A|X$6 25|VSS 25|VSS sg13_lv_nmos L=0.13u W=0.42u AS=0.1428p
+ AD=0.0798p PS=1.52u PD=0.8u
M$85 25|VSS \$196 \$197 25|VSS sg13_lv_nmos L=0.5u W=0.42u AS=0.0798p
+ AD=0.1428p PS=0.8u PD=1.52u
M$86 \$227 A|Y$9 25|VSS 25|VSS sg13_lv_nmos L=0.13u W=0.42u AS=0.1428p
+ AD=0.0798p PS=1.52u PD=0.8u
M$87 25|VSS \$227 \$229 25|VSS sg13_lv_nmos L=0.5u W=0.42u AS=0.0798p
+ AD=0.1428p PS=0.8u PD=1.52u
M$88 25|VSS \$229 \$230 25|VSS sg13_lv_nmos L=0.5u W=0.42u AS=0.1426p
+ AD=0.1428p PS=1.16u PD=1.52u
M$89 25|VSS \$230 A|X$14 25|VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.1426p
+ AD=0.2516p PS=1.16u PD=2.16u
M$90 25|VSS A|B|Y$2 A|Y$10 25|VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.259p
+ AD=0.259p PS=2.18u PD=2.18u
M$91 25|VSS A|X$11 A|Y$7 25|VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.2516p
+ AD=0.1406p PS=2.16u PD=1.12u
M$92 A|Y$7 A|B|Y$2 25|VSS 25|VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.1406p
+ AD=0.2516p PS=1.12u PD=2.16u
M$93 \$232 A|Y$11 25|VSS 25|VSS sg13_lv_nmos L=0.13u W=0.42u AS=0.1428p
+ AD=0.0798p PS=1.52u PD=0.8u
M$94 25|VSS \$232 \$233 25|VSS sg13_lv_nmos L=0.5u W=0.42u AS=0.0798p
+ AD=0.1428p PS=0.8u PD=1.52u
M$95 25|VSS \$233 \$234 25|VSS sg13_lv_nmos L=0.5u W=0.42u AS=0.1426p
+ AD=0.1428p PS=1.16u PD=1.52u
M$96 25|VSS \$234 A|X$15 25|VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.1426p
+ AD=0.2516p PS=1.16u PD=2.16u
M$97 \$235 A|X$17 25|VSS 25|VSS sg13_lv_nmos L=0.13u W=0.42u AS=0.1428p
+ AD=0.0798p PS=1.52u PD=0.8u
M$98 25|VSS \$235 \$236 25|VSS sg13_lv_nmos L=0.5u W=0.42u AS=0.0798p
+ AD=0.1428p PS=0.8u PD=1.52u
M$99 25|VSS \$236 \$237 25|VSS sg13_lv_nmos L=0.5u W=0.42u AS=0.1426p
+ AD=0.1428p PS=1.16u PD=1.52u
M$100 25|VSS \$237 A|X$16 25|VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.1426p
+ AD=0.2516p PS=1.16u PD=2.16u
M$101 25|VSS A|B|Y$4 A|Y$8 25|VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.259p
+ AD=0.259p PS=2.18u PD=2.18u
M$102 25|VSS A|X$18 A|B|Y$3 25|VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.259p
+ AD=0.259p PS=2.18u PD=2.18u
M$103 \$255 \$245 25|VSS 25|VSS sg13_lv_nmos L=0.5u W=0.42u AS=0.1428p
+ AD=0.1426p PS=1.52u PD=1.16u
M$104 25|VSS \$255 A|X$7 25|VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.1426p
+ AD=0.2516p PS=1.16u PD=2.16u
M$105 \$256 \$247 25|VSS 25|VSS sg13_lv_nmos L=0.5u W=0.42u AS=0.1428p
+ AD=0.1426p PS=1.52u PD=1.16u
M$106 25|VSS \$256 A|B|X 25|VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.1426p
+ AD=0.2516p PS=1.16u PD=2.16u
M$107 25|VSS A|Y$10 A|Y$9 25|VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.2516p
+ AD=0.1406p PS=2.16u PD=1.12u
M$108 A|Y$9 A|B|X 25|VSS 25|VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.1406p
+ AD=0.2516p PS=1.12u PD=2.16u
M$109 25|VSS A|B|Y$4 A|Y$11 25|VSS sg13_lv_nmos L=0.13u W=5.92u AS=1.2395p
+ AD=1.2395p PS=10.01u PD=10.01u
M$117 \$257 \$251 25|VSS 25|VSS sg13_lv_nmos L=0.5u W=0.42u AS=0.1428p
+ AD=0.1426p PS=1.52u PD=1.16u
M$118 25|VSS \$257 A|X$19 25|VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.1426p
+ AD=0.2516p PS=1.16u PD=2.16u
M$119 \$238 A|Y$8 \$239 25|VSS sg13_lv_nmos L=0.13u W=0.64u AS=0.2176p
+ AD=0.1216p PS=1.96u PD=1.02u
M$120 25|VSS A|B|Y$3 \$239 25|VSS sg13_lv_nmos L=0.13u W=0.64u AS=0.1331p
+ AD=0.1216p PS=1.12u PD=1.02u
M$121 25|VSS \$238 X 25|VSS sg13_lv_nmos L=0.13u W=1.48u AS=0.2737p AD=0.4218p
+ PS=2.24u PD=3.36u
M$123 \$258 \$254 25|VSS 25|VSS sg13_lv_nmos L=0.5u W=0.42u AS=0.1428p
+ AD=0.1426p PS=1.52u PD=1.16u
M$124 25|VSS \$258 A|X$18 25|VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.1426p
+ AD=0.2516p PS=1.16u PD=2.16u
M$125 \$244 A|X$14 25|VSS 25|VSS sg13_lv_nmos L=0.13u W=0.42u AS=0.1428p
+ AD=0.0798p PS=1.52u PD=0.8u
M$126 25|VSS \$244 \$245 25|VSS sg13_lv_nmos L=0.5u W=0.42u AS=0.0798p
+ AD=0.1428p PS=0.8u PD=1.52u
M$127 25|VSS A|Y$13 A|Y$14 25|VSS sg13_lv_nmos L=0.13u W=1.48u AS=0.3922p
+ AD=0.3959p PS=3.28u PD=3.29u
M$129 \$246 A|X$13 25|VSS 25|VSS sg13_lv_nmos L=0.13u W=0.42u AS=0.1428p
+ AD=0.0798p PS=1.52u PD=0.8u
M$130 25|VSS \$246 \$247 25|VSS sg13_lv_nmos L=0.5u W=0.42u AS=0.0798p
+ AD=0.1428p PS=0.8u PD=1.52u
M$131 25|VSS A|B|X A|Y$13 25|VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.259p
+ AD=0.259p PS=2.18u PD=2.18u
M$132 \$260 A|X$19 25|VSS 25|VSS sg13_lv_nmos L=0.13u W=0.42u AS=0.1428p
+ AD=0.0798p PS=1.52u PD=0.8u
M$133 25|VSS \$260 \$261 25|VSS sg13_lv_nmos L=0.5u W=0.42u AS=0.0798p
+ AD=0.1428p PS=0.8u PD=1.52u
M$134 25|VSS \$261 \$262 25|VSS sg13_lv_nmos L=0.5u W=0.42u AS=0.1426p
+ AD=0.1428p PS=1.16u PD=1.52u
M$135 25|VSS \$262 A|X$17 25|VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.1426p
+ AD=0.2516p PS=1.16u PD=2.16u
M$136 \$250 A|X$15 25|VSS 25|VSS sg13_lv_nmos L=0.13u W=0.42u AS=0.1428p
+ AD=0.0798p PS=1.52u PD=0.8u
M$137 25|VSS \$250 \$251 25|VSS sg13_lv_nmos L=0.5u W=0.42u AS=0.0798p
+ AD=0.1428p PS=0.8u PD=1.52u
M$138 25|VSS A|Y$12 A|B|Y$4 25|VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.259p
+ AD=0.259p PS=2.18u PD=2.18u
M$139 25|VSS 13|A|VINR A|Y$12 25|VSS sg13_lv_nmos L=0.13u W=1.48u AS=0.3922p
+ AD=0.3959p PS=3.28u PD=3.29u
M$141 \$253 A|X$16 25|VSS 25|VSS sg13_lv_nmos L=0.13u W=0.42u AS=0.1428p
+ AD=0.0798p PS=1.52u PD=0.8u
M$142 25|VSS \$253 \$254 25|VSS sg13_lv_nmos L=0.5u W=0.42u AS=0.0798p
+ AD=0.1428p PS=0.8u PD=1.52u
M$143 25|VSS A|Y$14 18|VCP|Y 25|VSS sg13_lv_nmos L=0.13u W=2.96u AS=0.6734p
+ AD=0.6734p PS=5.52u PD=5.52u
M$147 \$300 18|VCP|Y 25|VSS 25|VSS sg13_lv_nmos L=0.13u W=2.24u AS=1.0528p
+ AD=1.0528p PS=5.24u PD=5.24u
M$149 \$301 17|VCN|Y 25|VSS 25|VSS sg13_lv_nmos L=0.13u W=2.24u AS=1.0528p
+ AD=1.0528p PS=5.24u PD=5.24u
M$151 22 \$292 20 20 sg13_hv_nmos L=0.45u W=2000u AS=510.4p AD=510.4p
+ PS=2142.08u PD=2142.08u
M$251 21 \$293 20 20 sg13_hv_nmos L=0.45u W=2000u AS=510.4p AD=510.4p
+ PS=2142.08u PD=2142.08u
M$551 20 20 20 20 sg13_hv_nmos L=0.45u W=1160u AS=300.4p AD=300.4p PS=1260.08u
+ PD=1260.08u
M$608 20 18|VCP|Y \$292 20 sg13_hv_nmos L=0.45u W=250u AS=62.5p AD=62.5p
+ PS=262.5u PD=262.5u
M$633 \$292 20 20 20 sg13_hv_nmos L=0.45u W=10u AS=2.5p AD=2.5p PS=10.5u
+ PD=10.5u
M$634 20 20 \$296 20 sg13_hv_nmos L=0.45u W=20u AS=5p AD=5p PS=21u PD=21u
M$635 \$296 \$300 20 20 sg13_hv_nmos L=0.45u W=60u AS=15p AD=15p PS=63u PD=63u
M$642 20 20 \$297 20 sg13_hv_nmos L=0.45u W=20u AS=5p AD=5p PS=21u PD=21u
M$643 \$297 18|VCP|Y 20 20 sg13_hv_nmos L=0.45u W=60u AS=15p AD=15p PS=63u
+ PD=63u
M$708 20 17|VCN|Y \$293 20 sg13_hv_nmos L=0.45u W=250u AS=62.5p AD=62.5p
+ PS=262.5u PD=262.5u
M$733 \$293 20 20 20 sg13_hv_nmos L=0.45u W=10u AS=2.5p AD=2.5p PS=10.5u
+ PD=10.5u
M$734 20 20 \$298 20 sg13_hv_nmos L=0.45u W=20u AS=5p AD=5p PS=21u PD=21u
M$735 \$298 \$301 20 20 sg13_hv_nmos L=0.45u W=60u AS=15p AD=15p PS=63u PD=63u
M$742 20 20 \$299 20 sg13_hv_nmos L=0.45u W=20u AS=5p AD=5p PS=21u PD=21u
M$743 \$299 17|VCN|Y 20 20 sg13_hv_nmos L=0.45u W=60u AS=15p AD=15p PS=63u
+ PD=63u
M$751 27 21 26 26 sg13_hv_nmos L=0.45u W=40800u AS=14616p AD=14616p PS=44523.2u
+ PD=44523.2u
M$4831 19|VDD A|Y 17|VCN|Y 19|VDD sg13_lv_pmos L=0.13u W=4.48u AS=1.0192p
+ AD=1.0192p PS=7.42u PD=7.42u
M$4835 \$151 \$150 19|VDD 19|VDD sg13_lv_pmos L=0.5u W=1u AS=0.34p AD=0.2254p
+ PS=2.68u PD=1.53u
M$4836 19|VDD \$151 A|X 19|VDD sg13_lv_pmos L=0.13u W=1.12u AS=0.2254p
+ AD=0.4256p PS=1.53u PD=3u
M$4837 \$156 \$155 19|VDD 19|VDD sg13_lv_pmos L=0.5u W=1u AS=0.34p AD=0.2254p
+ PS=2.68u PD=1.53u
M$4838 19|VDD \$156 A|X$2 19|VDD sg13_lv_pmos L=0.13u W=1.12u AS=0.2254p
+ AD=0.4256p PS=1.53u PD=3u
M$4839 19|VDD 14|A|VINS A|Y$1 19|VDD sg13_lv_pmos L=0.13u W=2.24u AS=0.5964p
+ AD=0.5964p PS=4.425u PD=4.425u
M$4841 19|VDD A|Y$2 \$149 19|VDD sg13_lv_pmos L=0.13u W=0.42u AS=0.1523p
+ AD=0.1428p PS=1.38u PD=1.52u
M$4842 19|VDD \$149 \$150 19|VDD sg13_lv_pmos L=0.5u W=1u AS=0.1523p AD=0.34p
+ PS=1.38u PD=2.68u
M$4843 19|VDD A|X$1 \$153 19|VDD sg13_lv_pmos L=0.13u W=0.42u AS=0.1523p
+ AD=0.1428p PS=1.38u PD=1.52u
M$4844 19|VDD \$153 \$155 19|VDD sg13_lv_pmos L=0.5u W=1u AS=0.1523p AD=0.34p
+ PS=1.38u PD=2.68u
M$4845 19|VDD A|Y$1 A|B|Y 19|VDD sg13_lv_pmos L=0.13u W=1.12u AS=0.392p
+ AD=0.392p PS=2.94u PD=2.94u
M$4846 19|VDD A|X$3 A|Y 19|VDD sg13_lv_pmos L=0.13u W=2.24u AS=0.5964p
+ AD=0.5964p PS=4.425u PD=4.425u
M$4848 19|VDD A|B|Y A|Y$2 19|VDD sg13_lv_pmos L=0.13u W=8.96u AS=1.876p
+ AD=1.876p PS=13.43u PD=13.43u
M$4856 19|VDD A|X$4 \$161 19|VDD sg13_lv_pmos L=0.13u W=0.42u AS=0.1523p
+ AD=0.1428p PS=1.38u PD=1.52u
M$4857 19|VDD \$161 \$163 19|VDD sg13_lv_pmos L=0.5u W=1u AS=0.1523p AD=0.34p
+ PS=1.38u PD=2.68u
M$4858 19|VDD \$163 \$164 19|VDD sg13_lv_pmos L=0.5u W=1u AS=0.2254p AD=0.34p
+ PS=1.53u PD=2.68u
M$4859 19|VDD \$164 A|X$1 19|VDD sg13_lv_pmos L=0.13u W=1.12u AS=0.2254p
+ AD=0.4256p PS=1.53u PD=3u
M$4860 19|VDD A|X$5 A|B|Y$1 19|VDD sg13_lv_pmos L=0.13u W=1.12u AS=0.392p
+ AD=0.392p PS=2.94u PD=2.94u
M$4861 \$180 \$168 19|VDD 19|VDD sg13_lv_pmos L=0.5u W=1u AS=0.34p AD=0.2254p
+ PS=2.68u PD=1.53u
M$4862 19|VDD \$180 A|X$6 19|VDD sg13_lv_pmos L=0.13u W=1.12u AS=0.2254p
+ AD=0.4256p PS=1.53u PD=3u
M$4863 \$182 \$171 19|VDD 19|VDD sg13_lv_pmos L=0.5u W=1u AS=0.34p AD=0.2254p
+ PS=2.68u PD=1.53u
M$4864 19|VDD \$182 A|X$3 19|VDD sg13_lv_pmos L=0.13u W=1.12u AS=0.2254p
+ AD=0.4256p PS=1.53u PD=3u
M$4865 19|VDD A|Y$3 \$183 19|VDD sg13_lv_pmos L=0.13u W=0.84u AS=0.2856p
+ AD=0.1596p PS=2.36u PD=1.22u
M$4866 19|VDD A|B|Y \$183 19|VDD sg13_lv_pmos L=0.13u W=0.84u AS=0.1918p
+ AD=0.1596p PS=1.5u PD=1.22u
M$4867 19|VDD \$183 B|X 19|VDD sg13_lv_pmos L=0.13u W=2.24u AS=0.4046p
+ AD=0.6384p PS=3u PD=4.5u
M$4869 \$184 \$175 19|VDD 19|VDD sg13_lv_pmos L=0.5u W=1u AS=0.34p AD=0.2254p
+ PS=2.68u PD=1.53u
M$4870 19|VDD \$184 A|X$4 19|VDD sg13_lv_pmos L=0.13u W=1.12u AS=0.2254p
+ AD=0.4256p PS=1.53u PD=3u
M$4871 \$185 \$177 19|VDD 19|VDD sg13_lv_pmos L=0.5u W=1u AS=0.34p AD=0.2254p
+ PS=2.68u PD=1.53u
M$4872 19|VDD \$185 A|X$5 19|VDD sg13_lv_pmos L=0.13u W=1.12u AS=0.2254p
+ AD=0.4256p PS=1.53u PD=3u
M$4873 19|VDD A|B|Y$1 A|Y$3 19|VDD sg13_lv_pmos L=0.13u W=1.12u AS=0.392p
+ AD=0.392p PS=2.94u PD=2.94u
M$4874 19|VDD A|B|Y A|Y$4 19|VDD sg13_lv_pmos L=0.13u W=1.12u AS=0.392p
+ AD=0.392p PS=2.94u PD=2.94u
M$4875 19|VDD A|Y$5 \$190 19|VDD sg13_lv_pmos L=0.13u W=0.42u AS=0.1523p
+ AD=0.1428p PS=1.38u PD=1.52u
M$4876 19|VDD \$190 \$191 19|VDD sg13_lv_pmos L=0.5u W=1u AS=0.1523p AD=0.34p
+ PS=1.38u PD=2.68u
M$4877 19|VDD \$191 \$205 19|VDD sg13_lv_pmos L=0.5u W=1u AS=0.2254p AD=0.34p
+ PS=1.53u PD=2.68u
M$4878 19|VDD \$205 A|X$9 19|VDD sg13_lv_pmos L=0.13u W=1.12u AS=0.2254p
+ AD=0.4256p PS=1.53u PD=3u
M$4879 19|VDD A|X$7 \$167 19|VDD sg13_lv_pmos L=0.13u W=0.42u AS=0.1523p
+ AD=0.1428p PS=1.38u PD=1.52u
M$4880 19|VDD \$167 \$168 19|VDD sg13_lv_pmos L=0.5u W=1u AS=0.1523p AD=0.34p
+ PS=1.38u PD=2.68u
M$4881 19|VDD A|X$12 \$193 19|VDD sg13_lv_pmos L=0.13u W=0.42u AS=0.1523p
+ AD=0.1428p PS=1.38u PD=1.52u
M$4882 19|VDD \$193 \$194 19|VDD sg13_lv_pmos L=0.5u W=1u AS=0.1523p AD=0.34p
+ PS=1.38u PD=2.68u
M$4883 19|VDD \$194 \$207 19|VDD sg13_lv_pmos L=0.5u W=1u AS=0.2254p AD=0.34p
+ PS=1.53u PD=2.68u
M$4884 19|VDD \$207 A|X$10 19|VDD sg13_lv_pmos L=0.13u W=1.12u AS=0.2254p
+ AD=0.4256p PS=1.53u PD=3u
M$4885 19|VDD A|X$8 \$170 19|VDD sg13_lv_pmos L=0.13u W=0.42u AS=0.1523p
+ AD=0.1428p PS=1.38u PD=1.52u
M$4886 19|VDD \$170 \$171 19|VDD sg13_lv_pmos L=0.5u W=1u AS=0.1523p AD=0.34p
+ PS=1.38u PD=2.68u
M$4887 19|VDD A|X$6 \$196 19|VDD sg13_lv_pmos L=0.13u W=0.42u AS=0.1523p
+ AD=0.1428p PS=1.38u PD=1.52u
M$4888 19|VDD \$196 \$197 19|VDD sg13_lv_pmos L=0.5u W=1u AS=0.1523p AD=0.34p
+ PS=1.38u PD=2.68u
M$4889 19|VDD \$197 \$208 19|VDD sg13_lv_pmos L=0.5u W=1u AS=0.2254p AD=0.34p
+ PS=1.53u PD=2.68u
M$4890 19|VDD \$208 A|X$8 19|VDD sg13_lv_pmos L=0.13u W=1.12u AS=0.2254p
+ AD=0.4256p PS=1.53u PD=3u
M$4891 19|VDD A|X$3 \$213 19|VDD sg13_lv_pmos L=0.13u W=1.12u AS=0.4032p
+ AD=0.1176p PS=2.96u PD=1.33u
M$4892 \$213 A|B|Y$2 A|Y$5 19|VDD sg13_lv_pmos L=0.13u W=1.12u AS=0.1176p
+ AD=0.3808p PS=1.33u PD=2.92u
M$4893 19|VDD A|Y$7 \$212 19|VDD sg13_lv_pmos L=0.13u W=1.12u AS=0.4032p
+ AD=0.1176p PS=2.96u PD=1.33u
M$4894 \$212 B|X A|B|Y$2 19|VDD sg13_lv_pmos L=0.13u W=1.12u AS=0.1176p
+ AD=0.3808p PS=1.33u PD=2.92u
M$4895 19|VDD A|X \$174 19|VDD sg13_lv_pmos L=0.13u W=0.42u AS=0.1523p
+ AD=0.1428p PS=1.38u PD=1.52u
M$4896 19|VDD \$174 \$175 19|VDD sg13_lv_pmos L=0.5u W=1u AS=0.1523p AD=0.34p
+ PS=1.38u PD=2.68u
M$4897 19|VDD A|Y$6 \$199 19|VDD sg13_lv_pmos L=0.13u W=0.84u AS=0.2856p
+ AD=0.1596p PS=2.36u PD=1.22u
M$4898 \$199 A|B|Y$4 19|VDD 19|VDD sg13_lv_pmos L=0.13u W=0.84u AS=0.1596p
+ AD=0.1918p PS=1.22u PD=1.5u
M$4899 19|VDD \$199 A|X$11 19|VDD sg13_lv_pmos L=0.13u W=2.24u AS=0.4046p
+ AD=0.6384p PS=3u PD=4.5u
M$4901 19|VDD A|Y$4 \$201 19|VDD sg13_lv_pmos L=0.13u W=0.84u AS=0.2856p
+ AD=0.1596p PS=2.36u PD=1.22u
M$4902 \$201 A|B|Y$1 19|VDD 19|VDD sg13_lv_pmos L=0.13u W=0.84u AS=0.1596p
+ AD=0.1918p PS=1.22u PD=1.5u
M$4903 19|VDD \$201 X 19|VDD sg13_lv_pmos L=0.13u W=2.24u AS=0.4046p AD=0.6384p
+ PS=3u PD=4.5u
M$4905 19|VDD A|X$2 \$176 19|VDD sg13_lv_pmos L=0.13u W=0.42u AS=0.1523p
+ AD=0.1428p PS=1.38u PD=1.52u
M$4906 19|VDD \$176 \$177 19|VDD sg13_lv_pmos L=0.5u W=1u AS=0.1523p AD=0.34p
+ PS=1.38u PD=2.68u
M$4907 19|VDD A|B|Y$3 A|Y$6 19|VDD sg13_lv_pmos L=0.13u W=1.12u AS=0.392p
+ AD=0.392p PS=2.94u PD=2.94u
M$4908 \$223 \$222 19|VDD 19|VDD sg13_lv_pmos L=0.5u W=1u AS=0.34p AD=0.2254p
+ PS=2.68u PD=1.53u
M$4909 19|VDD \$223 A|X$12 19|VDD sg13_lv_pmos L=0.13u W=1.12u AS=0.2254p
+ AD=0.4256p PS=1.53u PD=3u
M$4910 \$226 \$225 19|VDD 19|VDD sg13_lv_pmos L=0.5u W=1u AS=0.34p AD=0.2254p
+ PS=2.68u PD=1.53u
M$4911 19|VDD \$226 A|X$13 19|VDD sg13_lv_pmos L=0.13u W=1.12u AS=0.2254p
+ AD=0.4256p PS=1.53u PD=3u
M$4912 \$230 \$229 19|VDD 19|VDD sg13_lv_pmos L=0.5u W=1u AS=0.34p AD=0.2254p
+ PS=2.68u PD=1.53u
M$4913 19|VDD \$230 A|X$14 19|VDD sg13_lv_pmos L=0.13u W=1.12u AS=0.2254p
+ AD=0.4256p PS=1.53u PD=3u
M$4914 19|VDD A|B|Y$2 A|Y$10 19|VDD sg13_lv_pmos L=0.13u W=1.12u AS=0.392p
+ AD=0.392p PS=2.94u PD=2.94u
M$4915 19|VDD A|X$11 \$242 19|VDD sg13_lv_pmos L=0.13u W=1.12u AS=0.4032p
+ AD=0.1176p PS=2.96u PD=1.33u
M$4916 \$242 A|B|Y$2 A|Y$7 19|VDD sg13_lv_pmos L=0.13u W=1.12u AS=0.1176p
+ AD=0.3808p PS=1.33u PD=2.92u
M$4917 \$234 \$233 19|VDD 19|VDD sg13_lv_pmos L=0.5u W=1u AS=0.34p AD=0.2254p
+ PS=2.68u PD=1.53u
M$4918 19|VDD \$234 A|X$15 19|VDD sg13_lv_pmos L=0.13u W=1.12u AS=0.2254p
+ AD=0.4256p PS=1.53u PD=3u
M$4919 \$237 \$236 19|VDD 19|VDD sg13_lv_pmos L=0.5u W=1u AS=0.34p AD=0.2254p
+ PS=2.68u PD=1.53u
M$4920 19|VDD \$237 A|X$16 19|VDD sg13_lv_pmos L=0.13u W=1.12u AS=0.2254p
+ AD=0.4256p PS=1.53u PD=3u
M$4921 19|VDD A|Y$8 \$238 19|VDD sg13_lv_pmos L=0.13u W=0.84u AS=0.2856p
+ AD=0.1596p PS=2.36u PD=1.22u
M$4922 19|VDD A|B|Y$3 \$238 19|VDD sg13_lv_pmos L=0.13u W=0.84u AS=0.1918p
+ AD=0.1596p PS=1.5u PD=1.22u
M$4923 19|VDD \$238 X 19|VDD sg13_lv_pmos L=0.13u W=2.24u AS=0.4046p AD=0.6384p
+ PS=3u PD=4.5u
M$4925 19|VDD A|B|Y$4 A|Y$8 19|VDD sg13_lv_pmos L=0.13u W=1.12u AS=0.392p
+ AD=0.392p PS=2.94u PD=2.94u
M$4926 19|VDD A|X$18 A|B|Y$3 19|VDD sg13_lv_pmos L=0.13u W=1.12u AS=0.392p
+ AD=0.392p PS=2.94u PD=2.94u
M$4927 19|VDD A|X$9 \$221 19|VDD sg13_lv_pmos L=0.13u W=0.42u AS=0.1523p
+ AD=0.1428p PS=1.38u PD=1.52u
M$4928 19|VDD \$221 \$222 19|VDD sg13_lv_pmos L=0.5u W=1u AS=0.1523p AD=0.34p
+ PS=1.38u PD=2.68u
M$4929 19|VDD A|X$14 \$244 19|VDD sg13_lv_pmos L=0.13u W=0.42u AS=0.1523p
+ AD=0.1428p PS=1.38u PD=1.52u
M$4930 19|VDD \$244 \$245 19|VDD sg13_lv_pmos L=0.5u W=1u AS=0.1523p AD=0.34p
+ PS=1.38u PD=2.68u
M$4931 19|VDD \$245 \$255 19|VDD sg13_lv_pmos L=0.5u W=1u AS=0.2254p AD=0.34p
+ PS=1.53u PD=2.68u
M$4932 19|VDD \$255 A|X$7 19|VDD sg13_lv_pmos L=0.13u W=1.12u AS=0.2254p
+ AD=0.4256p PS=1.53u PD=3u
M$4933 19|VDD A|X$10 \$224 19|VDD sg13_lv_pmos L=0.13u W=0.42u AS=0.1523p
+ AD=0.1428p PS=1.38u PD=1.52u
M$4934 19|VDD \$224 \$225 19|VDD sg13_lv_pmos L=0.5u W=1u AS=0.1523p AD=0.34p
+ PS=1.38u PD=2.68u
M$4935 19|VDD A|X$13 \$246 19|VDD sg13_lv_pmos L=0.13u W=0.42u AS=0.1523p
+ AD=0.1428p PS=1.38u PD=1.52u
M$4936 19|VDD \$246 \$247 19|VDD sg13_lv_pmos L=0.5u W=1u AS=0.1523p AD=0.34p
+ PS=1.38u PD=2.68u
M$4937 19|VDD \$247 \$256 19|VDD sg13_lv_pmos L=0.5u W=1u AS=0.2254p AD=0.34p
+ PS=1.53u PD=2.68u
M$4938 19|VDD \$256 A|B|X 19|VDD sg13_lv_pmos L=0.13u W=1.12u AS=0.2254p
+ AD=0.4256p PS=1.53u PD=3u
M$4939 19|VDD A|Y$9 \$227 19|VDD sg13_lv_pmos L=0.13u W=0.42u AS=0.1523p
+ AD=0.1428p PS=1.38u PD=1.52u
M$4940 19|VDD \$227 \$229 19|VDD sg13_lv_pmos L=0.5u W=1u AS=0.1523p AD=0.34p
+ PS=1.38u PD=2.68u
M$4941 19|VDD A|Y$10 \$259 19|VDD sg13_lv_pmos L=0.13u W=1.12u AS=0.4032p
+ AD=0.1176p PS=2.96u PD=1.33u
M$4942 \$259 A|B|X A|Y$9 19|VDD sg13_lv_pmos L=0.13u W=1.12u AS=0.1176p
+ AD=0.3808p PS=1.33u PD=2.92u
M$4943 19|VDD A|Y$11 \$232 19|VDD sg13_lv_pmos L=0.13u W=0.42u AS=0.1523p
+ AD=0.1428p PS=1.38u PD=1.52u
M$4944 19|VDD \$232 \$233 19|VDD sg13_lv_pmos L=0.5u W=1u AS=0.1523p AD=0.34p
+ PS=1.38u PD=2.68u
M$4945 19|VDD A|B|Y$4 A|Y$11 19|VDD sg13_lv_pmos L=0.13u W=8.96u AS=1.876p
+ AD=1.876p PS=13.43u PD=13.43u
M$4953 19|VDD A|X$17 \$235 19|VDD sg13_lv_pmos L=0.13u W=0.42u AS=0.1523p
+ AD=0.1428p PS=1.38u PD=1.52u
M$4954 19|VDD \$235 \$236 19|VDD sg13_lv_pmos L=0.5u W=1u AS=0.1523p AD=0.34p
+ PS=1.38u PD=2.68u
M$4955 19|VDD A|X$15 \$250 19|VDD sg13_lv_pmos L=0.13u W=0.42u AS=0.1523p
+ AD=0.1428p PS=1.38u PD=1.52u
M$4956 19|VDD \$250 \$251 19|VDD sg13_lv_pmos L=0.5u W=1u AS=0.1523p AD=0.34p
+ PS=1.38u PD=2.68u
M$4957 19|VDD \$251 \$257 19|VDD sg13_lv_pmos L=0.5u W=1u AS=0.2254p AD=0.34p
+ PS=1.53u PD=2.68u
M$4958 19|VDD \$257 A|X$19 19|VDD sg13_lv_pmos L=0.13u W=1.12u AS=0.2254p
+ AD=0.4256p PS=1.53u PD=3u
M$4959 19|VDD A|X$16 \$253 19|VDD sg13_lv_pmos L=0.13u W=0.42u AS=0.1523p
+ AD=0.1428p PS=1.38u PD=1.52u
M$4960 19|VDD \$253 \$254 19|VDD sg13_lv_pmos L=0.5u W=1u AS=0.1523p AD=0.34p
+ PS=1.38u PD=2.68u
M$4961 19|VDD \$254 \$258 19|VDD sg13_lv_pmos L=0.5u W=1u AS=0.2254p AD=0.34p
+ PS=1.53u PD=2.68u
M$4962 19|VDD \$258 A|X$18 19|VDD sg13_lv_pmos L=0.13u W=1.12u AS=0.2254p
+ AD=0.4256p PS=1.53u PD=3u
M$4963 19|VDD A|Y$14 18|VCP|Y 19|VDD sg13_lv_pmos L=0.13u W=4.48u AS=1.0192p
+ AD=1.0192p PS=7.42u PD=7.42u
M$4967 19|VDD A|Y$13 A|Y$14 19|VDD sg13_lv_pmos L=0.13u W=2.24u AS=0.5964p
+ AD=0.5964p PS=4.425u PD=4.425u
M$4969 19|VDD A|B|X A|Y$13 19|VDD sg13_lv_pmos L=0.13u W=1.12u AS=0.392p
+ AD=0.392p PS=2.94u PD=2.94u
M$4970 19|VDD A|X$19 \$260 19|VDD sg13_lv_pmos L=0.13u W=0.42u AS=0.1523p
+ AD=0.1428p PS=1.38u PD=1.52u
M$4971 19|VDD \$260 \$261 19|VDD sg13_lv_pmos L=0.5u W=1u AS=0.1523p AD=0.34p
+ PS=1.38u PD=2.68u
M$4972 \$262 \$261 19|VDD 19|VDD sg13_lv_pmos L=0.5u W=1u AS=0.34p AD=0.2254p
+ PS=2.68u PD=1.53u
M$4973 19|VDD \$262 A|X$17 19|VDD sg13_lv_pmos L=0.13u W=1.12u AS=0.2254p
+ AD=0.4256p PS=1.53u PD=3u
M$4974 19|VDD A|Y$12 A|B|Y$4 19|VDD sg13_lv_pmos L=0.13u W=1.12u AS=0.392p
+ AD=0.392p PS=2.94u PD=2.94u
M$4975 19|VDD 13|A|VINR A|Y$12 19|VDD sg13_lv_pmos L=0.13u W=2.24u AS=0.5964p
+ AD=0.5964p PS=4.425u PD=4.425u
M$4977 \$300 18|VCP|Y 19|VDD 19|VDD sg13_lv_pmos L=0.13u W=2.24u AS=1.0528p
+ AD=1.0528p PS=5.24u PD=5.24u
M$4979 \$301 17|VCN|Y 19|VDD 19|VDD sg13_lv_pmos L=0.13u W=2.24u AS=1.0528p
+ AD=1.0528p PS=5.24u PD=5.24u
M$4981 27 22 28 28 sg13_hv_pmos L=0.4u W=120960u AS=44217.6p AD=44217.6p
+ PS=134283.52u PD=134283.52u
M$8383 22 \$292 23 23 sg13_hv_pmos L=0.4u W=2500u AS=638p AD=638p PS=2677.6u
+ PD=2677.6u
M$8433 23 23 23 23 sg13_hv_pmos L=0.4u W=280u AS=75.2p AD=75.2p PS=315.04u
+ PD=315.04u
M$8436 23 23 \$292 23 sg13_hv_pmos L=0.4u W=20u AS=5p AD=5p PS=21u PD=21u
M$8437 \$292 \$296 23 23 sg13_hv_pmos L=0.4u W=300u AS=75p AD=75p PS=315u
+ PD=315u
M$8469 23 23 \$296 23 sg13_hv_pmos L=0.4u W=10u AS=2.5p AD=2.5p PS=10.5u
+ PD=10.5u
M$8470 \$296 \$297 23 23 sg13_hv_pmos L=0.4u W=10u AS=2.5p AD=2.5p PS=10.5u
+ PD=10.5u
M$8479 23 23 \$297 23 sg13_hv_pmos L=0.4u W=10u AS=2.5p AD=2.5p PS=10.5u
+ PD=10.5u
M$8480 \$297 \$296 23 23 sg13_hv_pmos L=0.4u W=10u AS=2.5p AD=2.5p PS=10.5u
+ PD=10.5u
M$8483 21 \$293 23 23 sg13_hv_pmos L=0.4u W=2500u AS=638p AD=638p PS=2677.6u
+ PD=2677.6u
M$8536 23 23 \$293 23 sg13_hv_pmos L=0.4u W=20u AS=5p AD=5p PS=21u PD=21u
M$8537 \$293 \$298 23 23 sg13_hv_pmos L=0.4u W=300u AS=75p AD=75p PS=315u
+ PD=315u
M$8569 23 23 \$298 23 sg13_hv_pmos L=0.4u W=10u AS=2.5p AD=2.5p PS=10.5u
+ PD=10.5u
M$8570 \$298 \$299 23 23 sg13_hv_pmos L=0.4u W=10u AS=2.5p AD=2.5p PS=10.5u
+ PD=10.5u
M$8579 23 23 \$299 23 sg13_hv_pmos L=0.4u W=10u AS=2.5p AD=2.5p PS=10.5u
+ PD=10.5u
M$8580 \$299 \$298 23 23 sg13_hv_pmos L=0.4u W=10u AS=2.5p AD=2.5p PS=10.5u
+ PD=10.5u
D$17677 25|VSS 28 8 diodevdd_2kv m=1
D$17678 25|VSS 28 9 diodevdd_2kv m=1
D$17679 25|VSS 28 10 diodevdd_2kv m=1
D$17680 25|VSS 28 11 diodevdd_2kv m=1
D$17681 25|VSS 28 12 diodevdd_2kv m=1
D$17682 25|VSS 28 13|A|VINR diodevdd_2kv m=1
D$17683 25|VSS 28 14|A|VINS diodevdd_2kv m=1
D$17684 25|VSS 28 7 diodevdd_2kv m=1
D$17685 25|VSS 28 15 diodevdd_2kv m=1
D$17686 25|VSS 28 6 diodevdd_2kv m=1
D$17687 25|VSS 28 16 diodevdd_2kv m=1
D$17688 25|VSS 28 5 diodevdd_2kv m=1
D$17689 25|VSS 28 17|VCN|Y diodevdd_2kv m=1
D$17690 25|VSS 28 4 diodevdd_2kv m=1
D$17691 25|VSS 28 18|VCP|Y diodevdd_2kv m=1
D$17692 25|VSS 28 3 diodevdd_2kv m=1
D$17693 25|VSS 28 19|VDD diodevdd_2kv m=1
D$17694 25|VSS 28 2 diodevdd_2kv m=1
D$17695 25|VSS 28 20 diodevdd_2kv m=1
D$17696 25|VSS 28 1 diodevdd_2kv m=1
D$17697 25|VSS 28 21 diodevdd_2kv m=1
D$17698 25|VSS 28 28 diodevdd_2kv m=1
D$17699 25|VSS 28 27 diodevdd_2kv m=1
D$17700 25|VSS 28 26 diodevdd_2kv m=1
D$17701 25|VSS 28 25|VSS diodevdd_2kv m=1
D$17702 25|VSS 28 24 diodevdd_2kv m=1
D$17703 25|VSS 28 23 diodevdd_2kv m=1
D$17704 25|VSS 28 22 diodevdd_2kv m=1
D$17705 28 25|VSS 8 diodevss_2kv m=1
D$17706 28 25|VSS 9 diodevss_2kv m=1
D$17707 28 25|VSS 10 diodevss_2kv m=1
D$17708 28 25|VSS 11 diodevss_2kv m=1
D$17709 28 25|VSS 12 diodevss_2kv m=1
D$17710 28 25|VSS 13|A|VINR diodevss_2kv m=1
D$17711 28 25|VSS 14|A|VINS diodevss_2kv m=1
D$17712 28 25|VSS 7 diodevss_2kv m=1
D$17713 28 25|VSS 15 diodevss_2kv m=1
D$17714 28 25|VSS 6 diodevss_2kv m=1
D$17715 28 25|VSS 16 diodevss_2kv m=1
D$17716 28 25|VSS 5 diodevss_2kv m=1
D$17717 28 25|VSS 17|VCN|Y diodevss_2kv m=1
D$17718 28 25|VSS 4 diodevss_2kv m=1
D$17719 28 25|VSS 18|VCP|Y diodevss_2kv m=1
D$17720 28 25|VSS 3 diodevss_2kv m=1
D$17721 28 25|VSS 19|VDD diodevss_2kv m=1
D$17722 28 25|VSS 2 diodevss_2kv m=1
D$17723 28 25|VSS 20 diodevss_2kv m=1
D$17724 28 25|VSS 1 diodevss_2kv m=1
D$17725 28 25|VSS 21 diodevss_2kv m=1
D$17726 28 25|VSS 28 diodevss_2kv m=1
D$17727 28 25|VSS 27 diodevss_2kv m=1
D$17728 28 25|VSS 26 diodevss_2kv m=1
D$17729 28 25|VSS 25|VSS diodevss_2kv m=1
D$17730 28 25|VSS 24 diodevss_2kv m=1
D$17731 28 25|VSS 23 diodevss_2kv m=1
D$17732 28 25|VSS 22 diodevss_2kv m=1
.ENDS AC3E_USM_TDBUCK
