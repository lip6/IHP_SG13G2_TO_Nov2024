** sch_path: /home/Joerdson/IHP-Open-PDK/ihp-sg13g2/libs.tech/xschem/CryoChip.sch
**.subckt CryoChip SN1 DN1 GN1 SN2 DN2 GN2 SN3 DN3 GN3 SN4 DN4 GN4 SN5 DN5 GN5 SN6 DN6 GN6 SN7 DN7 GN7 SN8 DN8 GN8 OUT IN VDD BP1
*+ SP1 DP1 GP1 BP2 SP2 DP2 GP2 BP3 SP3 DP3 GP3 BP4 SP4 DP4 GP4 BP5 SP5 DP5 GP5 BP6 SP6 DP6 GP6 BP7 SP7 DP7 GP7 BP8 SP8 DP8 GP8 GPN SDP1
*+ SDP2 SDP3 SDP4 SDP5 SDN5 SDN4 SDN3 SDN2 SDN1 SDN0 SDP6 SDP0 SDN6 BP BN
*.iopin SN1
*.iopin DN1
*.iopin GN1
*.iopin SN2
*.iopin DN2
*.iopin GN2
*.iopin SN3
*.iopin DN3
*.iopin GN3
*.iopin SN4
*.iopin DN4
*.iopin GN4
*.iopin SN5
*.iopin DN5
*.iopin GN5
*.iopin SN6
*.iopin DN6
*.iopin GN6
*.iopin SN7
*.iopin DN7
*.iopin GN7
*.iopin SN8
*.iopin DN8
*.iopin GN8
*.iopin OUT
*.iopin IN
*.iopin VDD
*.iopin BP1
*.iopin SP1
*.iopin DP1
*.iopin GP1
*.iopin BP2
*.iopin SP2
*.iopin DP2
*.iopin GP2
*.iopin BP3
*.iopin SP3
*.iopin DP3
*.iopin GP3
*.iopin BP4
*.iopin SP4
*.iopin DP4
*.iopin GP4
*.iopin BP5
*.iopin SP5
*.iopin DP5
*.iopin GP5
*.iopin BP6
*.iopin SP6
*.iopin DP6
*.iopin GP6
*.iopin BP7
*.iopin SP7
*.iopin DP7
*.iopin GP7
*.iopin BP8
*.iopin SP8
*.iopin DP8
*.iopin GP8
*.iopin GPN
*.iopin SDP1
*.iopin SDP2
*.iopin SDP3
*.iopin SDP4
*.iopin SDP5
*.iopin SDN5
*.iopin SDN4
*.iopin SDN3
*.iopin SDN2
*.iopin SDN1
*.iopin SDN0
*.iopin SDP6
*.iopin SDP0
*.iopin SDN6
*.iopin BP
*.iopin BN
XM13 DN1 GN1 SN1 BN sg13_lv_nmos w=0.15u l=0.13u ng=1 m=1
XM14 DN2 GN2 SN2 BN sg13_lv_nmos w=3u l=0.13u ng=1 m=1
XM15 DN3 GN3 SN3 BN sg13_lv_nmos w=3u l=0.3u ng=1 m=1
XM16 DN4 GN4 SN4 BN sg13_lv_nmos w=3u l=0.6u ng=1 m=1
XM17 DN5 GN5 SN5 BN sg13_lv_nmos w=3u l=1u ng=1 m=1
XM18 DN6 GN6 SN6 BN sg13_lv_nmos w=10u l=10u ng=1 m=1
XM19 DN7 GN7 SN7 BN sg13_lv_nmos w=1u l=1u ng=1 m=1
XM20 DN8 GN8 SN8 BN sg13_lv_nmos w=0.5u l=1u ng=1 m=1
XM21 DP1 GP1 SP1 BP1 sg13_lv_pmos w=0.15u l=0.13u ng=1 m=1
XM22 DP2 GP2 SP2 BP2 sg13_lv_pmos w=3.0u l=0.13u ng=1 m=1
XM23 DP3 GP3 SP3 BP3 sg13_lv_pmos w=3.0u l=0.3u ng=1 m=1
XM24 DP4 GP4 SP4 BP4 sg13_lv_pmos w=3.0u l=0.6u ng=1 m=1
XM25 DP5 GP5 SP5 BP5 sg13_lv_pmos w=3u l=1u ng=1 m=1
XM26 DP6 GP6 SP6 BP6 sg13_lv_pmos w=10u l=10u ng=1 m=1
XM27 DP7 GP7 SP7 BP7 sg13_lv_pmos w=1u l=1u ng=1 m=1
XM28 DP8 GP8 SP8 BP8 sg13_lv_pmos w=0.5u l=1u ng=1 m=1
XM29 BN IN OUT BN sg13_lv_nmos w=0.15u l=0.13u ng=1 m=1
XM30 OUT IN VDD VDD sg13_lv_pmos w=0.6u l=0.13u ng=1 m=1
XM1 SDN0 GPN SDN1 BN sg13_lv_nmos w=0.15u l=0.13u ng=1 m=1
XM2 SDP1 GPN SDP0 BP sg13_lv_pmos w=0.15u l=0.13u ng=1 m=1
XM3 SDN1 GPN SDN2 BN sg13_lv_nmos w=3.0u l=0.13u ng=1 m=1
XM4 SDP2 GPN SDP1 BP sg13_lv_pmos w=3.0u l=0.13u ng=1 m=1
XM5 SDN2 GPN SDN3 BN sg13_lv_nmos w=3.0u l=0.3u ng=1 m=1
XM6 SDP3 GPN SDP2 BP sg13_lv_pmos w=3.0u l=0.3u ng=1 m=1
XM7 SDN3 GPN SDN4 BN sg13_lv_nmos w=3.0u l=0.6u ng=1 m=1
XM8 SDP4 GPN SDP3 BP sg13_lv_pmos w=3.0u l=0.6u ng=1 m=1
XM9 SDN4 GPN SDN5 BN sg13_lv_nmos w=3.0u l=1.0u ng=1 m=1
XM10 SDP5 GPN SDP4 BP sg13_lv_pmos w=3.0u l=1.0u ng=1 m=1
XM11 SDN5 GPN SDN6 BN sg13_lv_nmos w=10u l=10u ng=1 m=1
XM12 SDP6 GPN SDP5 BP sg13_lv_pmos w=10u l=10u ng=1 m=1
**.ends
.end
