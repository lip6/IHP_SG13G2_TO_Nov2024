* Extracted by KLayout with SG13G2 LVS runset on : 22/11/2024 07:08

.SUBCKT top 15|25|VSS 24 8 10|A1|VINS_OL 11|A1|VINR_OL 12|S|VSEL_OL
+ 13|S|VSEL_DT 14|VINR_BUFF|X 7 6 16|PD_BUFF|X 2 9 5 17|NOC_N_BUFF|X 1 19|VDD A
+ A$1 A|Y A|Y$1 A|VINS|X A|VINR|X A|X A|X$1 A|X$2 VINS_BUFF|X A|X$3 A$2 A$3
+ A|B|Y A|X$4 A|B|Y$1 A|Y$2 A|X$5 A|X$6 A|Y$3 A|X$7 A|X$8 A|X$9 A|X$10 A|B|Y$2
+ A|X$11 A$4 4 A|X$12 A|Y$4 A|X$13 A|Y$5 A|Y$6 A|Y$7 A|B|Y$3 A|B|Y$4 A|Y$8
+ A|Y$9 X B|X A$5 A|Y$10 A|X$14 A|X$15 A|X$16 A|X$17 A|X$18 A|X$19 A|X$20
+ A|X$21 A|X$22 A|X$23 A|X$24 A$6 A|X$25 A|X$26 A|X$27 A|Y$11 A|X$28 A|X$29
+ A|Y$12 A|X$30 A|X$31 A|X$32 A|X$33 A|X$34 A|X$35 A|X$36 A|Y$13 A|B|X A|Y$14
+ A|Y$15 A|Y$16 A|X$37 A|X$38 A0|Y A|X$39 A|X$40 A|X$41 A|X$42 A|X$43 A0|X
+ A|X$44 A|X$45 A0|Y$1 A1|X A|X$46 A1|X$1 A|X$47 A0|X$1 27 28 18|NOC_P_BUFF|X
+ 23 20 NOC_P|X NOC_N|X 3 26 21 22
M$1 \$245 A|Y 15|25|VSS 15|25|VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.2664p
+ AD=0.3034p PS=2.2u PD=1.56u
M$2 15|25|VSS \$245 A|VINS|X 15|25|VSS sg13_lv_nmos L=0.13u W=2.96u AS=0.7252p
+ AD=0.6734p PS=4.92u PD=5.52u
M$6 15|25|VSS A A|Y 15|25|VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.259p AD=0.259p
+ PS=2.18u PD=2.18u
M$7 \$246 A|Y$1 15|25|VSS 15|25|VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.2664p
+ AD=0.3034p PS=2.2u PD=1.56u
M$8 15|25|VSS \$246 A|VINR|X 15|25|VSS sg13_lv_nmos L=0.13u W=2.96u AS=0.7252p
+ AD=0.6734p PS=4.92u PD=5.52u
M$12 15|25|VSS A$1 A|Y$1 15|25|VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.259p
+ AD=0.259p PS=2.18u PD=2.18u
M$13 15|25|VSS \$259 16|PD_BUFF|X 15|25|VSS sg13_lv_nmos L=0.13u W=11.84u
+ AS=2.3606p AD=2.2496p PS=18.96u PD=17.92u
M$29 15|25|VSS A|X \$259 15|25|VSS sg13_lv_nmos L=0.13u W=4.44u AS=0.8436p
+ AD=0.9546p PS=6.72u PD=7.76u
M$35 15|25|VSS \$261 VINS_BUFF|X 15|25|VSS sg13_lv_nmos L=0.13u W=11.84u
+ AS=2.3606p AD=2.2496p PS=18.96u PD=17.92u
M$51 15|25|VSS A|X$1 \$261 15|25|VSS sg13_lv_nmos L=0.13u W=4.44u AS=0.8436p
+ AD=0.9546p PS=6.72u PD=7.76u
M$57 15|25|VSS \$263 17|NOC_N_BUFF|X 15|25|VSS sg13_lv_nmos L=0.13u W=11.84u
+ AS=2.3606p AD=2.2496p PS=18.96u PD=17.92u
M$73 15|25|VSS A|X$2 \$263 15|25|VSS sg13_lv_nmos L=0.13u W=4.44u AS=0.8436p
+ AD=0.9546p PS=6.72u PD=7.76u
M$79 15|25|VSS \$266 16|PD_BUFF|X 15|25|VSS sg13_lv_nmos L=0.13u W=11.84u
+ AS=2.3606p AD=2.2496p PS=18.96u PD=17.92u
M$95 15|25|VSS A|X \$266 15|25|VSS sg13_lv_nmos L=0.13u W=4.44u AS=0.8436p
+ AD=0.9546p PS=6.72u PD=7.76u
M$101 15|25|VSS \$267 VINS_BUFF|X 15|25|VSS sg13_lv_nmos L=0.13u W=11.84u
+ AS=2.3606p AD=2.2496p PS=18.96u PD=17.92u
M$117 15|25|VSS A|X$1 \$267 15|25|VSS sg13_lv_nmos L=0.13u W=4.44u AS=0.8436p
+ AD=0.9546p PS=6.72u PD=7.76u
M$123 15|25|VSS \$268 17|NOC_N_BUFF|X 15|25|VSS sg13_lv_nmos L=0.13u W=11.84u
+ AS=2.3606p AD=2.2496p PS=18.96u PD=17.92u
M$139 15|25|VSS A|X$2 \$268 15|25|VSS sg13_lv_nmos L=0.13u W=4.44u AS=0.8436p
+ AD=0.9546p PS=6.72u PD=7.76u
M$145 15|25|VSS \$269 16|PD_BUFF|X 15|25|VSS sg13_lv_nmos L=0.13u W=11.84u
+ AS=2.3606p AD=2.2496p PS=18.96u PD=17.92u
M$161 15|25|VSS A|X \$269 15|25|VSS sg13_lv_nmos L=0.13u W=4.44u AS=0.8436p
+ AD=0.9546p PS=6.72u PD=7.76u
M$167 15|25|VSS \$270 VINS_BUFF|X 15|25|VSS sg13_lv_nmos L=0.13u W=11.84u
+ AS=2.3606p AD=2.2496p PS=18.96u PD=17.92u
M$183 15|25|VSS A|X$1 \$270 15|25|VSS sg13_lv_nmos L=0.13u W=4.44u AS=0.8436p
+ AD=0.9546p PS=6.72u PD=7.76u
M$189 15|25|VSS \$271 17|NOC_N_BUFF|X 15|25|VSS sg13_lv_nmos L=0.13u W=11.84u
+ AS=2.3606p AD=2.2496p PS=18.96u PD=17.92u
M$205 15|25|VSS A|X$2 \$271 15|25|VSS sg13_lv_nmos L=0.13u W=4.44u AS=0.8436p
+ AD=0.9546p PS=6.72u PD=7.76u
M$211 15|25|VSS \$272 16|PD_BUFF|X 15|25|VSS sg13_lv_nmos L=0.13u W=11.84u
+ AS=2.3606p AD=2.2496p PS=18.96u PD=17.92u
M$227 15|25|VSS A|X \$272 15|25|VSS sg13_lv_nmos L=0.13u W=4.44u AS=0.8436p
+ AD=0.9546p PS=6.72u PD=7.76u
M$233 15|25|VSS \$273 VINS_BUFF|X 15|25|VSS sg13_lv_nmos L=0.13u W=11.84u
+ AS=2.3606p AD=2.2496p PS=18.96u PD=17.92u
M$249 15|25|VSS A|X$1 \$273 15|25|VSS sg13_lv_nmos L=0.13u W=4.44u AS=0.8436p
+ AD=0.9546p PS=6.72u PD=7.76u
M$255 15|25|VSS \$274 17|NOC_N_BUFF|X 15|25|VSS sg13_lv_nmos L=0.13u W=11.84u
+ AS=2.3606p AD=2.2496p PS=18.96u PD=17.92u
M$271 15|25|VSS A|X$2 \$274 15|25|VSS sg13_lv_nmos L=0.13u W=4.44u AS=0.8436p
+ AD=0.9546p PS=6.72u PD=7.76u
M$277 15|25|VSS \$277 14|VINR_BUFF|X 15|25|VSS sg13_lv_nmos L=0.13u W=11.84u
+ AS=2.3606p AD=2.2496p PS=18.96u PD=17.92u
M$293 15|25|VSS A|X$4 \$277 15|25|VSS sg13_lv_nmos L=0.13u W=4.44u AS=0.8436p
+ AD=0.9546p PS=6.72u PD=7.76u
M$299 15|25|VSS \$275 A|X 15|25|VSS sg13_lv_nmos L=0.13u W=11.84u AS=2.3606p
+ AD=2.2496p PS=18.96u PD=17.92u
M$315 15|25|VSS A|X$3 \$275 15|25|VSS sg13_lv_nmos L=0.13u W=4.44u AS=0.8436p
+ AD=0.9546p PS=6.72u PD=7.76u
M$321 15|25|VSS \$278 A|X$3 15|25|VSS sg13_lv_nmos L=0.13u W=2.96u AS=0.6734p
+ AD=0.7252p PS=5.52u PD=4.92u
M$325 15|25|VSS A$2 \$278 15|25|VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.3034p
+ AD=0.2664p PS=1.56u PD=2.2u
M$326 15|25|VSS A|Y$2 A|B|Y 15|25|VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.259p
+ AD=0.259p PS=2.18u PD=2.18u
M$327 15|25|VSS \$279 A|X$1 15|25|VSS sg13_lv_nmos L=0.13u W=11.84u AS=2.3606p
+ AD=2.2496p PS=18.96u PD=17.92u
M$343 15|25|VSS A|X$5 \$279 15|25|VSS sg13_lv_nmos L=0.13u W=4.44u AS=0.8436p
+ AD=0.9546p PS=6.72u PD=7.76u
M$349 15|25|VSS \$289 14|VINR_BUFF|X 15|25|VSS sg13_lv_nmos L=0.13u W=11.84u
+ AS=2.3606p AD=2.2496p PS=18.96u PD=17.92u
M$365 15|25|VSS A|X$4 \$289 15|25|VSS sg13_lv_nmos L=0.13u W=4.44u AS=0.8436p
+ AD=0.9546p PS=6.72u PD=7.76u
M$371 15|25|VSS \$290 A|X$4 15|25|VSS sg13_lv_nmos L=0.13u W=11.84u AS=2.3606p
+ AD=2.2496p PS=18.96u PD=17.92u
M$387 15|25|VSS A|X$6 \$290 15|25|VSS sg13_lv_nmos L=0.13u W=4.44u AS=0.8436p
+ AD=0.9546p PS=6.72u PD=7.76u
M$393 15|25|VSS \$292 A|X$6 15|25|VSS sg13_lv_nmos L=0.13u W=2.96u AS=0.6734p
+ AD=0.7252p PS=5.52u PD=4.92u
M$397 15|25|VSS A$3 \$292 15|25|VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.3034p
+ AD=0.2664p PS=1.56u PD=2.2u
M$398 \$280 A|B|Y$1 15|25|VSS 15|25|VSS sg13_lv_nmos L=0.13u W=0.55u
+ AS=0.247625p AD=0.159375p PS=2.29u PD=1.19u
M$399 15|25|VSS \$280 A$2 15|25|VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.159375p
+ AD=0.2516p PS=1.19u PD=2.16u
M$400 \$297 A|X$10 15|25|VSS 15|25|VSS sg13_lv_nmos L=0.13u W=0.42u AS=0.1428p
+ AD=0.0798p PS=1.52u PD=0.8u
M$401 15|25|VSS \$297 \$298 15|25|VSS sg13_lv_nmos L=0.5u W=0.42u AS=0.0798p
+ AD=0.1428p PS=0.8u PD=1.52u
M$402 \$282 A|VINR|X 15|25|VSS 15|25|VSS sg13_lv_nmos L=0.13u W=0.55u
+ AS=0.247625p AD=0.159375p PS=2.29u PD=1.19u
M$403 15|25|VSS \$282 A$3 15|25|VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.159375p
+ AD=0.2516p PS=1.19u PD=2.16u
M$404 15|25|VSS \$298 \$299 15|25|VSS sg13_lv_nmos L=0.5u W=0.42u AS=0.1426p
+ AD=0.1428p PS=1.16u PD=1.52u
M$405 15|25|VSS \$299 A|X$8 15|25|VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.1426p
+ AD=0.2516p PS=1.16u PD=2.16u
M$406 15|25|VSS A|VINR|X A|Y$2 15|25|VSS sg13_lv_nmos L=0.13u W=1.48u
+ AS=0.3922p AD=0.3959p PS=3.28u PD=3.29u
M$408 15|25|VSS A|B|Y$2 A|Y$3 15|25|VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.259p
+ AD=0.259p PS=2.18u PD=2.18u
M$409 15|25|VSS A|X$11 A|B|Y$2 15|25|VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.259p
+ AD=0.259p PS=2.18u PD=2.18u
M$410 15|25|VSS \$294 A|X$5 15|25|VSS sg13_lv_nmos L=0.13u W=2.96u AS=0.6734p
+ AD=0.7252p PS=5.52u PD=4.92u
M$414 15|25|VSS A$4 \$294 15|25|VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.3034p
+ AD=0.2664p PS=1.56u PD=2.2u
M$415 15|25|VSS \$295 A|X$2 15|25|VSS sg13_lv_nmos L=0.13u W=11.84u AS=2.3606p
+ AD=2.2496p PS=18.96u PD=17.92u
M$431 15|25|VSS A|X$7 \$295 15|25|VSS sg13_lv_nmos L=0.13u W=4.44u AS=0.8436p
+ AD=0.9546p PS=6.72u PD=7.76u
M$437 15|25|VSS \$312 14|VINR_BUFF|X 15|25|VSS sg13_lv_nmos L=0.13u W=11.84u
+ AS=2.3606p AD=2.2496p PS=18.96u PD=17.92u
M$453 15|25|VSS A|X$4 \$312 15|25|VSS sg13_lv_nmos L=0.13u W=4.44u AS=0.8436p
+ AD=0.9546p PS=6.72u PD=7.76u
M$459 15|25|VSS \$332 14|VINR_BUFF|X 15|25|VSS sg13_lv_nmos L=0.13u W=11.84u
+ AS=2.3606p AD=2.2496p PS=18.96u PD=17.92u
M$475 15|25|VSS A|X$4 \$332 15|25|VSS sg13_lv_nmos L=0.13u W=4.44u AS=0.8436p
+ AD=0.9546p PS=6.72u PD=7.76u
M$481 \$313 A|Y$4 15|25|VSS 15|25|VSS sg13_lv_nmos L=0.13u W=0.42u AS=0.1428p
+ AD=0.0798p PS=1.52u PD=0.8u
M$482 15|25|VSS \$313 \$314 15|25|VSS sg13_lv_nmos L=0.5u W=0.42u AS=0.0798p
+ AD=0.1428p PS=0.8u PD=1.52u
M$483 \$326 \$314 15|25|VSS 15|25|VSS sg13_lv_nmos L=0.5u W=0.42u AS=0.1428p
+ AD=0.1426p PS=1.52u PD=1.16u
M$484 15|25|VSS \$326 A|X$12 15|25|VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.1426p
+ AD=0.2516p PS=1.16u PD=2.16u
M$485 15|25|VSS A|B|Y A|Y$4 15|25|VSS sg13_lv_nmos L=0.13u W=5.92u AS=1.2395p
+ AD=1.2395p PS=10.01u PD=10.01u
M$493 \$334 A|X$12 15|25|VSS 15|25|VSS sg13_lv_nmos L=0.13u W=0.42u AS=0.1428p
+ AD=0.0798p PS=1.52u PD=0.8u
M$494 15|25|VSS \$334 \$335 15|25|VSS sg13_lv_nmos L=0.5u W=0.42u AS=0.0798p
+ AD=0.1428p PS=0.8u PD=1.52u
M$495 15|25|VSS \$335 \$336 15|25|VSS sg13_lv_nmos L=0.5u W=0.42u AS=0.1426p
+ AD=0.1428p PS=1.16u PD=1.52u
M$496 15|25|VSS \$336 A|X$10 15|25|VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.1426p
+ AD=0.2516p PS=1.16u PD=2.16u
M$497 \$317 A|X$8 15|25|VSS 15|25|VSS sg13_lv_nmos L=0.13u W=0.42u AS=0.1428p
+ AD=0.0798p PS=1.52u PD=0.8u
M$498 15|25|VSS \$317 \$318 15|25|VSS sg13_lv_nmos L=0.5u W=0.42u AS=0.0798p
+ AD=0.1428p PS=0.8u PD=1.52u
M$499 \$327 \$318 15|25|VSS 15|25|VSS sg13_lv_nmos L=0.5u W=0.42u AS=0.1428p
+ AD=0.1426p PS=1.52u PD=1.16u
M$500 15|25|VSS \$327 A|X$13 15|25|VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.1426p
+ AD=0.2516p PS=1.16u PD=2.16u
M$501 15|25|VSS A|Y$9 A|B|Y$1 15|25|VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.2516p
+ AD=0.1406p PS=2.16u PD=1.12u
M$502 A|B|Y$1 B|X 15|25|VSS 15|25|VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.1406p
+ AD=0.2516p PS=1.12u PD=2.16u
M$503 \$303 A|Y$3 \$309 15|25|VSS sg13_lv_nmos L=0.13u W=0.64u AS=0.2176p
+ AD=0.1216p PS=1.96u PD=1.02u
M$504 15|25|VSS A|B|Y \$309 15|25|VSS sg13_lv_nmos L=0.13u W=0.64u AS=0.1331p
+ AD=0.1216p PS=1.12u PD=1.02u
M$505 15|25|VSS \$303 A|X$9 15|25|VSS sg13_lv_nmos L=0.13u W=1.48u AS=0.2737p
+ AD=0.4218p PS=2.24u PD=3.36u
M$507 \$320 A|X$13 15|25|VSS 15|25|VSS sg13_lv_nmos L=0.13u W=0.42u AS=0.1428p
+ AD=0.0798p PS=1.52u PD=0.8u
M$508 15|25|VSS \$320 \$321 15|25|VSS sg13_lv_nmos L=0.5u W=0.42u AS=0.0798p
+ AD=0.1428p PS=0.8u PD=1.52u
M$509 15|25|VSS A|X$9 A|Y$9 15|25|VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.2516p
+ AD=0.1406p PS=2.16u PD=1.12u
M$510 A|Y$9 A|B|Y$1 15|25|VSS 15|25|VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.1406p
+ AD=0.2516p PS=1.12u PD=2.16u
M$511 \$328 \$321 15|25|VSS 15|25|VSS sg13_lv_nmos L=0.5u W=0.42u AS=0.1428p
+ AD=0.1426p PS=1.52u PD=1.16u
M$512 15|25|VSS \$328 A|X$11 15|25|VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.1426p
+ AD=0.2516p PS=1.16u PD=2.16u
M$513 15|25|VSS A|B|Y A|Y$5 15|25|VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.259p
+ AD=0.259p PS=2.18u PD=2.18u
M$514 15|25|VSS A|B|Y$3 A|Y$6 15|25|VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.259p
+ AD=0.259p PS=2.18u PD=2.18u
M$515 15|25|VSS A|B|Y$4 A|Y$7 15|25|VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.259p
+ AD=0.259p PS=2.18u PD=2.18u
M$516 15|25|VSS A|Y$8 A|B|Y$3 15|25|VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.259p
+ AD=0.259p PS=2.18u PD=2.18u
M$517 15|25|VSS A|VINS|X A|Y$8 15|25|VSS sg13_lv_nmos L=0.13u W=1.48u
+ AS=0.3922p AD=0.3959p PS=3.28u PD=3.29u
M$519 \$325 A|VINS|X 15|25|VSS 15|25|VSS sg13_lv_nmos L=0.13u W=0.55u
+ AS=0.247625p AD=0.159375p PS=2.29u PD=1.19u
M$520 15|25|VSS \$325 A$4 15|25|VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.159375p
+ AD=0.2516p PS=1.19u PD=2.16u
M$521 15|25|VSS \$333 A|X$7 15|25|VSS sg13_lv_nmos L=0.13u W=2.96u AS=0.6734p
+ AD=0.7252p PS=5.52u PD=4.92u
M$525 15|25|VSS A$5 \$333 15|25|VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.3034p
+ AD=0.2664p PS=1.56u PD=2.2u
M$526 15|25|VSS \$349 18|NOC_P_BUFF|X 15|25|VSS sg13_lv_nmos L=0.13u W=11.84u
+ AS=2.3606p AD=2.2496p PS=18.96u PD=17.92u
M$542 15|25|VSS A|X$14 \$349 15|25|VSS sg13_lv_nmos L=0.13u W=4.44u AS=0.8436p
+ AD=0.9546p PS=6.72u PD=7.76u
M$548 \$338 A|Y$5 \$346 15|25|VSS sg13_lv_nmos L=0.13u W=0.64u AS=0.2176p
+ AD=0.1216p PS=1.96u PD=1.02u
M$549 15|25|VSS A|B|Y$2 \$346 15|25|VSS sg13_lv_nmos L=0.13u W=0.64u AS=0.1331p
+ AD=0.1216p PS=1.12u PD=1.02u
M$550 15|25|VSS \$338 X 15|25|VSS sg13_lv_nmos L=0.13u W=1.48u AS=0.2737p
+ AD=0.4218p PS=2.24u PD=3.36u
M$552 15|25|VSS A|B|Y$3 A|Y$10 15|25|VSS sg13_lv_nmos L=0.13u W=5.92u
+ AS=1.2395p AD=1.2395p PS=10.01u PD=10.01u
M$560 \$340 A|Y$7 \$345 15|25|VSS sg13_lv_nmos L=0.13u W=0.64u AS=0.2176p
+ AD=0.1216p PS=1.96u PD=1.02u
M$561 15|25|VSS A|B|Y$3 \$345 15|25|VSS sg13_lv_nmos L=0.13u W=0.64u AS=0.1331p
+ AD=0.1216p PS=1.12u PD=1.02u
M$562 15|25|VSS \$340 B|X 15|25|VSS sg13_lv_nmos L=0.13u W=1.48u AS=0.2737p
+ AD=0.4218p PS=2.24u PD=3.36u
M$564 \$341 A|Y$6 \$344 15|25|VSS sg13_lv_nmos L=0.13u W=0.64u AS=0.2176p
+ AD=0.1216p PS=1.96u PD=1.02u
M$565 15|25|VSS A|B|Y$4 \$344 15|25|VSS sg13_lv_nmos L=0.13u W=0.64u AS=0.1331p
+ AD=0.1216p PS=1.12u PD=1.02u
M$566 15|25|VSS \$341 X 15|25|VSS sg13_lv_nmos L=0.13u W=1.48u AS=0.2737p
+ AD=0.4218p PS=2.24u PD=3.36u
M$568 15|25|VSS A|X$15 A|B|Y$4 15|25|VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.259p
+ AD=0.259p PS=2.18u PD=2.18u
M$569 \$354 \$353 15|25|VSS 15|25|VSS sg13_lv_nmos L=0.5u W=0.42u AS=0.1428p
+ AD=0.1426p PS=1.52u PD=1.16u
M$570 15|25|VSS \$354 A|X$15 15|25|VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.1426p
+ AD=0.2516p PS=1.16u PD=2.16u
M$571 15|25|VSS \$358 18|NOC_P_BUFF|X 15|25|VSS sg13_lv_nmos L=0.13u W=11.84u
+ AS=2.3606p AD=2.2496p PS=18.96u PD=17.92u
M$587 15|25|VSS A|X$14 \$358 15|25|VSS sg13_lv_nmos L=0.13u W=4.44u AS=0.8436p
+ AD=0.9546p PS=6.72u PD=7.76u
M$593 \$359 A|Y$10 15|25|VSS 15|25|VSS sg13_lv_nmos L=0.13u W=0.42u AS=0.1428p
+ AD=0.0798p PS=1.52u PD=0.8u
M$594 15|25|VSS \$359 \$360 15|25|VSS sg13_lv_nmos L=0.5u W=0.42u AS=0.0798p
+ AD=0.1428p PS=0.8u PD=1.52u
M$595 15|25|VSS \$360 \$368 15|25|VSS sg13_lv_nmos L=0.5u W=0.42u AS=0.1426p
+ AD=0.1428p PS=1.16u PD=1.52u
M$596 15|25|VSS \$368 A|X$17 15|25|VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.1426p
+ AD=0.2516p PS=1.16u PD=2.16u
M$597 \$362 A|X$17 15|25|VSS 15|25|VSS sg13_lv_nmos L=0.13u W=0.42u AS=0.1428p
+ AD=0.0798p PS=1.52u PD=0.8u
M$598 15|25|VSS \$362 \$363 15|25|VSS sg13_lv_nmos L=0.5u W=0.42u AS=0.0798p
+ AD=0.1428p PS=0.8u PD=1.52u
M$599 \$352 A|X$16 15|25|VSS 15|25|VSS sg13_lv_nmos L=0.13u W=0.42u AS=0.1428p
+ AD=0.0798p PS=1.52u PD=0.8u
M$600 15|25|VSS \$352 \$353 15|25|VSS sg13_lv_nmos L=0.5u W=0.42u AS=0.0798p
+ AD=0.1428p PS=0.8u PD=1.52u
M$601 15|25|VSS \$363 \$369 15|25|VSS sg13_lv_nmos L=0.5u W=0.42u AS=0.1426p
+ AD=0.1428p PS=1.16u PD=1.52u
M$602 15|25|VSS \$369 A|X$18 15|25|VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.1426p
+ AD=0.2516p PS=1.16u PD=2.16u
M$603 \$365 A|X$18 15|25|VSS 15|25|VSS sg13_lv_nmos L=0.13u W=0.42u AS=0.1428p
+ AD=0.0798p PS=1.52u PD=0.8u
M$604 15|25|VSS \$365 \$366 15|25|VSS sg13_lv_nmos L=0.5u W=0.42u AS=0.0798p
+ AD=0.1428p PS=0.8u PD=1.52u
M$605 15|25|VSS \$366 \$370 15|25|VSS sg13_lv_nmos L=0.5u W=0.42u AS=0.1426p
+ AD=0.1428p PS=1.16u PD=1.52u
M$606 15|25|VSS \$370 A|X$19 15|25|VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.1426p
+ AD=0.2516p PS=1.16u PD=2.16u
M$607 \$351 NOC_N|X 15|25|VSS 15|25|VSS sg13_lv_nmos L=0.13u W=0.55u
+ AS=0.247625p AD=0.159375p PS=2.29u PD=1.19u
M$608 15|25|VSS \$351 A$5 15|25|VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.159375p
+ AD=0.2516p PS=1.19u PD=2.16u
M$609 15|25|VSS \$381 18|NOC_P_BUFF|X 15|25|VSS sg13_lv_nmos L=0.13u W=11.84u
+ AS=2.3606p AD=2.2496p PS=18.96u PD=17.92u
M$625 15|25|VSS A|X$14 \$381 15|25|VSS sg13_lv_nmos L=0.13u W=4.44u AS=0.8436p
+ AD=0.9546p PS=6.72u PD=7.76u
M$631 15|25|VSS \$372 18|NOC_P_BUFF|X 15|25|VSS sg13_lv_nmos L=0.13u W=11.84u
+ AS=2.3606p AD=2.2496p PS=18.96u PD=17.92u
M$647 15|25|VSS A|X$14 \$372 15|25|VSS sg13_lv_nmos L=0.13u W=4.44u AS=0.8436p
+ AD=0.9546p PS=6.72u PD=7.76u
M$653 15|25|VSS \$382 A|X$14 15|25|VSS sg13_lv_nmos L=0.13u W=11.84u AS=2.3606p
+ AD=2.2496p PS=18.96u PD=17.92u
M$669 15|25|VSS A|X$20 \$382 15|25|VSS sg13_lv_nmos L=0.13u W=4.44u AS=0.8436p
+ AD=0.9546p PS=6.72u PD=7.76u
M$675 15|25|VSS \$384 A|X$20 15|25|VSS sg13_lv_nmos L=0.13u W=2.96u AS=0.6734p
+ AD=0.7252p PS=5.52u PD=4.92u
M$679 15|25|VSS A$6 \$384 15|25|VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.3034p
+ AD=0.2664p PS=1.56u PD=2.2u
M$680 \$385 A|X$25 15|25|VSS 15|25|VSS sg13_lv_nmos L=0.13u W=0.42u AS=0.1428p
+ AD=0.0798p PS=1.52u PD=0.8u
M$681 15|25|VSS \$385 \$386 15|25|VSS sg13_lv_nmos L=0.5u W=0.42u AS=0.0798p
+ AD=0.1428p PS=0.8u PD=1.52u
M$682 15|25|VSS \$386 \$387 15|25|VSS sg13_lv_nmos L=0.5u W=0.42u AS=0.1426p
+ AD=0.1428p PS=1.16u PD=1.52u
M$683 15|25|VSS \$387 A|X$21 15|25|VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.1426p
+ AD=0.2516p PS=1.16u PD=2.16u
M$684 \$389 A|X$21 15|25|VSS 15|25|VSS sg13_lv_nmos L=0.13u W=0.42u AS=0.1428p
+ AD=0.0798p PS=1.52u PD=0.8u
M$685 15|25|VSS \$389 \$390 15|25|VSS sg13_lv_nmos L=0.5u W=0.42u AS=0.0798p
+ AD=0.1428p PS=0.8u PD=1.52u
M$686 15|25|VSS \$390 \$391 15|25|VSS sg13_lv_nmos L=0.5u W=0.42u AS=0.1426p
+ AD=0.1428p PS=1.16u PD=1.52u
M$687 15|25|VSS \$391 A|X$22 15|25|VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.1426p
+ AD=0.2516p PS=1.16u PD=2.16u
M$688 \$393 A|X$22 15|25|VSS 15|25|VSS sg13_lv_nmos L=0.13u W=0.42u AS=0.1428p
+ AD=0.0798p PS=1.52u PD=0.8u
M$689 15|25|VSS \$393 \$394 15|25|VSS sg13_lv_nmos L=0.5u W=0.42u AS=0.0798p
+ AD=0.1428p PS=0.8u PD=1.52u
M$690 15|25|VSS \$394 \$395 15|25|VSS sg13_lv_nmos L=0.5u W=0.42u AS=0.1426p
+ AD=0.1428p PS=1.16u PD=1.52u
M$691 15|25|VSS \$395 A|X$23 15|25|VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.1426p
+ AD=0.2516p PS=1.16u PD=2.16u
M$692 \$397 A|X$23 15|25|VSS 15|25|VSS sg13_lv_nmos L=0.13u W=0.42u AS=0.1428p
+ AD=0.0798p PS=1.52u PD=0.8u
M$693 15|25|VSS \$397 \$398 15|25|VSS sg13_lv_nmos L=0.5u W=0.42u AS=0.0798p
+ AD=0.1428p PS=0.8u PD=1.52u
M$694 \$375 A|X$19 15|25|VSS 15|25|VSS sg13_lv_nmos L=0.13u W=0.42u AS=0.1428p
+ AD=0.0798p PS=1.52u PD=0.8u
M$695 15|25|VSS \$375 \$376 15|25|VSS sg13_lv_nmos L=0.5u W=0.42u AS=0.0798p
+ AD=0.1428p PS=0.8u PD=1.52u
M$696 15|25|VSS \$398 \$399 15|25|VSS sg13_lv_nmos L=0.5u W=0.42u AS=0.1426p
+ AD=0.1428p PS=1.16u PD=1.52u
M$697 15|25|VSS \$399 A|X$24 15|25|VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.1426p
+ AD=0.2516p PS=1.16u PD=2.16u
M$698 \$379 \$376 15|25|VSS 15|25|VSS sg13_lv_nmos L=0.5u W=0.42u AS=0.1428p
+ AD=0.1426p PS=1.52u PD=1.16u
M$699 15|25|VSS \$379 A|X$16 15|25|VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.1426p
+ AD=0.2516p PS=1.16u PD=2.16u
M$700 \$416 A|X$28 15|25|VSS 15|25|VSS sg13_lv_nmos L=0.13u W=0.42u AS=0.1428p
+ AD=0.0798p PS=1.52u PD=0.8u
M$701 15|25|VSS \$416 \$418 15|25|VSS sg13_lv_nmos L=0.5u W=0.42u AS=0.0798p
+ AD=0.1428p PS=0.8u PD=1.52u
M$702 15|25|VSS \$418 \$419 15|25|VSS sg13_lv_nmos L=0.5u W=0.42u AS=0.1426p
+ AD=0.1428p PS=1.16u PD=1.52u
M$703 15|25|VSS \$419 A|X$29 15|25|VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.1426p
+ AD=0.2516p PS=1.16u PD=2.16u
M$704 \$421 A|Y$12 15|25|VSS 15|25|VSS sg13_lv_nmos L=0.13u W=0.42u AS=0.1428p
+ AD=0.0798p PS=1.52u PD=0.8u
M$705 15|25|VSS \$421 \$423 15|25|VSS sg13_lv_nmos L=0.5u W=0.42u AS=0.0798p
+ AD=0.1428p PS=0.8u PD=1.52u
M$706 15|25|VSS \$423 \$424 15|25|VSS sg13_lv_nmos L=0.5u W=0.42u AS=0.1426p
+ AD=0.1428p PS=1.16u PD=1.52u
M$707 15|25|VSS \$424 A|X$30 15|25|VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.1426p
+ AD=0.2516p PS=1.16u PD=2.16u
M$708 \$426 A|X$31 15|25|VSS 15|25|VSS sg13_lv_nmos L=0.13u W=0.42u AS=0.1428p
+ AD=0.0798p PS=1.52u PD=0.8u
M$709 15|25|VSS \$426 \$428 15|25|VSS sg13_lv_nmos L=0.5u W=0.42u AS=0.0798p
+ AD=0.1428p PS=0.8u PD=1.52u
M$710 15|25|VSS \$428 \$429 15|25|VSS sg13_lv_nmos L=0.5u W=0.42u AS=0.1426p
+ AD=0.1428p PS=1.16u PD=1.52u
M$711 15|25|VSS \$429 A|X$32 15|25|VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.1426p
+ AD=0.2516p PS=1.16u PD=2.16u
M$712 \$431 A|X$33 15|25|VSS 15|25|VSS sg13_lv_nmos L=0.13u W=0.42u AS=0.1428p
+ AD=0.0798p PS=1.52u PD=0.8u
M$713 15|25|VSS \$431 \$433 15|25|VSS sg13_lv_nmos L=0.5u W=0.42u AS=0.0798p
+ AD=0.1428p PS=0.8u PD=1.52u
M$714 15|25|VSS \$433 \$434 15|25|VSS sg13_lv_nmos L=0.5u W=0.42u AS=0.1426p
+ AD=0.1428p PS=1.16u PD=1.52u
M$715 15|25|VSS \$434 A|X$34 15|25|VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.1426p
+ AD=0.2516p PS=1.16u PD=2.16u
M$716 \$436 A|Y$11 15|25|VSS 15|25|VSS sg13_lv_nmos L=0.13u W=0.42u AS=0.1428p
+ AD=0.0798p PS=1.52u PD=0.8u
M$717 15|25|VSS \$436 \$437 15|25|VSS sg13_lv_nmos L=0.5u W=0.42u AS=0.0798p
+ AD=0.1428p PS=0.8u PD=1.52u
M$718 15|25|VSS \$437 \$438 15|25|VSS sg13_lv_nmos L=0.5u W=0.42u AS=0.1426p
+ AD=0.1428p PS=1.16u PD=1.52u
M$719 15|25|VSS \$438 A|X$35 15|25|VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.1426p
+ AD=0.2516p PS=1.16u PD=2.16u
M$720 \$403 A|Y$11 15|25|VSS 15|25|VSS sg13_lv_nmos L=0.13u W=0.42u AS=0.1428p
+ AD=0.0798p PS=1.52u PD=0.8u
M$721 15|25|VSS \$403 \$404 15|25|VSS sg13_lv_nmos L=0.5u W=0.42u AS=0.0798p
+ AD=0.1428p PS=0.8u PD=1.52u
M$722 \$411 \$404 15|25|VSS 15|25|VSS sg13_lv_nmos L=0.5u W=0.42u AS=0.1428p
+ AD=0.1426p PS=1.52u PD=1.16u
M$723 15|25|VSS \$411 A|X$25 15|25|VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.1426p
+ AD=0.2516p PS=1.16u PD=2.16u
M$724 15|25|VSS A|X$36 A|Y$11 15|25|VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.2516p
+ AD=0.1406p PS=2.16u PD=1.12u
M$725 A|Y$11 A|B|Y$1 15|25|VSS 15|25|VSS sg13_lv_nmos L=0.13u W=0.74u
+ AS=0.1406p AD=0.2516p PS=1.12u PD=2.16u
M$726 15|25|VSS A|X$36 A|Y$13 15|25|VSS sg13_lv_nmos L=0.13u W=1.48u AS=0.3922p
+ AD=0.3959p PS=3.28u PD=3.29u
M$728 15|25|VSS A|Y$14 A|Y$12 15|25|VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.2516p
+ AD=0.1406p PS=2.16u PD=1.12u
M$729 A|Y$12 A|B|X 15|25|VSS 15|25|VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.1406p
+ AD=0.2516p PS=1.12u PD=2.16u
M$730 15|25|VSS A|B|Y$1 A|Y$14 15|25|VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.259p
+ AD=0.259p PS=2.18u PD=2.18u
M$731 15|25|VSS NOC_P|X \$444 15|25|VSS sg13_lv_nmos L=0.13u W=0.55u
+ AS=0.159375p AD=0.247625p PS=1.19u PD=2.29u
M$732 15|25|VSS \$444 A$6 15|25|VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.159375p
+ AD=0.2516p PS=1.19u PD=2.16u
M$733 15|25|VSS A|Y$15 A0|Y 15|25|VSS sg13_lv_nmos L=0.13u W=2.96u AS=0.6734p
+ AD=0.6734p PS=5.52u PD=5.52u
M$737 15|25|VSS A|B|X A|Y$16 15|25|VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.259p
+ AD=0.259p PS=2.18u PD=2.18u
M$738 \$405 A|X$24 15|25|VSS 15|25|VSS sg13_lv_nmos L=0.13u W=0.42u AS=0.1428p
+ AD=0.0798p PS=1.52u PD=0.8u
M$739 15|25|VSS \$405 \$406 15|25|VSS sg13_lv_nmos L=0.5u W=0.42u AS=0.0798p
+ AD=0.1428p PS=0.8u PD=1.52u
M$740 \$412 \$406 15|25|VSS 15|25|VSS sg13_lv_nmos L=0.5u W=0.42u AS=0.1428p
+ AD=0.1426p PS=1.52u PD=1.16u
M$741 15|25|VSS \$412 A|X$26 15|25|VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.1426p
+ AD=0.2516p PS=1.16u PD=2.16u
M$742 \$447 A|X$27 15|25|VSS 15|25|VSS sg13_lv_nmos L=0.13u W=0.42u AS=0.1428p
+ AD=0.0798p PS=1.52u PD=0.8u
M$743 15|25|VSS \$447 \$448 15|25|VSS sg13_lv_nmos L=0.5u W=0.42u AS=0.0798p
+ AD=0.1428p PS=0.8u PD=1.52u
M$744 \$408 A|X$26 15|25|VSS 15|25|VSS sg13_lv_nmos L=0.13u W=0.42u AS=0.1428p
+ AD=0.0798p PS=1.52u PD=0.8u
M$745 15|25|VSS \$408 \$409 15|25|VSS sg13_lv_nmos L=0.5u W=0.42u AS=0.0798p
+ AD=0.1428p PS=0.8u PD=1.52u
M$746 \$413 \$409 15|25|VSS 15|25|VSS sg13_lv_nmos L=0.5u W=0.42u AS=0.1428p
+ AD=0.1426p PS=1.52u PD=1.16u
M$747 15|25|VSS \$413 A|X$27 15|25|VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.1426p
+ AD=0.2516p PS=1.16u PD=2.16u
M$748 15|25|VSS \$448 \$449 15|25|VSS sg13_lv_nmos L=0.5u W=0.42u AS=0.1426p
+ AD=0.1428p PS=1.16u PD=1.52u
M$749 15|25|VSS \$449 A|X$37 15|25|VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.1426p
+ AD=0.2516p PS=1.16u PD=2.16u
M$750 \$451 A|X$37 15|25|VSS 15|25|VSS sg13_lv_nmos L=0.13u W=0.42u AS=0.1428p
+ AD=0.0798p PS=1.52u PD=0.8u
M$751 15|25|VSS \$451 \$452 15|25|VSS sg13_lv_nmos L=0.5u W=0.42u AS=0.0798p
+ AD=0.1428p PS=0.8u PD=1.52u
M$752 15|25|VSS \$452 \$453 15|25|VSS sg13_lv_nmos L=0.5u W=0.42u AS=0.1426p
+ AD=0.1428p PS=1.16u PD=1.52u
M$753 15|25|VSS \$453 A|X$38 15|25|VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.1426p
+ AD=0.2516p PS=1.16u PD=2.16u
M$754 \$458 A|Y$12 15|25|VSS 15|25|VSS sg13_lv_nmos L=0.13u W=0.42u AS=0.1428p
+ AD=0.0798p PS=1.52u PD=0.8u
M$755 15|25|VSS \$458 \$459 15|25|VSS sg13_lv_nmos L=0.5u W=0.42u AS=0.0798p
+ AD=0.1428p PS=0.8u PD=1.52u
M$756 \$490 \$459 15|25|VSS 15|25|VSS sg13_lv_nmos L=0.5u W=0.42u AS=0.1428p
+ AD=0.1426p PS=1.52u PD=1.16u
M$757 15|25|VSS \$490 A|X$39 15|25|VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.1426p
+ AD=0.2516p PS=1.16u PD=2.16u
M$758 \$461 A|X$46 15|25|VSS 15|25|VSS sg13_lv_nmos L=0.13u W=0.42u AS=0.1428p
+ AD=0.0798p PS=1.52u PD=0.8u
M$759 15|25|VSS \$461 \$462 15|25|VSS sg13_lv_nmos L=0.5u W=0.42u AS=0.0798p
+ AD=0.1428p PS=0.8u PD=1.52u
M$760 \$492 \$462 15|25|VSS 15|25|VSS sg13_lv_nmos L=0.5u W=0.42u AS=0.1428p
+ AD=0.1426p PS=1.52u PD=1.16u
M$761 15|25|VSS \$492 A|X$40 15|25|VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.1426p
+ AD=0.2516p PS=1.16u PD=2.16u
M$762 \$464 A|X$30 15|25|VSS 15|25|VSS sg13_lv_nmos L=0.13u W=0.42u AS=0.1428p
+ AD=0.0798p PS=1.52u PD=0.8u
M$763 15|25|VSS \$464 \$465 15|25|VSS sg13_lv_nmos L=0.5u W=0.42u AS=0.0798p
+ AD=0.1428p PS=0.8u PD=1.52u
M$764 \$493 \$465 15|25|VSS 15|25|VSS sg13_lv_nmos L=0.5u W=0.42u AS=0.1428p
+ AD=0.1426p PS=1.52u PD=1.16u
M$765 15|25|VSS \$493 A|X$41 15|25|VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.1426p
+ AD=0.2516p PS=1.16u PD=2.16u
M$766 \$467 A|X$32 15|25|VSS 15|25|VSS sg13_lv_nmos L=0.13u W=0.42u AS=0.1428p
+ AD=0.0798p PS=1.52u PD=0.8u
M$767 15|25|VSS \$467 \$468 15|25|VSS sg13_lv_nmos L=0.5u W=0.42u AS=0.0798p
+ AD=0.1428p PS=0.8u PD=1.52u
M$768 \$494 \$468 15|25|VSS 15|25|VSS sg13_lv_nmos L=0.5u W=0.42u AS=0.1428p
+ AD=0.1426p PS=1.52u PD=1.16u
M$769 15|25|VSS \$494 A|X$42 15|25|VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.1426p
+ AD=0.2516p PS=1.16u PD=2.16u
M$770 \$470 A|X$42 15|25|VSS 15|25|VSS sg13_lv_nmos L=0.13u W=0.42u AS=0.1428p
+ AD=0.0798p PS=1.52u PD=0.8u
M$771 15|25|VSS \$470 \$471 15|25|VSS sg13_lv_nmos L=0.5u W=0.42u AS=0.0798p
+ AD=0.1428p PS=0.8u PD=1.52u
M$772 \$495 \$471 15|25|VSS 15|25|VSS sg13_lv_nmos L=0.5u W=0.42u AS=0.1428p
+ AD=0.1426p PS=1.52u PD=1.16u
M$773 15|25|VSS \$495 A|X$43 15|25|VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.1426p
+ AD=0.2516p PS=1.16u PD=2.16u
M$774 \$473 A|X$34 15|25|VSS 15|25|VSS sg13_lv_nmos L=0.13u W=0.42u AS=0.1428p
+ AD=0.0798p PS=1.52u PD=0.8u
M$775 15|25|VSS \$473 \$474 15|25|VSS sg13_lv_nmos L=0.5u W=0.42u AS=0.0798p
+ AD=0.1428p PS=0.8u PD=1.52u
M$776 \$496 \$474 15|25|VSS 15|25|VSS sg13_lv_nmos L=0.5u W=0.42u AS=0.1428p
+ AD=0.1426p PS=1.52u PD=1.16u
M$777 15|25|VSS \$496 A0|X 15|25|VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.1426p
+ AD=0.2516p PS=1.16u PD=2.16u
M$778 \$476 A|X$35 15|25|VSS 15|25|VSS sg13_lv_nmos L=0.13u W=0.42u AS=0.1428p
+ AD=0.0798p PS=1.52u PD=0.8u
M$779 15|25|VSS \$476 \$477 15|25|VSS sg13_lv_nmos L=0.5u W=0.42u AS=0.0798p
+ AD=0.1428p PS=0.8u PD=1.52u
M$780 \$497 \$477 15|25|VSS 15|25|VSS sg13_lv_nmos L=0.5u W=0.42u AS=0.1428p
+ AD=0.1426p PS=1.52u PD=1.16u
M$781 15|25|VSS \$497 A|X$44 15|25|VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.1426p
+ AD=0.2516p PS=1.16u PD=2.16u
M$782 \$479 A|X$44 15|25|VSS 15|25|VSS sg13_lv_nmos L=0.13u W=0.42u AS=0.1428p
+ AD=0.0798p PS=1.52u PD=0.8u
M$783 15|25|VSS \$479 \$480 15|25|VSS sg13_lv_nmos L=0.5u W=0.42u AS=0.0798p
+ AD=0.1428p PS=0.8u PD=1.52u
M$784 \$498 \$480 15|25|VSS 15|25|VSS sg13_lv_nmos L=0.5u W=0.42u AS=0.1428p
+ AD=0.1426p PS=1.52u PD=1.16u
M$785 15|25|VSS \$498 A|X$45 15|25|VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.1426p
+ AD=0.2516p PS=1.16u PD=2.16u
M$786 15|25|VSS A|Y$13 A0|Y$1 15|25|VSS sg13_lv_nmos L=0.13u W=2.96u AS=0.6734p
+ AD=0.6734p PS=5.52u PD=5.52u
M$790 \$483 12|S|VSEL_OL 15|25|VSS 15|25|VSS sg13_lv_nmos L=0.13u W=0.55u
+ AS=0.187p AD=0.18945p PS=1.78u PD=1.27u
M$791 15|25|VSS 12|S|VSEL_OL \$508 15|25|VSS sg13_lv_nmos L=0.13u W=0.74u
+ AS=0.18945p AD=0.13135p PS=1.27u PD=1.095u
M$792 \$508 11|A1|VINR_OL \$484 15|25|VSS sg13_lv_nmos L=0.13u W=0.74u
+ AS=0.13135p AD=0.1628p PS=1.095u PD=1.18u
M$793 \$484 A0|Y$1 \$507 15|25|VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.1628p
+ AD=0.3367p PS=1.18u PD=1.65u
M$794 \$507 \$483 15|25|VSS 15|25|VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.3367p
+ AD=0.148p PS=1.65u PD=1.14u
M$795 15|25|VSS \$484 NOC_N|X 15|25|VSS sg13_lv_nmos L=0.13u W=1.48u AS=0.3515p
+ AD=0.518p PS=2.43u PD=3.62u
M$797 \$485 12|S|VSEL_OL 15|25|VSS 15|25|VSS sg13_lv_nmos L=0.13u W=0.55u
+ AS=0.187p AD=0.18945p PS=1.78u PD=1.27u
M$798 15|25|VSS 12|S|VSEL_OL \$506 15|25|VSS sg13_lv_nmos L=0.13u W=0.74u
+ AS=0.18945p AD=0.13135p PS=1.27u PD=1.095u
M$799 \$506 10|A1|VINS_OL \$486 15|25|VSS sg13_lv_nmos L=0.13u W=0.74u
+ AS=0.13135p AD=0.1628p PS=1.095u PD=1.18u
M$800 \$486 A0|Y \$505 15|25|VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.1628p
+ AD=0.3367p PS=1.18u PD=1.65u
M$801 \$505 \$485 15|25|VSS 15|25|VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.3367p
+ AD=0.148p PS=1.65u PD=1.14u
M$802 15|25|VSS \$486 NOC_P|X 15|25|VSS sg13_lv_nmos L=0.13u W=1.48u AS=0.3515p
+ AD=0.518p PS=2.43u PD=3.62u
M$804 \$487 A|X$38 15|25|VSS 15|25|VSS sg13_lv_nmos L=0.13u W=0.42u AS=0.1428p
+ AD=0.0798p PS=1.52u PD=0.8u
M$805 15|25|VSS \$487 \$488 15|25|VSS sg13_lv_nmos L=0.5u W=0.42u AS=0.0798p
+ AD=0.1428p PS=0.8u PD=1.52u
M$806 \$499 \$488 15|25|VSS 15|25|VSS sg13_lv_nmos L=0.5u W=0.42u AS=0.1428p
+ AD=0.1426p PS=1.52u PD=1.16u
M$807 15|25|VSS \$499 A1|X 15|25|VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.1426p
+ AD=0.2516p PS=1.16u PD=2.16u
M$808 \$509 A|X$39 15|25|VSS 15|25|VSS sg13_lv_nmos L=0.13u W=0.42u AS=0.1428p
+ AD=0.0798p PS=1.52u PD=0.8u
M$809 15|25|VSS \$509 \$510 15|25|VSS sg13_lv_nmos L=0.5u W=0.42u AS=0.0798p
+ AD=0.1428p PS=0.8u PD=1.52u
M$810 15|25|VSS \$510 \$511 15|25|VSS sg13_lv_nmos L=0.5u W=0.42u AS=0.1426p
+ AD=0.1428p PS=1.16u PD=1.52u
M$811 15|25|VSS \$511 A|X$28 15|25|VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.1426p
+ AD=0.2516p PS=1.16u PD=2.16u
M$812 \$512 A|X$29 15|25|VSS 15|25|VSS sg13_lv_nmos L=0.13u W=0.42u AS=0.1428p
+ AD=0.0798p PS=1.52u PD=0.8u
M$813 15|25|VSS \$512 \$513 15|25|VSS sg13_lv_nmos L=0.5u W=0.42u AS=0.0798p
+ AD=0.1428p PS=0.8u PD=1.52u
M$814 15|25|VSS \$513 \$514 15|25|VSS sg13_lv_nmos L=0.5u W=0.42u AS=0.1426p
+ AD=0.1428p PS=1.16u PD=1.52u
M$815 15|25|VSS \$514 A|X$46 15|25|VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.1426p
+ AD=0.2516p PS=1.16u PD=2.16u
M$816 \$515 A|X$40 15|25|VSS 15|25|VSS sg13_lv_nmos L=0.13u W=0.42u AS=0.1428p
+ AD=0.0798p PS=1.52u PD=0.8u
M$817 15|25|VSS \$515 \$516 15|25|VSS sg13_lv_nmos L=0.5u W=0.42u AS=0.0798p
+ AD=0.1428p PS=0.8u PD=1.52u
M$818 15|25|VSS \$516 \$517 15|25|VSS sg13_lv_nmos L=0.5u W=0.42u AS=0.1426p
+ AD=0.1428p PS=1.16u PD=1.52u
M$819 15|25|VSS \$517 A|X$31 15|25|VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.1426p
+ AD=0.2516p PS=1.16u PD=2.16u
M$820 \$518 A|X$41 15|25|VSS 15|25|VSS sg13_lv_nmos L=0.13u W=0.42u AS=0.1428p
+ AD=0.0798p PS=1.52u PD=0.8u
M$821 15|25|VSS \$518 \$519 15|25|VSS sg13_lv_nmos L=0.5u W=0.42u AS=0.0798p
+ AD=0.1428p PS=0.8u PD=1.52u
M$822 15|25|VSS \$519 \$520 15|25|VSS sg13_lv_nmos L=0.5u W=0.42u AS=0.1426p
+ AD=0.1428p PS=1.16u PD=1.52u
M$823 15|25|VSS \$520 A|X$33 15|25|VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.1426p
+ AD=0.2516p PS=1.16u PD=2.16u
M$824 \$521 A|X$43 15|25|VSS 15|25|VSS sg13_lv_nmos L=0.13u W=0.42u AS=0.1428p
+ AD=0.0798p PS=1.52u PD=0.8u
M$825 15|25|VSS \$521 \$522 15|25|VSS sg13_lv_nmos L=0.5u W=0.42u AS=0.0798p
+ AD=0.1428p PS=0.8u PD=1.52u
M$826 15|25|VSS \$522 \$523 15|25|VSS sg13_lv_nmos L=0.5u W=0.42u AS=0.1426p
+ AD=0.1428p PS=1.16u PD=1.52u
M$827 15|25|VSS \$523 A1|X$1 15|25|VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.1426p
+ AD=0.2516p PS=1.16u PD=2.16u
M$828 15|25|VSS 13|S|VSEL_DT \$525 15|25|VSS sg13_lv_nmos L=0.13u W=0.55u
+ AS=0.18945p AD=0.187p PS=1.27u PD=1.78u
M$829 15|25|VSS 13|S|VSEL_DT \$537 15|25|VSS sg13_lv_nmos L=0.13u W=0.74u
+ AS=0.18945p AD=0.13135p PS=1.27u PD=1.095u
M$830 \$537 A1|X$1 \$526 15|25|VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.13135p
+ AD=0.1628p PS=1.095u PD=1.18u
M$831 \$526 A0|X \$536 15|25|VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.1628p
+ AD=0.3367p PS=1.18u PD=1.65u
M$832 \$536 \$525 15|25|VSS 15|25|VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.3367p
+ AD=0.148p PS=1.65u PD=1.14u
M$833 15|25|VSS \$526 A|X$36 15|25|VSS sg13_lv_nmos L=0.13u W=1.48u AS=0.3515p
+ AD=0.518p PS=2.43u PD=3.62u
M$835 \$527 A|X$45 15|25|VSS 15|25|VSS sg13_lv_nmos L=0.13u W=0.42u AS=0.1428p
+ AD=0.0798p PS=1.52u PD=0.8u
M$836 15|25|VSS \$527 \$528 15|25|VSS sg13_lv_nmos L=0.5u W=0.42u AS=0.0798p
+ AD=0.1428p PS=0.8u PD=1.52u
M$837 15|25|VSS \$528 \$529 15|25|VSS sg13_lv_nmos L=0.5u W=0.42u AS=0.1426p
+ AD=0.1428p PS=1.16u PD=1.52u
M$838 15|25|VSS \$529 A|X$47 15|25|VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.1426p
+ AD=0.2516p PS=1.16u PD=2.16u
M$839 \$544 A|X$47 15|25|VSS 15|25|VSS sg13_lv_nmos L=0.13u W=0.42u AS=0.1428p
+ AD=0.0798p PS=1.52u PD=0.8u
M$840 15|25|VSS \$544 \$545 15|25|VSS sg13_lv_nmos L=0.5u W=0.42u AS=0.0798p
+ AD=0.1428p PS=0.8u PD=1.52u
M$841 15|25|VSS 13|S|VSEL_DT \$531 15|25|VSS sg13_lv_nmos L=0.13u W=0.55u
+ AS=0.18945p AD=0.187p PS=1.27u PD=1.78u
M$842 15|25|VSS 13|S|VSEL_DT \$535 15|25|VSS sg13_lv_nmos L=0.13u W=0.74u
+ AS=0.18945p AD=0.13135p PS=1.27u PD=1.095u
M$843 \$535 A1|X \$532 15|25|VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.13135p
+ AD=0.1628p PS=1.095u PD=1.18u
M$844 \$532 A0|X$1 \$534 15|25|VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.1628p
+ AD=0.3367p PS=1.18u PD=1.65u
M$845 \$534 \$531 15|25|VSS 15|25|VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.3367p
+ AD=0.148p PS=1.65u PD=1.14u
M$846 15|25|VSS \$532 A|B|X 15|25|VSS sg13_lv_nmos L=0.13u W=1.48u AS=0.3515p
+ AD=0.518p PS=2.43u PD=3.62u
M$848 \$546 \$545 15|25|VSS 15|25|VSS sg13_lv_nmos L=0.5u W=0.42u AS=0.1428p
+ AD=0.1426p PS=1.52u PD=1.16u
M$849 15|25|VSS \$546 A0|X$1 15|25|VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.1426p
+ AD=0.2516p PS=1.16u PD=2.16u
M$850 15|25|VSS A|Y$16 A|Y$15 15|25|VSS sg13_lv_nmos L=0.13u W=1.48u AS=0.3922p
+ AD=0.3959p PS=3.28u PD=3.29u
M$852 \$572 NOC_P|X 15|25|VSS 15|25|VSS sg13_lv_nmos L=0.13u W=2.24u AS=1.0528p
+ AD=1.0528p PS=5.24u PD=5.24u
M$854 \$574 NOC_N|X 15|25|VSS 15|25|VSS sg13_lv_nmos L=0.13u W=2.24u AS=1.0528p
+ AD=1.0528p PS=5.24u PD=5.24u
M$856 6 6 6 6 sg13_hv_nmos L=0.45u W=88u AS=23.04p AD=23.04p PS=138.08u
+ PD=138.08u
M$857 6 \$81 8 6 sg13_hv_nmos L=0.45u W=32u AS=8p AD=8p PS=48u PD=48u
M$890 6 \$82 \$81 6 sg13_hv_nmos L=0.45u W=16u AS=4p AD=4p PS=24u PD=24u
M$907 6 \$83 \$82 6 sg13_hv_nmos L=0.45u W=8u AS=2p AD=2p PS=12u PD=12u
M$916 6 \$84 \$83 6 sg13_hv_nmos L=0.45u W=4u AS=1p AD=1p PS=6u PD=6u
M$921 6 \$85 \$84 6 sg13_hv_nmos L=0.45u W=2u AS=0.5p AD=0.5p PS=3u PD=3u
M$924 6 6 \$85 6 sg13_hv_nmos L=0.45u W=1u AS=0.25p AD=0.25p PS=1.5u PD=1.5u
M$925 \$85 \$86 6 6 sg13_hv_nmos L=0.45u W=1u AS=0.25p AD=0.25p PS=1.5u PD=1.5u
M$998 5 5 5 5 sg13_hv_nmos L=0.45u W=88u AS=23.04p AD=23.04p PS=138.08u
+ PD=138.08u
M$999 5 \$93 \$102 5 sg13_hv_nmos L=0.45u W=1u AS=0.25p AD=0.25p PS=1.5u PD=1.5u
M$1000 \$102 5 5 5 sg13_hv_nmos L=0.45u W=1u AS=0.25p AD=0.25p PS=1.5u PD=1.5u
M$1002 5 \$102 \$103 5 sg13_hv_nmos L=0.45u W=2u AS=0.5p AD=0.5p PS=3u PD=3u
M$1005 5 \$103 \$104 5 sg13_hv_nmos L=0.45u W=4u AS=1p AD=1p PS=6u PD=6u
M$1010 5 \$104 \$106 5 sg13_hv_nmos L=0.45u W=8u AS=2p AD=2p PS=12u PD=12u
M$1019 5 \$106 \$107 5 sg13_hv_nmos L=0.45u W=16u AS=4p AD=4p PS=24u PD=24u
M$1036 5 \$107 7 5 sg13_hv_nmos L=0.45u W=32u AS=8p AD=8p PS=48u PD=48u
M$1140 6 6 \$172 6 sg13_hv_nmos L=5u W=2u AS=1.02p AD=0.5p PS=5.02u PD=2.5u
M$1141 \$172 6 \$164 6 sg13_hv_nmos L=5u W=2u AS=0.5p AD=0.5p PS=2.5u PD=2.5u
M$1142 \$164 6 6 6 sg13_hv_nmos L=5u W=2u AS=0.5p AD=1.02p PS=2.5u PD=5.02u
M$1143 6 6 \$173 6 sg13_hv_nmos L=5u W=2u AS=1.02p AD=0.5p PS=5.02u PD=2.5u
M$1144 \$173 \$170 \$165 6 sg13_hv_nmos L=5u W=2u AS=0.5p AD=0.5p PS=2.5u
+ PD=2.5u
M$1145 \$165 6 6 6 sg13_hv_nmos L=5u W=2u AS=0.5p AD=1.02p PS=2.5u PD=5.02u
M$1146 6 6 \$174 6 sg13_hv_nmos L=5u W=2u AS=1.02p AD=0.5p PS=5.02u PD=2.5u
M$1147 \$174 \$165 \$166 6 sg13_hv_nmos L=5u W=2u AS=0.5p AD=0.5p PS=2.5u
+ PD=2.5u
M$1148 \$166 6 6 6 sg13_hv_nmos L=5u W=2u AS=0.5p AD=1.02p PS=2.5u PD=5.02u
M$1149 6 6 \$175 6 sg13_hv_nmos L=5u W=2u AS=1.02p AD=0.5p PS=5.02u PD=2.5u
M$1150 \$175 \$166 \$167 6 sg13_hv_nmos L=5u W=2u AS=0.5p AD=0.5p PS=2.5u
+ PD=2.5u
M$1151 \$167 6 6 6 sg13_hv_nmos L=5u W=2u AS=0.5p AD=1.02p PS=2.5u PD=5.02u
M$1152 6 6 \$176 6 sg13_hv_nmos L=5u W=2u AS=1.02p AD=0.5p PS=5.02u PD=2.5u
M$1153 \$176 \$167 \$168 6 sg13_hv_nmos L=5u W=2u AS=0.5p AD=0.5p PS=2.5u
+ PD=2.5u
M$1154 \$168 6 6 6 sg13_hv_nmos L=5u W=2u AS=0.5p AD=1.02p PS=2.5u PD=5.02u
M$1155 6 6 \$177 6 sg13_hv_nmos L=5u W=2u AS=1.02p AD=0.5p PS=5.02u PD=2.5u
M$1156 \$177 \$168 \$170 6 sg13_hv_nmos L=5u W=2u AS=0.5p AD=0.5p PS=2.5u
+ PD=2.5u
M$1157 \$170 6 6 6 sg13_hv_nmos L=5u W=2u AS=0.5p AD=1.02p PS=2.5u PD=5.02u
M$1158 6 6 \$178 6 sg13_hv_nmos L=5u W=2u AS=1.02p AD=0.5p PS=5.02u PD=2.5u
M$1159 \$178 6 \$169 6 sg13_hv_nmos L=5u W=2u AS=0.5p AD=0.5p PS=2.5u PD=2.5u
M$1160 \$169 6 6 6 sg13_hv_nmos L=5u W=2u AS=0.5p AD=1.02p PS=2.5u PD=5.02u
M$1161 6 6 6 6 sg13_hv_nmos L=0.5u W=35u AS=14.21p AD=10.57p PS=84.42u PD=63.14u
M$1162 6 \$140 \$150 6 sg13_hv_nmos L=0.5u W=5u AS=1.25p AD=1.25p PS=7.5u
+ PD=7.5u
M$1167 \$150 6 6 6 sg13_hv_nmos L=0.5u W=1u AS=0.25p AD=0.51p PS=1.5u PD=3.02u
M$1169 6 \$141 \$151 6 sg13_hv_nmos L=0.5u W=5u AS=1.25p AD=1.25p PS=7.5u
+ PD=7.5u
M$1174 \$151 6 6 6 sg13_hv_nmos L=0.5u W=1u AS=0.25p AD=0.51p PS=1.5u PD=3.02u
M$1176 6 \$142 \$152 6 sg13_hv_nmos L=0.5u W=5u AS=1.25p AD=1.25p PS=7.5u
+ PD=7.5u
M$1181 \$152 6 6 6 sg13_hv_nmos L=0.5u W=1u AS=0.25p AD=0.51p PS=1.5u PD=3.02u
M$1183 6 \$143 \$153 6 sg13_hv_nmos L=0.5u W=5u AS=1.25p AD=1.25p PS=7.5u
+ PD=7.5u
M$1188 \$153 6 6 6 sg13_hv_nmos L=0.5u W=1u AS=0.25p AD=0.51p PS=1.5u PD=3.02u
M$1190 6 \$144 \$154 6 sg13_hv_nmos L=0.5u W=5u AS=1.25p AD=1.25p PS=7.5u
+ PD=7.5u
M$1195 \$154 6 6 6 sg13_hv_nmos L=0.5u W=1u AS=0.25p AD=0.51p PS=1.5u PD=3.02u
M$1197 6 \$145 \$155 6 sg13_hv_nmos L=0.5u W=5u AS=1.25p AD=1.25p PS=7.5u
+ PD=7.5u
M$1202 \$155 6 6 6 sg13_hv_nmos L=0.5u W=1u AS=0.25p AD=0.51p PS=1.5u PD=3.02u
M$1204 6 \$146 \$156 6 sg13_hv_nmos L=0.5u W=5u AS=1.25p AD=1.25p PS=7.5u
+ PD=7.5u
M$1209 \$156 6 6 6 sg13_hv_nmos L=0.5u W=1u AS=0.25p AD=0.51p PS=1.5u PD=3.02u
M$1211 6 6 \$172 6 sg13_hv_nmos L=0.5u W=1u AS=0.25p AD=0.25p PS=1.5u PD=1.5u
M$1212 \$172 \$140 6 6 sg13_hv_nmos L=0.5u W=3u AS=0.75p AD=0.75p PS=4.5u
+ PD=4.5u
M$1218 6 6 \$173 6 sg13_hv_nmos L=0.5u W=1u AS=0.25p AD=0.25p PS=1.5u PD=1.5u
M$1219 \$173 \$141 6 6 sg13_hv_nmos L=0.5u W=3u AS=0.75p AD=0.75p PS=4.5u
+ PD=4.5u
M$1225 6 6 \$174 6 sg13_hv_nmos L=0.5u W=1u AS=0.25p AD=0.25p PS=1.5u PD=1.5u
M$1226 \$174 \$142 6 6 sg13_hv_nmos L=0.5u W=3u AS=0.75p AD=0.75p PS=4.5u
+ PD=4.5u
M$1232 6 6 \$175 6 sg13_hv_nmos L=0.5u W=1u AS=0.25p AD=0.25p PS=1.5u PD=1.5u
M$1233 \$175 \$143 6 6 sg13_hv_nmos L=0.5u W=3u AS=0.75p AD=0.75p PS=4.5u
+ PD=4.5u
M$1239 6 6 \$176 6 sg13_hv_nmos L=0.5u W=1u AS=0.25p AD=0.25p PS=1.5u PD=1.5u
M$1240 \$176 \$144 6 6 sg13_hv_nmos L=0.5u W=3u AS=0.75p AD=0.75p PS=4.5u
+ PD=4.5u
M$1246 6 6 \$177 6 sg13_hv_nmos L=0.5u W=1u AS=0.25p AD=0.25p PS=1.5u PD=1.5u
M$1247 \$177 \$145 6 6 sg13_hv_nmos L=0.5u W=3u AS=0.75p AD=0.75p PS=4.5u
+ PD=4.5u
M$1253 6 6 \$178 6 sg13_hv_nmos L=0.5u W=1u AS=0.25p AD=0.25p PS=1.5u PD=1.5u
M$1254 \$178 \$146 6 6 sg13_hv_nmos L=0.5u W=3u AS=0.75p AD=0.75p PS=4.5u
+ PD=4.5u
M$1260 6 \$140 \$140 6 sg13_hv_nmos L=0.5u W=5u AS=1.25p AD=1.25p PS=7.5u
+ PD=7.5u
M$1265 \$140 6 6 6 sg13_hv_nmos L=0.5u W=1u AS=0.25p AD=0.51p PS=1.5u PD=3.02u
M$1267 6 \$141 \$141 6 sg13_hv_nmos L=0.5u W=5u AS=1.25p AD=1.25p PS=7.5u
+ PD=7.5u
M$1272 \$141 6 6 6 sg13_hv_nmos L=0.5u W=1u AS=0.25p AD=0.51p PS=1.5u PD=3.02u
M$1274 6 \$142 \$142 6 sg13_hv_nmos L=0.5u W=5u AS=1.25p AD=1.25p PS=7.5u
+ PD=7.5u
M$1279 \$142 6 6 6 sg13_hv_nmos L=0.5u W=1u AS=0.25p AD=0.51p PS=1.5u PD=3.02u
M$1281 6 \$143 \$143 6 sg13_hv_nmos L=0.5u W=5u AS=1.25p AD=1.25p PS=7.5u
+ PD=7.5u
M$1286 \$143 6 6 6 sg13_hv_nmos L=0.5u W=1u AS=0.25p AD=0.51p PS=1.5u PD=3.02u
M$1288 6 \$144 \$144 6 sg13_hv_nmos L=0.5u W=5u AS=1.25p AD=1.25p PS=7.5u
+ PD=7.5u
M$1293 \$144 6 6 6 sg13_hv_nmos L=0.5u W=1u AS=0.25p AD=0.51p PS=1.5u PD=3.02u
M$1295 6 \$145 \$145 6 sg13_hv_nmos L=0.5u W=5u AS=1.25p AD=1.25p PS=7.5u
+ PD=7.5u
M$1300 \$145 6 6 6 sg13_hv_nmos L=0.5u W=1u AS=0.25p AD=0.51p PS=1.5u PD=3.02u
M$1302 6 \$146 \$146 6 sg13_hv_nmos L=0.5u W=5u AS=1.25p AD=1.25p PS=7.5u
+ PD=7.5u
M$1307 \$146 6 6 6 sg13_hv_nmos L=0.5u W=1u AS=0.25p AD=0.51p PS=1.5u PD=3.02u
M$1308 5 5 5 5 sg13_hv_nmos L=0.5u W=35u AS=14.21p AD=10.57p PS=84.42u PD=63.14u
M$1309 5 \$204 \$204 5 sg13_hv_nmos L=0.5u W=5u AS=1.25p AD=1.25p PS=7.5u
+ PD=7.5u
M$1314 \$204 5 5 5 sg13_hv_nmos L=0.5u W=1u AS=0.25p AD=0.51p PS=1.5u PD=3.02u
M$1316 5 \$205 \$205 5 sg13_hv_nmos L=0.5u W=5u AS=1.25p AD=1.25p PS=7.5u
+ PD=7.5u
M$1321 \$205 5 5 5 sg13_hv_nmos L=0.5u W=1u AS=0.25p AD=0.51p PS=1.5u PD=3.02u
M$1323 5 \$206 \$206 5 sg13_hv_nmos L=0.5u W=5u AS=1.25p AD=1.25p PS=7.5u
+ PD=7.5u
M$1328 \$206 5 5 5 sg13_hv_nmos L=0.5u W=1u AS=0.25p AD=0.51p PS=1.5u PD=3.02u
M$1330 5 \$207 \$207 5 sg13_hv_nmos L=0.5u W=5u AS=1.25p AD=1.25p PS=7.5u
+ PD=7.5u
M$1335 \$207 5 5 5 sg13_hv_nmos L=0.5u W=1u AS=0.25p AD=0.51p PS=1.5u PD=3.02u
M$1337 5 \$208 \$208 5 sg13_hv_nmos L=0.5u W=5u AS=1.25p AD=1.25p PS=7.5u
+ PD=7.5u
M$1342 \$208 5 5 5 sg13_hv_nmos L=0.5u W=1u AS=0.25p AD=0.51p PS=1.5u PD=3.02u
M$1351 6 6 \$184 6 sg13_hv_nmos L=0.45u W=1u AS=0.25p AD=0.25p PS=1.5u PD=1.5u
M$1352 \$184 \$168 6 6 sg13_hv_nmos L=0.45u W=1u AS=0.25p AD=0.25p PS=1.5u
+ PD=1.5u
M$1354 6 \$184 \$86 6 sg13_hv_nmos L=0.45u W=2u AS=0.5p AD=0.5p PS=3u PD=3u
M$1365 5 5 \$195 5 sg13_hv_nmos L=0.45u W=1u AS=0.25p AD=0.25p PS=1.5u PD=1.5u
M$1366 \$195 \$194 5 5 sg13_hv_nmos L=0.45u W=1u AS=0.25p AD=0.25p PS=1.5u
+ PD=1.5u
M$1368 5 \$195 \$93 5 sg13_hv_nmos L=0.45u W=2u AS=0.5p AD=0.5p PS=3u PD=3u
M$1372 5 \$209 \$209 5 sg13_hv_nmos L=0.5u W=5u AS=1.25p AD=1.25p PS=7.5u
+ PD=7.5u
M$1377 \$209 5 5 5 sg13_hv_nmos L=0.5u W=1u AS=0.25p AD=0.51p PS=1.5u PD=3.02u
M$1379 5 \$210 \$210 5 sg13_hv_nmos L=0.5u W=5u AS=1.25p AD=1.25p PS=7.5u
+ PD=7.5u
M$1384 \$210 5 5 5 sg13_hv_nmos L=0.5u W=1u AS=0.25p AD=0.51p PS=1.5u PD=3.02u
M$1386 5 5 \$214 5 sg13_hv_nmos L=0.5u W=1u AS=0.25p AD=0.25p PS=1.5u PD=1.5u
M$1387 \$214 \$204 5 5 sg13_hv_nmos L=0.5u W=3u AS=0.75p AD=0.75p PS=4.5u
+ PD=4.5u
M$1393 5 5 \$215 5 sg13_hv_nmos L=0.5u W=1u AS=0.25p AD=0.25p PS=1.5u PD=1.5u
M$1394 \$215 \$205 5 5 sg13_hv_nmos L=0.5u W=3u AS=0.75p AD=0.75p PS=4.5u
+ PD=4.5u
M$1400 5 5 \$216 5 sg13_hv_nmos L=0.5u W=1u AS=0.25p AD=0.25p PS=1.5u PD=1.5u
M$1401 \$216 \$206 5 5 sg13_hv_nmos L=0.5u W=3u AS=0.75p AD=0.75p PS=4.5u
+ PD=4.5u
M$1407 5 5 \$217 5 sg13_hv_nmos L=0.5u W=1u AS=0.25p AD=0.25p PS=1.5u PD=1.5u
M$1408 \$217 \$207 5 5 sg13_hv_nmos L=0.5u W=3u AS=0.75p AD=0.75p PS=4.5u
+ PD=4.5u
M$1414 5 5 \$218 5 sg13_hv_nmos L=0.5u W=1u AS=0.25p AD=0.25p PS=1.5u PD=1.5u
M$1415 \$218 \$208 5 5 sg13_hv_nmos L=0.5u W=3u AS=0.75p AD=0.75p PS=4.5u
+ PD=4.5u
M$1421 5 5 \$219 5 sg13_hv_nmos L=0.5u W=1u AS=0.25p AD=0.25p PS=1.5u PD=1.5u
M$1422 \$219 \$209 5 5 sg13_hv_nmos L=0.5u W=3u AS=0.75p AD=0.75p PS=4.5u
+ PD=4.5u
M$1428 5 5 \$220 5 sg13_hv_nmos L=0.5u W=1u AS=0.25p AD=0.25p PS=1.5u PD=1.5u
M$1429 \$220 \$210 5 5 sg13_hv_nmos L=0.5u W=3u AS=0.75p AD=0.75p PS=4.5u
+ PD=4.5u
M$1435 5 \$204 \$224 5 sg13_hv_nmos L=0.5u W=5u AS=1.25p AD=1.25p PS=7.5u
+ PD=7.5u
M$1440 \$224 5 5 5 sg13_hv_nmos L=0.5u W=1u AS=0.25p AD=0.51p PS=1.5u PD=3.02u
M$1442 5 \$205 \$225 5 sg13_hv_nmos L=0.5u W=5u AS=1.25p AD=1.25p PS=7.5u
+ PD=7.5u
M$1447 \$225 5 5 5 sg13_hv_nmos L=0.5u W=1u AS=0.25p AD=0.51p PS=1.5u PD=3.02u
M$1449 5 \$206 \$226 5 sg13_hv_nmos L=0.5u W=5u AS=1.25p AD=1.25p PS=7.5u
+ PD=7.5u
M$1454 \$226 5 5 5 sg13_hv_nmos L=0.5u W=1u AS=0.25p AD=0.51p PS=1.5u PD=3.02u
M$1456 5 \$207 \$227 5 sg13_hv_nmos L=0.5u W=5u AS=1.25p AD=1.25p PS=7.5u
+ PD=7.5u
M$1461 \$227 5 5 5 sg13_hv_nmos L=0.5u W=1u AS=0.25p AD=0.51p PS=1.5u PD=3.02u
M$1463 5 \$208 \$228 5 sg13_hv_nmos L=0.5u W=5u AS=1.25p AD=1.25p PS=7.5u
+ PD=7.5u
M$1468 \$228 5 5 5 sg13_hv_nmos L=0.5u W=1u AS=0.25p AD=0.51p PS=1.5u PD=3.02u
M$1470 5 \$209 \$229 5 sg13_hv_nmos L=0.5u W=5u AS=1.25p AD=1.25p PS=7.5u
+ PD=7.5u
M$1475 \$229 5 5 5 sg13_hv_nmos L=0.5u W=1u AS=0.25p AD=0.51p PS=1.5u PD=3.02u
M$1477 5 \$210 \$230 5 sg13_hv_nmos L=0.5u W=5u AS=1.25p AD=1.25p PS=7.5u
+ PD=7.5u
M$1482 \$230 5 5 5 sg13_hv_nmos L=0.5u W=1u AS=0.25p AD=0.51p PS=1.5u PD=3.02u
M$1483 5 5 \$214 5 sg13_hv_nmos L=5u W=2u AS=1.02p AD=0.5p PS=5.02u PD=2.5u
M$1484 \$214 5 \$236 5 sg13_hv_nmos L=5u W=2u AS=0.5p AD=0.5p PS=2.5u PD=2.5u
M$1485 \$236 5 5 5 sg13_hv_nmos L=5u W=2u AS=0.5p AD=1.02p PS=2.5u PD=5.02u
M$1486 5 5 \$215 5 sg13_hv_nmos L=5u W=2u AS=1.02p AD=0.5p PS=5.02u PD=2.5u
M$1487 \$215 \$199 \$238 5 sg13_hv_nmos L=5u W=2u AS=0.5p AD=0.5p PS=2.5u
+ PD=2.5u
M$1488 \$238 5 5 5 sg13_hv_nmos L=5u W=2u AS=0.5p AD=1.02p PS=2.5u PD=5.02u
M$1489 5 5 \$216 5 sg13_hv_nmos L=5u W=2u AS=1.02p AD=0.5p PS=5.02u PD=2.5u
M$1490 \$216 \$238 \$239 5 sg13_hv_nmos L=5u W=2u AS=0.5p AD=0.5p PS=2.5u
+ PD=2.5u
M$1491 \$239 5 5 5 sg13_hv_nmos L=5u W=2u AS=0.5p AD=1.02p PS=2.5u PD=5.02u
M$1492 5 5 \$217 5 sg13_hv_nmos L=5u W=2u AS=1.02p AD=0.5p PS=5.02u PD=2.5u
M$1493 \$217 \$239 \$240 5 sg13_hv_nmos L=5u W=2u AS=0.5p AD=0.5p PS=2.5u
+ PD=2.5u
M$1494 \$240 5 5 5 sg13_hv_nmos L=5u W=2u AS=0.5p AD=1.02p PS=2.5u PD=5.02u
M$1495 5 5 \$218 5 sg13_hv_nmos L=5u W=2u AS=1.02p AD=0.5p PS=5.02u PD=2.5u
M$1496 \$218 \$240 \$194 5 sg13_hv_nmos L=5u W=2u AS=0.5p AD=0.5p PS=2.5u
+ PD=2.5u
M$1497 \$194 5 5 5 sg13_hv_nmos L=5u W=2u AS=0.5p AD=1.02p PS=2.5u PD=5.02u
M$1498 5 5 \$219 5 sg13_hv_nmos L=5u W=2u AS=1.02p AD=0.5p PS=5.02u PD=2.5u
M$1499 \$219 \$194 \$199 5 sg13_hv_nmos L=5u W=2u AS=0.5p AD=0.5p PS=2.5u
+ PD=2.5u
M$1500 \$199 5 5 5 sg13_hv_nmos L=5u W=2u AS=0.5p AD=1.02p PS=2.5u PD=5.02u
M$1501 5 5 \$220 5 sg13_hv_nmos L=5u W=2u AS=1.02p AD=0.5p PS=5.02u PD=2.5u
M$1502 \$220 5 \$237 5 sg13_hv_nmos L=5u W=2u AS=0.5p AD=0.5p PS=2.5u PD=2.5u
M$1503 \$237 5 5 5 sg13_hv_nmos L=5u W=2u AS=0.5p AD=1.02p PS=2.5u PD=5.02u
M$1504 A \$93 15|25|VSS 15|25|VSS sg13_hv_nmos L=0.45u W=1u AS=0.77p AD=0.77p
+ PS=3.54u PD=3.54u
M$1505 A$1 \$86 15|25|VSS 15|25|VSS sg13_hv_nmos L=0.45u W=1u AS=0.77p AD=0.77p
+ PS=3.54u PD=3.54u
M$1506 \$414 \$563 20 20 sg13_hv_nmos L=0.45u W=2000u AS=510.4p AD=510.4p
+ PS=2142.08u PD=2142.08u
M$1606 \$562 \$564 20 20 sg13_hv_nmos L=0.45u W=2000u AS=510.4p AD=510.4p
+ PS=2142.08u PD=2142.08u
M$1906 20 20 20 20 sg13_hv_nmos L=0.45u W=1316u AS=340.44p AD=340.44p
+ PS=1500.16u PD=1500.16u
M$1963 20 NOC_P|X \$563 20 sg13_hv_nmos L=0.45u W=250u AS=62.5p AD=62.5p
+ PS=262.5u PD=262.5u
M$1988 \$563 20 20 20 sg13_hv_nmos L=0.45u W=10u AS=2.5p AD=2.5p PS=10.5u
+ PD=10.5u
M$1989 20 20 \$567 20 sg13_hv_nmos L=0.45u W=20u AS=5p AD=5p PS=21u PD=21u
M$1990 \$567 \$572 20 20 sg13_hv_nmos L=0.45u W=60u AS=15p AD=15p PS=63u PD=63u
M$1997 20 20 \$568 20 sg13_hv_nmos L=0.45u W=20u AS=5p AD=5p PS=21u PD=21u
M$1998 \$568 NOC_P|X 20 20 sg13_hv_nmos L=0.45u W=60u AS=15p AD=15p PS=63u
+ PD=63u
M$2063 20 NOC_N|X \$564 20 sg13_hv_nmos L=0.45u W=250u AS=62.5p AD=62.5p
+ PS=262.5u PD=262.5u
M$2088 \$564 20 20 20 sg13_hv_nmos L=0.45u W=10u AS=2.5p AD=2.5p PS=10.5u
+ PD=10.5u
M$2089 20 20 \$569 20 sg13_hv_nmos L=0.45u W=20u AS=5p AD=5p PS=21u PD=21u
M$2090 \$569 \$574 20 20 sg13_hv_nmos L=0.45u W=60u AS=15p AD=15p PS=63u PD=63u
M$2097 20 20 \$570 20 sg13_hv_nmos L=0.45u W=20u AS=5p AD=5p PS=21u PD=21u
M$2098 \$570 NOC_N|X 20 20 sg13_hv_nmos L=0.45u W=60u AS=15p AD=15p PS=63u
+ PD=63u
M$2106 27 \$562 26 26 sg13_hv_nmos L=0.45u W=40800u AS=14616p AD=14616p
+ PS=44523.2u PD=44523.2u
M$5442 20 \$623 21 20 sg13_hv_nmos L=0.45u W=32u AS=8p AD=8p PS=48u PD=48u
M$5475 20 \$627 \$623 20 sg13_hv_nmos L=0.45u W=16u AS=4p AD=4p PS=24u PD=24u
M$5492 20 \$634 \$627 20 sg13_hv_nmos L=0.45u W=8u AS=2p AD=2p PS=12u PD=12u
M$5501 20 \$635 \$634 20 sg13_hv_nmos L=0.45u W=4u AS=1p AD=1p PS=6u PD=6u
M$5506 20 \$637 \$635 20 sg13_hv_nmos L=0.45u W=2u AS=0.5p AD=0.5p PS=3u PD=3u
M$5509 20 20 \$637 20 sg13_hv_nmos L=0.45u W=1u AS=0.25p AD=0.25p PS=1.5u
+ PD=1.5u
M$5510 \$637 \$562 20 20 sg13_hv_nmos L=0.45u W=1u AS=0.25p AD=0.25p PS=1.5u
+ PD=1.5u
M$6400 20 \$414 \$651 20 sg13_hv_nmos L=0.45u W=1u AS=0.25p AD=0.25p PS=1.5u
+ PD=1.5u
M$6401 \$651 20 20 20 sg13_hv_nmos L=0.45u W=1u AS=0.25p AD=0.25p PS=1.5u
+ PD=1.5u
M$6403 20 \$651 \$652 20 sg13_hv_nmos L=0.45u W=2u AS=0.5p AD=0.5p PS=3u PD=3u
M$6406 20 \$652 \$653 20 sg13_hv_nmos L=0.45u W=4u AS=1p AD=1p PS=6u PD=6u
M$6411 20 \$653 \$654 20 sg13_hv_nmos L=0.45u W=8u AS=2p AD=2p PS=12u PD=12u
M$6420 20 \$654 \$655 20 sg13_hv_nmos L=0.45u W=16u AS=4p AD=4p PS=24u PD=24u
M$6437 20 \$655 22 20 sg13_hv_nmos L=0.45u W=32u AS=8p AD=8p PS=48u PD=48u
M$6470 19|VDD A A|Y 19|VDD sg13_lv_pmos L=0.13u W=1.12u AS=0.392p AD=0.392p
+ PS=2.94u PD=2.94u
M$6471 19|VDD A$1 A|Y$1 19|VDD sg13_lv_pmos L=0.13u W=1.12u AS=0.392p AD=0.392p
+ PS=2.94u PD=2.94u
M$6472 19|VDD A|Y \$245 19|VDD sg13_lv_pmos L=0.13u W=1.68u AS=0.4452p
+ AD=0.3626p PS=3.58u PD=2.72u
M$6474 19|VDD \$245 A|VINS|X 19|VDD sg13_lv_pmos L=0.13u W=4.48u AS=0.8414p
+ AD=1.0192p PS=6u PD=7.42u
M$6478 19|VDD A|Y$1 \$246 19|VDD sg13_lv_pmos L=0.13u W=1.68u AS=0.4452p
+ AD=0.3626p PS=3.58u PD=2.72u
M$6480 19|VDD \$246 A|VINR|X 19|VDD sg13_lv_pmos L=0.13u W=4.48u AS=0.8414p
+ AD=1.0192p PS=6u PD=7.42u
M$6484 19|VDD \$259 16|PD_BUFF|X 19|VDD sg13_lv_pmos L=0.13u W=17.92u
+ AS=3.5896p AD=3.4048p PS=25.45u PD=24u
M$6500 19|VDD A|X \$259 19|VDD sg13_lv_pmos L=0.13u W=6.72u AS=1.2768p
+ AD=1.4448p PS=9u PD=10.42u
M$6506 19|VDD \$261 VINS_BUFF|X 19|VDD sg13_lv_pmos L=0.13u W=17.92u AS=3.5896p
+ AD=3.4048p PS=25.45u PD=24u
M$6522 19|VDD A|X$1 \$261 19|VDD sg13_lv_pmos L=0.13u W=6.72u AS=1.2768p
+ AD=1.4448p PS=9u PD=10.42u
M$6528 19|VDD \$263 17|NOC_N_BUFF|X 19|VDD sg13_lv_pmos L=0.13u W=17.92u
+ AS=3.5896p AD=3.4048p PS=25.45u PD=24u
M$6544 19|VDD A|X$2 \$263 19|VDD sg13_lv_pmos L=0.13u W=6.72u AS=1.2768p
+ AD=1.4448p PS=9u PD=10.42u
M$6550 19|VDD \$266 16|PD_BUFF|X 19|VDD sg13_lv_pmos L=0.13u W=17.92u
+ AS=3.5896p AD=3.4048p PS=25.45u PD=24u
M$6566 19|VDD A|X \$266 19|VDD sg13_lv_pmos L=0.13u W=6.72u AS=1.2768p
+ AD=1.4448p PS=9u PD=10.42u
M$6572 19|VDD \$267 VINS_BUFF|X 19|VDD sg13_lv_pmos L=0.13u W=17.92u AS=3.5896p
+ AD=3.4048p PS=25.45u PD=24u
M$6588 19|VDD A|X$1 \$267 19|VDD sg13_lv_pmos L=0.13u W=6.72u AS=1.2768p
+ AD=1.4448p PS=9u PD=10.42u
M$6594 19|VDD \$268 17|NOC_N_BUFF|X 19|VDD sg13_lv_pmos L=0.13u W=17.92u
+ AS=3.5896p AD=3.4048p PS=25.45u PD=24u
M$6610 19|VDD A|X$2 \$268 19|VDD sg13_lv_pmos L=0.13u W=6.72u AS=1.2768p
+ AD=1.4448p PS=9u PD=10.42u
M$6616 19|VDD \$269 16|PD_BUFF|X 19|VDD sg13_lv_pmos L=0.13u W=17.92u
+ AS=3.5896p AD=3.4048p PS=25.45u PD=24u
M$6632 19|VDD A|X \$269 19|VDD sg13_lv_pmos L=0.13u W=6.72u AS=1.2768p
+ AD=1.4448p PS=9u PD=10.42u
M$6638 19|VDD \$270 VINS_BUFF|X 19|VDD sg13_lv_pmos L=0.13u W=17.92u AS=3.5896p
+ AD=3.4048p PS=25.45u PD=24u
M$6654 19|VDD A|X$1 \$270 19|VDD sg13_lv_pmos L=0.13u W=6.72u AS=1.2768p
+ AD=1.4448p PS=9u PD=10.42u
M$6660 19|VDD \$271 17|NOC_N_BUFF|X 19|VDD sg13_lv_pmos L=0.13u W=17.92u
+ AS=3.5896p AD=3.4048p PS=25.45u PD=24u
M$6676 19|VDD A|X$2 \$271 19|VDD sg13_lv_pmos L=0.13u W=6.72u AS=1.2768p
+ AD=1.4448p PS=9u PD=10.42u
M$6682 19|VDD \$272 16|PD_BUFF|X 19|VDD sg13_lv_pmos L=0.13u W=17.92u
+ AS=3.5896p AD=3.4048p PS=25.45u PD=24u
M$6698 19|VDD A|X \$272 19|VDD sg13_lv_pmos L=0.13u W=6.72u AS=1.2768p
+ AD=1.4448p PS=9u PD=10.42u
M$6704 19|VDD \$275 A|X 19|VDD sg13_lv_pmos L=0.13u W=17.92u AS=3.5896p
+ AD=3.4048p PS=25.45u PD=24u
M$6720 19|VDD A|X$3 \$275 19|VDD sg13_lv_pmos L=0.13u W=6.72u AS=1.2768p
+ AD=1.4448p PS=9u PD=10.42u
M$6726 19|VDD \$273 VINS_BUFF|X 19|VDD sg13_lv_pmos L=0.13u W=17.92u AS=3.5896p
+ AD=3.4048p PS=25.45u PD=24u
M$6742 19|VDD A|X$1 \$273 19|VDD sg13_lv_pmos L=0.13u W=6.72u AS=1.2768p
+ AD=1.4448p PS=9u PD=10.42u
M$6748 19|VDD \$274 17|NOC_N_BUFF|X 19|VDD sg13_lv_pmos L=0.13u W=17.92u
+ AS=3.5896p AD=3.4048p PS=25.45u PD=24u
M$6764 19|VDD A|X$2 \$274 19|VDD sg13_lv_pmos L=0.13u W=6.72u AS=1.2768p
+ AD=1.4448p PS=9u PD=10.42u
M$6770 19|VDD \$277 14|VINR_BUFF|X 19|VDD sg13_lv_pmos L=0.13u W=17.92u
+ AS=3.5896p AD=3.4048p PS=25.45u PD=24u
M$6786 19|VDD A|X$4 \$277 19|VDD sg13_lv_pmos L=0.13u W=6.72u AS=1.2768p
+ AD=1.4448p PS=9u PD=10.42u
M$6792 19|VDD \$278 A|X$3 19|VDD sg13_lv_pmos L=0.13u W=4.48u AS=1.0192p
+ AD=0.8414p PS=7.42u PD=6u
M$6796 19|VDD A$2 \$278 19|VDD sg13_lv_pmos L=0.13u W=1.68u AS=0.3626p
+ AD=0.4452p PS=2.72u PD=3.58u
M$6798 \$280 A|B|Y$1 19|VDD 19|VDD sg13_lv_pmos L=0.13u W=0.84u AS=0.3024p
+ AD=0.2051p PS=2.4u PD=1.52u
M$6799 19|VDD \$280 A$2 19|VDD sg13_lv_pmos L=0.13u W=1.12u AS=0.2051p
+ AD=0.4032p PS=1.52u PD=2.96u
M$6800 \$282 A|VINR|X 19|VDD 19|VDD sg13_lv_pmos L=0.13u W=0.84u AS=0.3024p
+ AD=0.2051p PS=2.4u PD=1.52u
M$6801 19|VDD \$282 A$3 19|VDD sg13_lv_pmos L=0.13u W=1.12u AS=0.2051p
+ AD=0.4032p PS=1.52u PD=2.96u
M$6802 19|VDD A|Y$2 A|B|Y 19|VDD sg13_lv_pmos L=0.13u W=1.12u AS=0.392p
+ AD=0.392p PS=2.94u PD=2.94u
M$6803 19|VDD \$279 A|X$1 19|VDD sg13_lv_pmos L=0.13u W=17.92u AS=3.5896p
+ AD=3.4048p PS=25.45u PD=24u
M$6819 19|VDD A|X$5 \$279 19|VDD sg13_lv_pmos L=0.13u W=6.72u AS=1.2768p
+ AD=1.4448p PS=9u PD=10.42u
M$6825 19|VDD \$289 14|VINR_BUFF|X 19|VDD sg13_lv_pmos L=0.13u W=17.92u
+ AS=3.5896p AD=3.4048p PS=25.45u PD=24u
M$6841 19|VDD A|X$4 \$289 19|VDD sg13_lv_pmos L=0.13u W=6.72u AS=1.2768p
+ AD=1.4448p PS=9u PD=10.42u
M$6847 19|VDD \$290 A|X$4 19|VDD sg13_lv_pmos L=0.13u W=17.92u AS=3.5896p
+ AD=3.4048p PS=25.45u PD=24u
M$6863 19|VDD A|X$6 \$290 19|VDD sg13_lv_pmos L=0.13u W=6.72u AS=1.2768p
+ AD=1.4448p PS=9u PD=10.42u
M$6869 19|VDD A$3 \$292 19|VDD sg13_lv_pmos L=0.13u W=1.68u AS=0.3626p
+ AD=0.4452p PS=2.72u PD=3.58u
M$6871 19|VDD \$292 A|X$6 19|VDD sg13_lv_pmos L=0.13u W=4.48u AS=1.0192p
+ AD=0.8414p PS=7.42u PD=6u
M$6875 \$299 \$298 19|VDD 19|VDD sg13_lv_pmos L=0.5u W=1u AS=0.34p AD=0.2254p
+ PS=2.68u PD=1.53u
M$6876 19|VDD \$299 A|X$8 19|VDD sg13_lv_pmos L=0.13u W=1.12u AS=0.2254p
+ AD=0.4256p PS=1.53u PD=3u
M$6877 19|VDD A|VINR|X A|Y$2 19|VDD sg13_lv_pmos L=0.13u W=2.24u AS=0.5964p
+ AD=0.5964p PS=4.425u PD=4.425u
M$6879 19|VDD A|Y$3 \$303 19|VDD sg13_lv_pmos L=0.13u W=0.84u AS=0.2856p
+ AD=0.1596p PS=2.36u PD=1.22u
M$6880 19|VDD A|B|Y \$303 19|VDD sg13_lv_pmos L=0.13u W=0.84u AS=0.1918p
+ AD=0.1596p PS=1.5u PD=1.22u
M$6881 19|VDD \$303 A|X$9 19|VDD sg13_lv_pmos L=0.13u W=2.24u AS=0.4046p
+ AD=0.6384p PS=3u PD=4.5u
M$6883 19|VDD A$4 \$294 19|VDD sg13_lv_pmos L=0.13u W=1.68u AS=0.3626p
+ AD=0.4452p PS=2.72u PD=3.58u
M$6885 19|VDD \$294 A|X$5 19|VDD sg13_lv_pmos L=0.13u W=4.48u AS=1.0192p
+ AD=0.8414p PS=7.42u PD=6u
M$6889 19|VDD \$295 A|X$2 19|VDD sg13_lv_pmos L=0.13u W=17.92u AS=3.5896p
+ AD=3.4048p PS=25.45u PD=24u
M$6905 19|VDD A|X$7 \$295 19|VDD sg13_lv_pmos L=0.13u W=6.72u AS=1.2768p
+ AD=1.4448p PS=9u PD=10.42u
M$6911 19|VDD \$312 14|VINR_BUFF|X 19|VDD sg13_lv_pmos L=0.13u W=17.92u
+ AS=3.5896p AD=3.4048p PS=25.45u PD=24u
M$6927 19|VDD A|X$4 \$312 19|VDD sg13_lv_pmos L=0.13u W=6.72u AS=1.2768p
+ AD=1.4448p PS=9u PD=10.42u
M$6933 19|VDD \$332 14|VINR_BUFF|X 19|VDD sg13_lv_pmos L=0.13u W=17.92u
+ AS=3.5896p AD=3.4048p PS=25.45u PD=24u
M$6949 19|VDD A|X$4 \$332 19|VDD sg13_lv_pmos L=0.13u W=6.72u AS=1.2768p
+ AD=1.4448p PS=9u PD=10.42u
M$6955 19|VDD A|Y$4 \$313 19|VDD sg13_lv_pmos L=0.13u W=0.42u AS=0.1523p
+ AD=0.1428p PS=1.38u PD=1.52u
M$6956 19|VDD \$313 \$314 19|VDD sg13_lv_pmos L=0.5u W=1u AS=0.1523p AD=0.34p
+ PS=1.38u PD=2.68u
M$6957 19|VDD \$314 \$326 19|VDD sg13_lv_pmos L=0.5u W=1u AS=0.2254p AD=0.34p
+ PS=1.53u PD=2.68u
M$6958 19|VDD \$326 A|X$12 19|VDD sg13_lv_pmos L=0.13u W=1.12u AS=0.2254p
+ AD=0.4256p PS=1.53u PD=3u
M$6959 19|VDD A|B|Y A|Y$4 19|VDD sg13_lv_pmos L=0.13u W=8.96u AS=1.876p
+ AD=1.876p PS=13.43u PD=13.43u
M$6967 \$336 \$335 19|VDD 19|VDD sg13_lv_pmos L=0.5u W=1u AS=0.34p AD=0.2254p
+ PS=2.68u PD=1.53u
M$6968 19|VDD \$336 A|X$10 19|VDD sg13_lv_pmos L=0.13u W=1.12u AS=0.2254p
+ AD=0.4256p PS=1.53u PD=3u
M$6969 19|VDD A|X$10 \$297 19|VDD sg13_lv_pmos L=0.13u W=0.42u AS=0.1523p
+ AD=0.1428p PS=1.38u PD=1.52u
M$6970 19|VDD \$297 \$298 19|VDD sg13_lv_pmos L=0.5u W=1u AS=0.1523p AD=0.34p
+ PS=1.38u PD=2.68u
M$6971 19|VDD A|X$8 \$317 19|VDD sg13_lv_pmos L=0.13u W=0.42u AS=0.1523p
+ AD=0.1428p PS=1.38u PD=1.52u
M$6972 19|VDD \$317 \$318 19|VDD sg13_lv_pmos L=0.5u W=1u AS=0.1523p AD=0.34p
+ PS=1.38u PD=2.68u
M$6973 19|VDD \$318 \$327 19|VDD sg13_lv_pmos L=0.5u W=1u AS=0.2254p AD=0.34p
+ PS=1.53u PD=2.68u
M$6974 19|VDD \$327 A|X$13 19|VDD sg13_lv_pmos L=0.13u W=1.12u AS=0.2254p
+ AD=0.4256p PS=1.53u PD=3u
M$6975 19|VDD A|Y$9 \$348 19|VDD sg13_lv_pmos L=0.13u W=1.12u AS=0.4032p
+ AD=0.1176p PS=2.96u PD=1.33u
M$6976 \$348 B|X A|B|Y$1 19|VDD sg13_lv_pmos L=0.13u W=1.12u AS=0.1176p
+ AD=0.3808p PS=1.33u PD=2.92u
M$6977 19|VDD A|X$13 \$320 19|VDD sg13_lv_pmos L=0.13u W=0.42u AS=0.1523p
+ AD=0.1428p PS=1.38u PD=1.52u
M$6978 19|VDD \$320 \$321 19|VDD sg13_lv_pmos L=0.5u W=1u AS=0.1523p AD=0.34p
+ PS=1.38u PD=2.68u
M$6979 19|VDD A|X$9 \$347 19|VDD sg13_lv_pmos L=0.13u W=1.12u AS=0.4032p
+ AD=0.1176p PS=2.96u PD=1.33u
M$6980 \$347 A|B|Y$1 A|Y$9 19|VDD sg13_lv_pmos L=0.13u W=1.12u AS=0.1176p
+ AD=0.3808p PS=1.33u PD=2.92u
M$6981 19|VDD \$321 \$328 19|VDD sg13_lv_pmos L=0.5u W=1u AS=0.2254p AD=0.34p
+ PS=1.53u PD=2.68u
M$6982 19|VDD \$328 A|X$11 19|VDD sg13_lv_pmos L=0.13u W=1.12u AS=0.2254p
+ AD=0.4256p PS=1.53u PD=3u
M$6983 19|VDD A|B|Y$2 A|Y$3 19|VDD sg13_lv_pmos L=0.13u W=1.12u AS=0.392p
+ AD=0.392p PS=2.94u PD=2.94u
M$6984 19|VDD A|Y$5 \$338 19|VDD sg13_lv_pmos L=0.13u W=0.84u AS=0.2856p
+ AD=0.1596p PS=2.36u PD=1.22u
M$6985 19|VDD A|B|Y$2 \$338 19|VDD sg13_lv_pmos L=0.13u W=0.84u AS=0.1918p
+ AD=0.1596p PS=1.5u PD=1.22u
M$6986 19|VDD \$338 X 19|VDD sg13_lv_pmos L=0.13u W=2.24u AS=0.4046p AD=0.6384p
+ PS=3u PD=4.5u
M$6988 19|VDD A|X$11 A|B|Y$2 19|VDD sg13_lv_pmos L=0.13u W=1.12u AS=0.392p
+ AD=0.392p PS=2.94u PD=2.94u
M$6989 19|VDD A|B|Y A|Y$5 19|VDD sg13_lv_pmos L=0.13u W=1.12u AS=0.392p
+ AD=0.392p PS=2.94u PD=2.94u
M$6990 19|VDD A|Y$7 \$340 19|VDD sg13_lv_pmos L=0.13u W=0.84u AS=0.2856p
+ AD=0.1596p PS=2.36u PD=1.22u
M$6991 19|VDD A|B|Y$3 \$340 19|VDD sg13_lv_pmos L=0.13u W=0.84u AS=0.1918p
+ AD=0.1596p PS=1.5u PD=1.22u
M$6992 19|VDD \$340 B|X 19|VDD sg13_lv_pmos L=0.13u W=2.24u AS=0.4046p
+ AD=0.6384p PS=3u PD=4.5u
M$6994 19|VDD A|B|Y$3 A|Y$6 19|VDD sg13_lv_pmos L=0.13u W=1.12u AS=0.392p
+ AD=0.392p PS=2.94u PD=2.94u
M$6995 19|VDD A|B|Y$4 A|Y$7 19|VDD sg13_lv_pmos L=0.13u W=1.12u AS=0.392p
+ AD=0.392p PS=2.94u PD=2.94u
M$6996 19|VDD A|Y$6 \$341 19|VDD sg13_lv_pmos L=0.13u W=0.84u AS=0.2856p
+ AD=0.1596p PS=2.36u PD=1.22u
M$6997 19|VDD A|B|Y$4 \$341 19|VDD sg13_lv_pmos L=0.13u W=0.84u AS=0.1918p
+ AD=0.1596p PS=1.5u PD=1.22u
M$6998 19|VDD \$341 X 19|VDD sg13_lv_pmos L=0.13u W=2.24u AS=0.4046p AD=0.6384p
+ PS=3u PD=4.5u
M$7000 19|VDD A|Y$8 A|B|Y$3 19|VDD sg13_lv_pmos L=0.13u W=1.12u AS=0.392p
+ AD=0.392p PS=2.94u PD=2.94u
M$7001 19|VDD A|VINS|X A|Y$8 19|VDD sg13_lv_pmos L=0.13u W=2.24u AS=0.5964p
+ AD=0.5964p PS=4.425u PD=4.425u
M$7003 \$325 A|VINS|X 19|VDD 19|VDD sg13_lv_pmos L=0.13u W=0.84u AS=0.3024p
+ AD=0.2051p PS=2.4u PD=1.52u
M$7004 19|VDD \$325 A$4 19|VDD sg13_lv_pmos L=0.13u W=1.12u AS=0.2051p
+ AD=0.4032p PS=1.52u PD=2.96u
M$7005 19|VDD A$5 \$333 19|VDD sg13_lv_pmos L=0.13u W=1.68u AS=0.3626p
+ AD=0.4452p PS=2.72u PD=3.58u
M$7007 19|VDD \$333 A|X$7 19|VDD sg13_lv_pmos L=0.13u W=4.48u AS=1.0192p
+ AD=0.8414p PS=7.42u PD=6u
M$7011 19|VDD \$349 18|NOC_P_BUFF|X 19|VDD sg13_lv_pmos L=0.13u W=17.92u
+ AS=3.5896p AD=3.4048p PS=25.45u PD=24u
M$7027 19|VDD A|X$14 \$349 19|VDD sg13_lv_pmos L=0.13u W=6.72u AS=1.2768p
+ AD=1.4448p PS=9u PD=10.42u
M$7033 19|VDD A|X$12 \$334 19|VDD sg13_lv_pmos L=0.13u W=0.42u AS=0.1523p
+ AD=0.1428p PS=1.38u PD=1.52u
M$7034 19|VDD \$334 \$335 19|VDD sg13_lv_pmos L=0.5u W=1u AS=0.1523p AD=0.34p
+ PS=1.38u PD=2.68u
M$7035 19|VDD A|B|Y$3 A|Y$10 19|VDD sg13_lv_pmos L=0.13u W=8.96u AS=1.876p
+ AD=1.876p PS=13.43u PD=13.43u
M$7043 19|VDD A|X$15 A|B|Y$4 19|VDD sg13_lv_pmos L=0.13u W=1.12u AS=0.392p
+ AD=0.392p PS=2.94u PD=2.94u
M$7044 19|VDD A|X$16 \$352 19|VDD sg13_lv_pmos L=0.13u W=0.42u AS=0.1523p
+ AD=0.1428p PS=1.38u PD=1.52u
M$7045 19|VDD \$352 \$353 19|VDD sg13_lv_pmos L=0.5u W=1u AS=0.1523p AD=0.34p
+ PS=1.38u PD=2.68u
M$7046 19|VDD \$353 \$354 19|VDD sg13_lv_pmos L=0.5u W=1u AS=0.2254p AD=0.34p
+ PS=1.53u PD=2.68u
M$7047 19|VDD \$354 A|X$15 19|VDD sg13_lv_pmos L=0.13u W=1.12u AS=0.2254p
+ AD=0.4256p PS=1.53u PD=3u
M$7048 \$351 NOC_N|X 19|VDD 19|VDD sg13_lv_pmos L=0.13u W=0.84u AS=0.3024p
+ AD=0.2051p PS=2.4u PD=1.52u
M$7049 19|VDD \$351 A$5 19|VDD sg13_lv_pmos L=0.13u W=1.12u AS=0.2051p
+ AD=0.4032p PS=1.52u PD=2.96u
M$7050 19|VDD \$358 18|NOC_P_BUFF|X 19|VDD sg13_lv_pmos L=0.13u W=17.92u
+ AS=3.5896p AD=3.4048p PS=25.45u PD=24u
M$7066 19|VDD A|X$14 \$358 19|VDD sg13_lv_pmos L=0.13u W=6.72u AS=1.2768p
+ AD=1.4448p PS=9u PD=10.42u
M$7072 19|VDD A|Y$10 \$359 19|VDD sg13_lv_pmos L=0.13u W=0.42u AS=0.1523p
+ AD=0.1428p PS=1.38u PD=1.52u
M$7073 19|VDD \$359 \$360 19|VDD sg13_lv_pmos L=0.5u W=1u AS=0.1523p AD=0.34p
+ PS=1.38u PD=2.68u
M$7074 \$368 \$360 19|VDD 19|VDD sg13_lv_pmos L=0.5u W=1u AS=0.34p AD=0.2254p
+ PS=2.68u PD=1.53u
M$7075 19|VDD \$368 A|X$17 19|VDD sg13_lv_pmos L=0.13u W=1.12u AS=0.2254p
+ AD=0.4256p PS=1.53u PD=3u
M$7076 19|VDD A|X$17 \$362 19|VDD sg13_lv_pmos L=0.13u W=0.42u AS=0.1523p
+ AD=0.1428p PS=1.38u PD=1.52u
M$7077 19|VDD \$362 \$363 19|VDD sg13_lv_pmos L=0.5u W=1u AS=0.1523p AD=0.34p
+ PS=1.38u PD=2.68u
M$7078 \$369 \$363 19|VDD 19|VDD sg13_lv_pmos L=0.5u W=1u AS=0.34p AD=0.2254p
+ PS=2.68u PD=1.53u
M$7079 19|VDD \$369 A|X$18 19|VDD sg13_lv_pmos L=0.13u W=1.12u AS=0.2254p
+ AD=0.4256p PS=1.53u PD=3u
M$7080 19|VDD A|X$18 \$365 19|VDD sg13_lv_pmos L=0.13u W=0.42u AS=0.1523p
+ AD=0.1428p PS=1.38u PD=1.52u
M$7081 19|VDD \$365 \$366 19|VDD sg13_lv_pmos L=0.5u W=1u AS=0.1523p AD=0.34p
+ PS=1.38u PD=2.68u
M$7082 \$370 \$366 19|VDD 19|VDD sg13_lv_pmos L=0.5u W=1u AS=0.34p AD=0.2254p
+ PS=2.68u PD=1.53u
M$7083 19|VDD \$370 A|X$19 19|VDD sg13_lv_pmos L=0.13u W=1.12u AS=0.2254p
+ AD=0.4256p PS=1.53u PD=3u
M$7084 19|VDD \$372 18|NOC_P_BUFF|X 19|VDD sg13_lv_pmos L=0.13u W=17.92u
+ AS=3.5896p AD=3.4048p PS=25.45u PD=24u
M$7100 19|VDD A|X$14 \$372 19|VDD sg13_lv_pmos L=0.13u W=6.72u AS=1.2768p
+ AD=1.4448p PS=9u PD=10.42u
M$7106 19|VDD \$381 18|NOC_P_BUFF|X 19|VDD sg13_lv_pmos L=0.13u W=17.92u
+ AS=3.5896p AD=3.4048p PS=25.45u PD=24u
M$7122 19|VDD A|X$14 \$381 19|VDD sg13_lv_pmos L=0.13u W=6.72u AS=1.2768p
+ AD=1.4448p PS=9u PD=10.42u
M$7128 19|VDD \$382 A|X$14 19|VDD sg13_lv_pmos L=0.13u W=17.92u AS=3.5896p
+ AD=3.4048p PS=25.45u PD=24u
M$7144 19|VDD A|X$20 \$382 19|VDD sg13_lv_pmos L=0.13u W=6.72u AS=1.2768p
+ AD=1.4448p PS=9u PD=10.42u
M$7150 19|VDD A$6 \$384 19|VDD sg13_lv_pmos L=0.13u W=1.68u AS=0.3626p
+ AD=0.4452p PS=2.72u PD=3.58u
M$7152 19|VDD \$384 A|X$20 19|VDD sg13_lv_pmos L=0.13u W=4.48u AS=1.0192p
+ AD=0.8414p PS=7.42u PD=6u
M$7156 \$387 \$386 19|VDD 19|VDD sg13_lv_pmos L=0.5u W=1u AS=0.34p AD=0.2254p
+ PS=2.68u PD=1.53u
M$7157 19|VDD \$387 A|X$21 19|VDD sg13_lv_pmos L=0.13u W=1.12u AS=0.2254p
+ AD=0.4256p PS=1.53u PD=3u
M$7158 \$391 \$390 19|VDD 19|VDD sg13_lv_pmos L=0.5u W=1u AS=0.34p AD=0.2254p
+ PS=2.68u PD=1.53u
M$7159 19|VDD \$391 A|X$22 19|VDD sg13_lv_pmos L=0.13u W=1.12u AS=0.2254p
+ AD=0.4256p PS=1.53u PD=3u
M$7160 \$395 \$394 19|VDD 19|VDD sg13_lv_pmos L=0.5u W=1u AS=0.34p AD=0.2254p
+ PS=2.68u PD=1.53u
M$7161 19|VDD \$395 A|X$23 19|VDD sg13_lv_pmos L=0.13u W=1.12u AS=0.2254p
+ AD=0.4256p PS=1.53u PD=3u
M$7162 \$399 \$398 19|VDD 19|VDD sg13_lv_pmos L=0.5u W=1u AS=0.34p AD=0.2254p
+ PS=2.68u PD=1.53u
M$7163 19|VDD \$399 A|X$24 19|VDD sg13_lv_pmos L=0.13u W=1.12u AS=0.2254p
+ AD=0.4256p PS=1.53u PD=3u
M$7164 19|VDD A|X$19 \$375 19|VDD sg13_lv_pmos L=0.13u W=0.42u AS=0.1523p
+ AD=0.1428p PS=1.38u PD=1.52u
M$7165 19|VDD \$375 \$376 19|VDD sg13_lv_pmos L=0.5u W=1u AS=0.1523p AD=0.34p
+ PS=1.38u PD=2.68u
M$7166 19|VDD \$376 \$379 19|VDD sg13_lv_pmos L=0.5u W=1u AS=0.2254p AD=0.34p
+ PS=1.53u PD=2.68u
M$7167 19|VDD \$379 A|X$16 19|VDD sg13_lv_pmos L=0.13u W=1.12u AS=0.2254p
+ AD=0.4256p PS=1.53u PD=3u
M$7168 19|VDD A|X$28 \$416 19|VDD sg13_lv_pmos L=0.13u W=0.42u AS=0.1523p
+ AD=0.1428p PS=1.38u PD=1.52u
M$7169 19|VDD \$416 \$418 19|VDD sg13_lv_pmos L=0.5u W=1u AS=0.1523p AD=0.34p
+ PS=1.38u PD=2.68u
M$7170 \$419 \$418 19|VDD 19|VDD sg13_lv_pmos L=0.5u W=1u AS=0.34p AD=0.2254p
+ PS=2.68u PD=1.53u
M$7171 19|VDD \$419 A|X$29 19|VDD sg13_lv_pmos L=0.13u W=1.12u AS=0.2254p
+ AD=0.4256p PS=1.53u PD=3u
M$7172 19|VDD A|Y$12 \$421 19|VDD sg13_lv_pmos L=0.13u W=0.42u AS=0.1523p
+ AD=0.1428p PS=1.38u PD=1.52u
M$7173 19|VDD \$421 \$423 19|VDD sg13_lv_pmos L=0.5u W=1u AS=0.1523p AD=0.34p
+ PS=1.38u PD=2.68u
M$7174 \$424 \$423 19|VDD 19|VDD sg13_lv_pmos L=0.5u W=1u AS=0.34p AD=0.2254p
+ PS=2.68u PD=1.53u
M$7175 19|VDD \$424 A|X$30 19|VDD sg13_lv_pmos L=0.13u W=1.12u AS=0.2254p
+ AD=0.4256p PS=1.53u PD=3u
M$7176 19|VDD A|X$31 \$426 19|VDD sg13_lv_pmos L=0.13u W=0.42u AS=0.1523p
+ AD=0.1428p PS=1.38u PD=1.52u
M$7177 19|VDD \$426 \$428 19|VDD sg13_lv_pmos L=0.5u W=1u AS=0.1523p AD=0.34p
+ PS=1.38u PD=2.68u
M$7178 \$429 \$428 19|VDD 19|VDD sg13_lv_pmos L=0.5u W=1u AS=0.34p AD=0.2254p
+ PS=2.68u PD=1.53u
M$7179 19|VDD \$429 A|X$32 19|VDD sg13_lv_pmos L=0.13u W=1.12u AS=0.2254p
+ AD=0.4256p PS=1.53u PD=3u
M$7180 19|VDD A|X$33 \$431 19|VDD sg13_lv_pmos L=0.13u W=0.42u AS=0.1523p
+ AD=0.1428p PS=1.38u PD=1.52u
M$7181 19|VDD \$431 \$433 19|VDD sg13_lv_pmos L=0.5u W=1u AS=0.1523p AD=0.34p
+ PS=1.38u PD=2.68u
M$7182 \$434 \$433 19|VDD 19|VDD sg13_lv_pmos L=0.5u W=1u AS=0.34p AD=0.2254p
+ PS=2.68u PD=1.53u
M$7183 19|VDD \$434 A|X$34 19|VDD sg13_lv_pmos L=0.13u W=1.12u AS=0.2254p
+ AD=0.4256p PS=1.53u PD=3u
M$7184 19|VDD A|Y$11 \$436 19|VDD sg13_lv_pmos L=0.13u W=0.42u AS=0.1523p
+ AD=0.1428p PS=1.38u PD=1.52u
M$7185 19|VDD \$436 \$437 19|VDD sg13_lv_pmos L=0.5u W=1u AS=0.1523p AD=0.34p
+ PS=1.38u PD=2.68u
M$7186 \$438 \$437 19|VDD 19|VDD sg13_lv_pmos L=0.5u W=1u AS=0.34p AD=0.2254p
+ PS=2.68u PD=1.53u
M$7187 19|VDD \$438 A|X$35 19|VDD sg13_lv_pmos L=0.13u W=1.12u AS=0.2254p
+ AD=0.4256p PS=1.53u PD=3u
M$7188 19|VDD A|Y$11 \$403 19|VDD sg13_lv_pmos L=0.13u W=0.42u AS=0.1523p
+ AD=0.1428p PS=1.38u PD=1.52u
M$7189 19|VDD \$403 \$404 19|VDD sg13_lv_pmos L=0.5u W=1u AS=0.1523p AD=0.34p
+ PS=1.38u PD=2.68u
M$7190 19|VDD \$404 \$411 19|VDD sg13_lv_pmos L=0.5u W=1u AS=0.2254p AD=0.34p
+ PS=1.53u PD=2.68u
M$7191 19|VDD \$411 A|X$25 19|VDD sg13_lv_pmos L=0.13u W=1.12u AS=0.2254p
+ AD=0.4256p PS=1.53u PD=3u
M$7192 19|VDD A|X$36 \$457 19|VDD sg13_lv_pmos L=0.13u W=1.12u AS=0.4032p
+ AD=0.1176p PS=2.96u PD=1.33u
M$7193 \$457 A|B|Y$1 A|Y$11 19|VDD sg13_lv_pmos L=0.13u W=1.12u AS=0.1176p
+ AD=0.3808p PS=1.33u PD=2.92u
M$7194 19|VDD A|X$25 \$385 19|VDD sg13_lv_pmos L=0.13u W=0.42u AS=0.1523p
+ AD=0.1428p PS=1.38u PD=1.52u
M$7195 19|VDD \$385 \$386 19|VDD sg13_lv_pmos L=0.5u W=1u AS=0.1523p AD=0.34p
+ PS=1.38u PD=2.68u
M$7196 19|VDD A|X$36 A|Y$13 19|VDD sg13_lv_pmos L=0.13u W=2.24u AS=0.5964p
+ AD=0.5964p PS=4.425u PD=4.425u
M$7198 19|VDD A|Y$14 \$456 19|VDD sg13_lv_pmos L=0.13u W=1.12u AS=0.4032p
+ AD=0.1176p PS=2.96u PD=1.33u
M$7199 \$456 A|B|X A|Y$12 19|VDD sg13_lv_pmos L=0.13u W=1.12u AS=0.1176p
+ AD=0.3808p PS=1.33u PD=2.92u
M$7200 19|VDD A|X$21 \$389 19|VDD sg13_lv_pmos L=0.13u W=0.42u AS=0.1523p
+ AD=0.1428p PS=1.38u PD=1.52u
M$7201 19|VDD \$389 \$390 19|VDD sg13_lv_pmos L=0.5u W=1u AS=0.1523p AD=0.34p
+ PS=1.38u PD=2.68u
M$7202 19|VDD A|B|Y$1 A|Y$14 19|VDD sg13_lv_pmos L=0.13u W=1.12u AS=0.392p
+ AD=0.392p PS=2.94u PD=2.94u
M$7203 19|VDD NOC_P|X \$444 19|VDD sg13_lv_pmos L=0.13u W=0.84u AS=0.2051p
+ AD=0.3024p PS=1.52u PD=2.4u
M$7204 19|VDD \$444 A$6 19|VDD sg13_lv_pmos L=0.13u W=1.12u AS=0.2051p
+ AD=0.4032p PS=1.52u PD=2.96u
M$7205 19|VDD A|X$22 \$393 19|VDD sg13_lv_pmos L=0.13u W=0.42u AS=0.1523p
+ AD=0.1428p PS=1.38u PD=1.52u
M$7206 19|VDD \$393 \$394 19|VDD sg13_lv_pmos L=0.5u W=1u AS=0.1523p AD=0.34p
+ PS=1.38u PD=2.68u
M$7207 19|VDD A|Y$15 A0|Y 19|VDD sg13_lv_pmos L=0.13u W=4.48u AS=1.0192p
+ AD=1.0192p PS=7.42u PD=7.42u
M$7211 19|VDD A|X$23 \$397 19|VDD sg13_lv_pmos L=0.13u W=0.42u AS=0.1523p
+ AD=0.1428p PS=1.38u PD=1.52u
M$7212 19|VDD \$397 \$398 19|VDD sg13_lv_pmos L=0.5u W=1u AS=0.1523p AD=0.34p
+ PS=1.38u PD=2.68u
M$7213 19|VDD A|B|X A|Y$16 19|VDD sg13_lv_pmos L=0.13u W=1.12u AS=0.392p
+ AD=0.392p PS=2.94u PD=2.94u
M$7214 19|VDD A|X$24 \$405 19|VDD sg13_lv_pmos L=0.13u W=0.42u AS=0.1523p
+ AD=0.1428p PS=1.38u PD=1.52u
M$7215 19|VDD \$405 \$406 19|VDD sg13_lv_pmos L=0.5u W=1u AS=0.1523p AD=0.34p
+ PS=1.38u PD=2.68u
M$7216 19|VDD \$406 \$412 19|VDD sg13_lv_pmos L=0.5u W=1u AS=0.2254p AD=0.34p
+ PS=1.53u PD=2.68u
M$7217 19|VDD \$412 A|X$26 19|VDD sg13_lv_pmos L=0.13u W=1.12u AS=0.2254p
+ AD=0.4256p PS=1.53u PD=3u
M$7218 19|VDD A|X$26 \$408 19|VDD sg13_lv_pmos L=0.13u W=0.42u AS=0.1523p
+ AD=0.1428p PS=1.38u PD=1.52u
M$7219 19|VDD \$408 \$409 19|VDD sg13_lv_pmos L=0.5u W=1u AS=0.1523p AD=0.34p
+ PS=1.38u PD=2.68u
M$7220 19|VDD A|X$27 \$447 19|VDD sg13_lv_pmos L=0.13u W=0.42u AS=0.1523p
+ AD=0.1428p PS=1.38u PD=1.52u
M$7221 19|VDD \$447 \$448 19|VDD sg13_lv_pmos L=0.5u W=1u AS=0.1523p AD=0.34p
+ PS=1.38u PD=2.68u
M$7222 19|VDD \$409 \$413 19|VDD sg13_lv_pmos L=0.5u W=1u AS=0.2254p AD=0.34p
+ PS=1.53u PD=2.68u
M$7223 19|VDD \$413 A|X$27 19|VDD sg13_lv_pmos L=0.13u W=1.12u AS=0.2254p
+ AD=0.4256p PS=1.53u PD=3u
M$7224 \$449 \$448 19|VDD 19|VDD sg13_lv_pmos L=0.5u W=1u AS=0.34p AD=0.2254p
+ PS=2.68u PD=1.53u
M$7225 19|VDD \$449 A|X$37 19|VDD sg13_lv_pmos L=0.13u W=1.12u AS=0.2254p
+ AD=0.4256p PS=1.53u PD=3u
M$7226 19|VDD A|X$37 \$451 19|VDD sg13_lv_pmos L=0.13u W=0.42u AS=0.1523p
+ AD=0.1428p PS=1.38u PD=1.52u
M$7227 19|VDD \$451 \$452 19|VDD sg13_lv_pmos L=0.5u W=1u AS=0.1523p AD=0.34p
+ PS=1.38u PD=2.68u
M$7228 \$453 \$452 19|VDD 19|VDD sg13_lv_pmos L=0.5u W=1u AS=0.34p AD=0.2254p
+ PS=2.68u PD=1.53u
M$7229 19|VDD \$453 A|X$38 19|VDD sg13_lv_pmos L=0.13u W=1.12u AS=0.2254p
+ AD=0.4256p PS=1.53u PD=3u
M$7230 19|VDD A|Y$12 \$458 19|VDD sg13_lv_pmos L=0.13u W=0.42u AS=0.1523p
+ AD=0.1428p PS=1.38u PD=1.52u
M$7231 19|VDD \$458 \$459 19|VDD sg13_lv_pmos L=0.5u W=1u AS=0.1523p AD=0.34p
+ PS=1.38u PD=2.68u
M$7232 19|VDD \$459 \$490 19|VDD sg13_lv_pmos L=0.5u W=1u AS=0.2254p AD=0.34p
+ PS=1.53u PD=2.68u
M$7233 19|VDD \$490 A|X$39 19|VDD sg13_lv_pmos L=0.13u W=1.12u AS=0.2254p
+ AD=0.4256p PS=1.53u PD=3u
M$7234 19|VDD A|X$46 \$461 19|VDD sg13_lv_pmos L=0.13u W=0.42u AS=0.1523p
+ AD=0.1428p PS=1.38u PD=1.52u
M$7235 19|VDD \$461 \$462 19|VDD sg13_lv_pmos L=0.5u W=1u AS=0.1523p AD=0.34p
+ PS=1.38u PD=2.68u
M$7236 19|VDD \$462 \$492 19|VDD sg13_lv_pmos L=0.5u W=1u AS=0.2254p AD=0.34p
+ PS=1.53u PD=2.68u
M$7237 19|VDD \$492 A|X$40 19|VDD sg13_lv_pmos L=0.13u W=1.12u AS=0.2254p
+ AD=0.4256p PS=1.53u PD=3u
M$7238 19|VDD A|X$30 \$464 19|VDD sg13_lv_pmos L=0.13u W=0.42u AS=0.1523p
+ AD=0.1428p PS=1.38u PD=1.52u
M$7239 19|VDD \$464 \$465 19|VDD sg13_lv_pmos L=0.5u W=1u AS=0.1523p AD=0.34p
+ PS=1.38u PD=2.68u
M$7240 19|VDD \$465 \$493 19|VDD sg13_lv_pmos L=0.5u W=1u AS=0.2254p AD=0.34p
+ PS=1.53u PD=2.68u
M$7241 19|VDD \$493 A|X$41 19|VDD sg13_lv_pmos L=0.13u W=1.12u AS=0.2254p
+ AD=0.4256p PS=1.53u PD=3u
M$7242 19|VDD A|X$32 \$467 19|VDD sg13_lv_pmos L=0.13u W=0.42u AS=0.1523p
+ AD=0.1428p PS=1.38u PD=1.52u
M$7243 19|VDD \$467 \$468 19|VDD sg13_lv_pmos L=0.5u W=1u AS=0.1523p AD=0.34p
+ PS=1.38u PD=2.68u
M$7244 19|VDD \$468 \$494 19|VDD sg13_lv_pmos L=0.5u W=1u AS=0.2254p AD=0.34p
+ PS=1.53u PD=2.68u
M$7245 19|VDD \$494 A|X$42 19|VDD sg13_lv_pmos L=0.13u W=1.12u AS=0.2254p
+ AD=0.4256p PS=1.53u PD=3u
M$7246 19|VDD A|X$42 \$470 19|VDD sg13_lv_pmos L=0.13u W=0.42u AS=0.1523p
+ AD=0.1428p PS=1.38u PD=1.52u
M$7247 19|VDD \$470 \$471 19|VDD sg13_lv_pmos L=0.5u W=1u AS=0.1523p AD=0.34p
+ PS=1.38u PD=2.68u
M$7248 19|VDD \$471 \$495 19|VDD sg13_lv_pmos L=0.5u W=1u AS=0.2254p AD=0.34p
+ PS=1.53u PD=2.68u
M$7249 19|VDD \$495 A|X$43 19|VDD sg13_lv_pmos L=0.13u W=1.12u AS=0.2254p
+ AD=0.4256p PS=1.53u PD=3u
M$7250 19|VDD A|X$34 \$473 19|VDD sg13_lv_pmos L=0.13u W=0.42u AS=0.1523p
+ AD=0.1428p PS=1.38u PD=1.52u
M$7251 19|VDD \$473 \$474 19|VDD sg13_lv_pmos L=0.5u W=1u AS=0.1523p AD=0.34p
+ PS=1.38u PD=2.68u
M$7252 19|VDD \$474 \$496 19|VDD sg13_lv_pmos L=0.5u W=1u AS=0.2254p AD=0.34p
+ PS=1.53u PD=2.68u
M$7253 19|VDD \$496 A0|X 19|VDD sg13_lv_pmos L=0.13u W=1.12u AS=0.2254p
+ AD=0.4256p PS=1.53u PD=3u
M$7254 19|VDD A|X$35 \$476 19|VDD sg13_lv_pmos L=0.13u W=0.42u AS=0.1523p
+ AD=0.1428p PS=1.38u PD=1.52u
M$7255 19|VDD \$476 \$477 19|VDD sg13_lv_pmos L=0.5u W=1u AS=0.1523p AD=0.34p
+ PS=1.38u PD=2.68u
M$7256 19|VDD \$477 \$497 19|VDD sg13_lv_pmos L=0.5u W=1u AS=0.2254p AD=0.34p
+ PS=1.53u PD=2.68u
M$7257 19|VDD \$497 A|X$44 19|VDD sg13_lv_pmos L=0.13u W=1.12u AS=0.2254p
+ AD=0.4256p PS=1.53u PD=3u
M$7258 19|VDD A|X$44 \$479 19|VDD sg13_lv_pmos L=0.13u W=0.42u AS=0.1523p
+ AD=0.1428p PS=1.38u PD=1.52u
M$7259 19|VDD \$479 \$480 19|VDD sg13_lv_pmos L=0.5u W=1u AS=0.1523p AD=0.34p
+ PS=1.38u PD=2.68u
M$7260 19|VDD \$480 \$498 19|VDD sg13_lv_pmos L=0.5u W=1u AS=0.2254p AD=0.34p
+ PS=1.53u PD=2.68u
M$7261 19|VDD \$498 A|X$45 19|VDD sg13_lv_pmos L=0.13u W=1.12u AS=0.2254p
+ AD=0.4256p PS=1.53u PD=3u
M$7262 19|VDD A|Y$13 A0|Y$1 19|VDD sg13_lv_pmos L=0.13u W=4.48u AS=1.0192p
+ AD=1.0192p PS=7.42u PD=7.42u
M$7266 19|VDD A|X$38 \$487 19|VDD sg13_lv_pmos L=0.13u W=0.42u AS=0.1523p
+ AD=0.1428p PS=1.38u PD=1.52u
M$7267 19|VDD \$487 \$488 19|VDD sg13_lv_pmos L=0.5u W=1u AS=0.1523p AD=0.34p
+ PS=1.38u PD=2.68u
M$7268 19|VDD \$488 \$499 19|VDD sg13_lv_pmos L=0.5u W=1u AS=0.2254p AD=0.34p
+ PS=1.53u PD=2.68u
M$7269 19|VDD \$499 A1|X 19|VDD sg13_lv_pmos L=0.13u W=1.12u AS=0.2254p
+ AD=0.4256p PS=1.53u PD=3u
M$7270 \$511 \$510 19|VDD 19|VDD sg13_lv_pmos L=0.5u W=1u AS=0.34p AD=0.2254p
+ PS=2.68u PD=1.53u
M$7271 19|VDD \$511 A|X$28 19|VDD sg13_lv_pmos L=0.13u W=1.12u AS=0.2254p
+ AD=0.4256p PS=1.53u PD=3u
M$7272 \$514 \$513 19|VDD 19|VDD sg13_lv_pmos L=0.5u W=1u AS=0.34p AD=0.2254p
+ PS=2.68u PD=1.53u
M$7273 19|VDD \$514 A|X$46 19|VDD sg13_lv_pmos L=0.13u W=1.12u AS=0.2254p
+ AD=0.4256p PS=1.53u PD=3u
M$7274 \$517 \$516 19|VDD 19|VDD sg13_lv_pmos L=0.5u W=1u AS=0.34p AD=0.2254p
+ PS=2.68u PD=1.53u
M$7275 19|VDD \$517 A|X$31 19|VDD sg13_lv_pmos L=0.13u W=1.12u AS=0.2254p
+ AD=0.4256p PS=1.53u PD=3u
M$7276 \$520 \$519 19|VDD 19|VDD sg13_lv_pmos L=0.5u W=1u AS=0.34p AD=0.2254p
+ PS=2.68u PD=1.53u
M$7277 19|VDD \$520 A|X$33 19|VDD sg13_lv_pmos L=0.13u W=1.12u AS=0.2254p
+ AD=0.4256p PS=1.53u PD=3u
M$7278 \$523 \$522 19|VDD 19|VDD sg13_lv_pmos L=0.5u W=1u AS=0.34p AD=0.2254p
+ PS=2.68u PD=1.53u
M$7279 19|VDD \$523 A1|X$1 19|VDD sg13_lv_pmos L=0.13u W=1.12u AS=0.2254p
+ AD=0.4256p PS=1.53u PD=3u
M$7280 \$525 13|S|VSEL_DT 19|VDD 19|VDD sg13_lv_pmos L=0.13u W=0.84u AS=0.2856p
+ AD=0.253p PS=2.36u PD=1.53u
M$7281 19|VDD 13|S|VSEL_DT \$543 19|VDD sg13_lv_pmos L=0.13u W=1u AS=0.253p
+ AD=0.3325p PS=1.53u PD=1.665u
M$7282 \$543 A0|X \$526 19|VDD sg13_lv_pmos L=0.13u W=1u AS=0.3325p AD=0.2225p
+ PS=1.665u PD=1.445u
M$7283 \$526 A1|X$1 \$542 19|VDD sg13_lv_pmos L=0.13u W=1u AS=0.2225p
+ AD=0.2975p PS=1.445u PD=1.595u
M$7284 \$542 \$525 19|VDD 19|VDD sg13_lv_pmos L=0.13u W=1u AS=0.2975p
+ AD=0.2198p PS=1.595u PD=1.52u
M$7285 19|VDD \$526 A|X$36 19|VDD sg13_lv_pmos L=0.13u W=2.24u AS=0.5278p
+ AD=0.784p PS=3.19u PD=4.76u
M$7287 \$529 \$528 19|VDD 19|VDD sg13_lv_pmos L=0.5u W=1u AS=0.34p AD=0.2254p
+ PS=2.68u PD=1.53u
M$7288 19|VDD \$529 A|X$47 19|VDD sg13_lv_pmos L=0.13u W=1.12u AS=0.2254p
+ AD=0.4256p PS=1.53u PD=3u
M$7289 \$531 13|S|VSEL_DT 19|VDD 19|VDD sg13_lv_pmos L=0.13u W=0.84u AS=0.2856p
+ AD=0.253p PS=2.36u PD=1.53u
M$7290 19|VDD 13|S|VSEL_DT \$541 19|VDD sg13_lv_pmos L=0.13u W=1u AS=0.253p
+ AD=0.3325p PS=1.53u PD=1.665u
M$7291 \$541 A0|X$1 \$532 19|VDD sg13_lv_pmos L=0.13u W=1u AS=0.3325p
+ AD=0.2225p PS=1.665u PD=1.445u
M$7292 \$532 A1|X \$540 19|VDD sg13_lv_pmos L=0.13u W=1u AS=0.2225p AD=0.2975p
+ PS=1.445u PD=1.595u
M$7293 \$540 \$531 19|VDD 19|VDD sg13_lv_pmos L=0.13u W=1u AS=0.2975p
+ AD=0.2198p PS=1.595u PD=1.52u
M$7294 19|VDD \$532 A|B|X 19|VDD sg13_lv_pmos L=0.13u W=2.24u AS=0.5278p
+ AD=0.784p PS=3.19u PD=4.76u
M$7296 19|VDD 12|S|VSEL_OL \$483 19|VDD sg13_lv_pmos L=0.13u W=0.84u AS=0.253p
+ AD=0.2856p PS=1.53u PD=2.36u
M$7297 19|VDD 12|S|VSEL_OL \$504 19|VDD sg13_lv_pmos L=0.13u W=1u AS=0.253p
+ AD=0.3325p PS=1.53u PD=1.665u
M$7298 \$504 A0|Y$1 \$484 19|VDD sg13_lv_pmos L=0.13u W=1u AS=0.3325p
+ AD=0.2225p PS=1.665u PD=1.445u
M$7299 \$484 11|A1|VINR_OL \$503 19|VDD sg13_lv_pmos L=0.13u W=1u AS=0.2225p
+ AD=0.2975p PS=1.445u PD=1.595u
M$7300 19|VDD \$483 \$503 19|VDD sg13_lv_pmos L=0.13u W=1u AS=0.2198p
+ AD=0.2975p PS=1.52u PD=1.595u
M$7301 19|VDD \$484 NOC_N|X 19|VDD sg13_lv_pmos L=0.13u W=2.24u AS=0.5278p
+ AD=0.784p PS=3.19u PD=4.76u
M$7303 19|VDD A|Y$16 A|Y$15 19|VDD sg13_lv_pmos L=0.13u W=2.24u AS=0.5964p
+ AD=0.5964p PS=4.425u PD=4.425u
M$7305 19|VDD 12|S|VSEL_OL \$485 19|VDD sg13_lv_pmos L=0.13u W=0.84u AS=0.253p
+ AD=0.2856p PS=1.53u PD=2.36u
M$7306 19|VDD 12|S|VSEL_OL \$502 19|VDD sg13_lv_pmos L=0.13u W=1u AS=0.253p
+ AD=0.3325p PS=1.53u PD=1.665u
M$7307 \$502 A0|Y \$486 19|VDD sg13_lv_pmos L=0.13u W=1u AS=0.3325p AD=0.2225p
+ PS=1.665u PD=1.445u
M$7308 \$486 10|A1|VINS_OL \$501 19|VDD sg13_lv_pmos L=0.13u W=1u AS=0.2225p
+ AD=0.2975p PS=1.445u PD=1.595u
M$7309 19|VDD \$485 \$501 19|VDD sg13_lv_pmos L=0.13u W=1u AS=0.2198p
+ AD=0.2975p PS=1.52u PD=1.595u
M$7310 19|VDD \$486 NOC_P|X 19|VDD sg13_lv_pmos L=0.13u W=2.24u AS=0.5278p
+ AD=0.784p PS=3.19u PD=4.76u
M$7312 19|VDD A|X$39 \$509 19|VDD sg13_lv_pmos L=0.13u W=0.42u AS=0.1523p
+ AD=0.1428p PS=1.38u PD=1.52u
M$7313 19|VDD \$509 \$510 19|VDD sg13_lv_pmos L=0.5u W=1u AS=0.1523p AD=0.34p
+ PS=1.38u PD=2.68u
M$7314 19|VDD A|X$29 \$512 19|VDD sg13_lv_pmos L=0.13u W=0.42u AS=0.1523p
+ AD=0.1428p PS=1.38u PD=1.52u
M$7315 19|VDD \$512 \$513 19|VDD sg13_lv_pmos L=0.5u W=1u AS=0.1523p AD=0.34p
+ PS=1.38u PD=2.68u
M$7316 19|VDD A|X$40 \$515 19|VDD sg13_lv_pmos L=0.13u W=0.42u AS=0.1523p
+ AD=0.1428p PS=1.38u PD=1.52u
M$7317 19|VDD \$515 \$516 19|VDD sg13_lv_pmos L=0.5u W=1u AS=0.1523p AD=0.34p
+ PS=1.38u PD=2.68u
M$7318 19|VDD A|X$41 \$518 19|VDD sg13_lv_pmos L=0.13u W=0.42u AS=0.1523p
+ AD=0.1428p PS=1.38u PD=1.52u
M$7319 19|VDD \$518 \$519 19|VDD sg13_lv_pmos L=0.5u W=1u AS=0.1523p AD=0.34p
+ PS=1.38u PD=2.68u
M$7320 19|VDD A|X$43 \$521 19|VDD sg13_lv_pmos L=0.13u W=0.42u AS=0.1523p
+ AD=0.1428p PS=1.38u PD=1.52u
M$7321 19|VDD \$521 \$522 19|VDD sg13_lv_pmos L=0.5u W=1u AS=0.1523p AD=0.34p
+ PS=1.38u PD=2.68u
M$7322 19|VDD A|X$45 \$527 19|VDD sg13_lv_pmos L=0.13u W=0.42u AS=0.1523p
+ AD=0.1428p PS=1.38u PD=1.52u
M$7323 19|VDD \$527 \$528 19|VDD sg13_lv_pmos L=0.5u W=1u AS=0.1523p AD=0.34p
+ PS=1.38u PD=2.68u
M$7324 19|VDD A|X$47 \$544 19|VDD sg13_lv_pmos L=0.13u W=0.42u AS=0.1523p
+ AD=0.1428p PS=1.38u PD=1.52u
M$7325 19|VDD \$544 \$545 19|VDD sg13_lv_pmos L=0.5u W=1u AS=0.1523p AD=0.34p
+ PS=1.38u PD=2.68u
M$7326 19|VDD \$545 \$546 19|VDD sg13_lv_pmos L=0.5u W=1u AS=0.2254p AD=0.34p
+ PS=1.53u PD=2.68u
M$7327 19|VDD \$546 A0|X$1 19|VDD sg13_lv_pmos L=0.13u W=1.12u AS=0.2254p
+ AD=0.4256p PS=1.53u PD=3u
M$7328 \$572 NOC_P|X 19|VDD 19|VDD sg13_lv_pmos L=0.13u W=2.24u AS=1.0528p
+ AD=1.0528p PS=5.24u PD=5.24u
M$7330 \$574 NOC_N|X 19|VDD 19|VDD sg13_lv_pmos L=0.13u W=2.24u AS=1.0528p
+ AD=1.0528p PS=5.24u PD=5.24u
M$7332 9 9 9 9 sg13_hv_pmos L=0.45u W=24u AS=7.04p AD=7.04p PS=42.08u PD=42.08u
M$7333 9 \$81 8 9 sg13_hv_pmos L=0.45u W=64u AS=16p AD=16p PS=96u PD=96u
M$7366 9 \$82 \$81 9 sg13_hv_pmos L=0.45u W=32u AS=8p AD=8p PS=48u PD=48u
M$7383 9 \$83 \$82 9 sg13_hv_pmos L=0.45u W=16u AS=4p AD=4p PS=24u PD=24u
M$7392 9 \$84 \$83 9 sg13_hv_pmos L=0.45u W=8u AS=2p AD=2p PS=12u PD=12u
M$7397 9 \$85 \$84 9 sg13_hv_pmos L=0.45u W=4u AS=1p AD=1p PS=6u PD=6u
M$7471 9 \$86 \$85 9 sg13_hv_pmos L=0.45u W=2u AS=0.5p AD=0.5p PS=3u PD=3u
M$7474 1 1 1 1 sg13_hv_pmos L=0.45u W=24u AS=7.04p AD=7.04p PS=42.08u PD=42.08u
M$7478 1 \$102 \$103 1 sg13_hv_pmos L=0.45u W=4u AS=1p AD=1p PS=6u PD=6u
M$7481 1 \$103 \$104 1 sg13_hv_pmos L=0.45u W=8u AS=2p AD=2p PS=12u PD=12u
M$7486 1 \$104 \$106 1 sg13_hv_pmos L=0.45u W=16u AS=4p AD=4p PS=24u PD=24u
M$7495 1 \$106 \$107 1 sg13_hv_pmos L=0.45u W=32u AS=8p AD=8p PS=48u PD=48u
M$7512 1 \$107 7 1 sg13_hv_pmos L=0.45u W=64u AS=16p AD=16p PS=96u PD=96u
M$7546 1 \$93 \$102 1 sg13_hv_pmos L=0.45u W=2u AS=0.5p AD=0.5p PS=3u PD=3u
M$7616 9 9 9 9 sg13_hv_pmos L=7u W=33.6u AS=26.2374p AD=26.2374p PS=183.54u
+ PD=183.54u
M$7617 9 9 \$140 9 sg13_hv_pmos L=7u W=4.8u AS=2.3868p AD=2.3868p PS=16.92u
+ PD=16.92u
M$7621 9 2 \$141 9 sg13_hv_pmos L=7u W=3.6u AS=1.7901p AD=1.7901p PS=12.69u
+ PD=12.69u
M$7625 9 2 \$142 9 sg13_hv_pmos L=7u W=3.6u AS=1.7901p AD=1.7901p PS=12.69u
+ PD=12.69u
M$7629 9 2 \$143 9 sg13_hv_pmos L=7u W=3.6u AS=1.7901p AD=1.7901p PS=12.69u
+ PD=12.69u
M$7633 9 2 \$144 9 sg13_hv_pmos L=7u W=3.6u AS=1.7901p AD=1.7901p PS=12.69u
+ PD=12.69u
M$7637 9 2 \$145 9 sg13_hv_pmos L=7u W=3.6u AS=1.7901p AD=1.7901p PS=12.69u
+ PD=12.69u
M$7641 9 9 \$146 9 sg13_hv_pmos L=7u W=4.8u AS=2.3868p AD=2.3868p PS=16.92u
+ PD=16.92u
M$7678 \$141 9 9 9 sg13_hv_pmos L=7u W=0.8u AS=0.3978p AD=0.3978p PS=2.82u
+ PD=2.82u
M$7682 \$142 9 9 9 sg13_hv_pmos L=7u W=0.8u AS=0.3978p AD=0.3978p PS=2.82u
+ PD=2.82u
M$7686 \$143 9 9 9 sg13_hv_pmos L=7u W=0.8u AS=0.3978p AD=0.3978p PS=2.82u
+ PD=2.82u
M$7690 \$144 9 9 9 sg13_hv_pmos L=7u W=0.8u AS=0.3978p AD=0.3978p PS=2.82u
+ PD=2.82u
M$7694 \$145 9 9 9 sg13_hv_pmos L=7u W=0.8u AS=0.3978p AD=0.3978p PS=2.82u
+ PD=2.82u
M$7706 \$141 6 9 9 sg13_hv_pmos L=7u W=0.4u AS=0.1989p AD=0.1989p PS=1.41u
+ PD=1.41u
M$7710 \$142 6 9 9 sg13_hv_pmos L=7u W=0.4u AS=0.1989p AD=0.1989p PS=1.41u
+ PD=1.41u
M$7714 \$143 4 9 9 sg13_hv_pmos L=7u W=0.4u AS=0.1989p AD=0.1989p PS=1.41u
+ PD=1.41u
M$7718 \$144 4 9 9 sg13_hv_pmos L=7u W=0.4u AS=0.1989p AD=0.1989p PS=1.41u
+ PD=1.41u
M$7722 \$145 6 9 9 sg13_hv_pmos L=7u W=0.4u AS=0.1989p AD=0.1989p PS=1.41u
+ PD=1.41u
M$7756 9 9 9 9 sg13_hv_pmos L=4u W=49u AS=17.71p AD=15.89p PS=105.42u PD=94.78u
M$7757 9 \$150 \$150 9 sg13_hv_pmos L=4u W=8u AS=2p AD=2p PS=12u PD=12u
M$7768 9 \$151 \$151 9 sg13_hv_pmos L=4u W=8u AS=2p AD=2p PS=12u PD=12u
M$7779 9 \$152 \$152 9 sg13_hv_pmos L=4u W=8u AS=2p AD=2p PS=12u PD=12u
M$7790 9 \$153 \$153 9 sg13_hv_pmos L=4u W=8u AS=2p AD=2p PS=12u PD=12u
M$7801 9 \$154 \$154 9 sg13_hv_pmos L=4u W=8u AS=2p AD=2p PS=12u PD=12u
M$7812 9 \$155 \$155 9 sg13_hv_pmos L=4u W=8u AS=2p AD=2p PS=12u PD=12u
M$7823 9 \$156 \$156 9 sg13_hv_pmos L=4u W=8u AS=2p AD=2p PS=12u PD=12u
M$7834 9 \$150 \$157 9 sg13_hv_pmos L=4u W=5u AS=1.25p AD=1.25p PS=7.5u PD=7.5u
M$7839 \$157 9 9 9 sg13_hv_pmos L=4u W=1u AS=0.25p AD=0.51p PS=1.5u PD=3.02u
M$7841 9 \$151 \$158 9 sg13_hv_pmos L=4u W=5u AS=1.25p AD=1.25p PS=7.5u PD=7.5u
M$7846 \$158 9 9 9 sg13_hv_pmos L=4u W=1u AS=0.25p AD=0.51p PS=1.5u PD=3.02u
M$7848 9 \$152 \$159 9 sg13_hv_pmos L=4u W=5u AS=1.25p AD=1.25p PS=7.5u PD=7.5u
M$7853 \$159 9 9 9 sg13_hv_pmos L=4u W=1u AS=0.25p AD=0.51p PS=1.5u PD=3.02u
M$7855 9 \$153 \$160 9 sg13_hv_pmos L=4u W=5u AS=1.25p AD=1.25p PS=7.5u PD=7.5u
M$7860 \$160 9 9 9 sg13_hv_pmos L=4u W=1u AS=0.25p AD=0.51p PS=1.5u PD=3.02u
M$7862 9 \$154 \$161 9 sg13_hv_pmos L=4u W=5u AS=1.25p AD=1.25p PS=7.5u PD=7.5u
M$7867 \$161 9 9 9 sg13_hv_pmos L=4u W=1u AS=0.25p AD=0.51p PS=1.5u PD=3.02u
M$7869 9 \$155 \$162 9 sg13_hv_pmos L=4u W=5u AS=1.25p AD=1.25p PS=7.5u PD=7.5u
M$7874 \$162 9 9 9 sg13_hv_pmos L=4u W=1u AS=0.25p AD=0.51p PS=1.5u PD=3.02u
M$7876 9 \$156 \$163 9 sg13_hv_pmos L=4u W=5u AS=1.25p AD=1.25p PS=7.5u PD=7.5u
M$7881 \$163 9 9 9 sg13_hv_pmos L=4u W=1u AS=0.25p AD=0.51p PS=1.5u PD=3.02u
M$7931 9 9 \$157 9 sg13_hv_pmos L=5u W=5u AS=2.55p AD=1.25p PS=11.02u PD=5.5u
M$7932 \$157 6 \$164 9 sg13_hv_pmos L=5u W=5u AS=1.25p AD=1.25p PS=5.5u PD=5.5u
M$7933 \$164 9 9 9 sg13_hv_pmos L=5u W=5u AS=1.25p AD=2.55p PS=5.5u PD=11.02u
M$7934 9 9 \$158 9 sg13_hv_pmos L=5u W=5u AS=2.55p AD=1.25p PS=11.02u PD=5.5u
M$7935 \$158 \$170 \$165 9 sg13_hv_pmos L=5u W=5u AS=1.25p AD=1.25p PS=5.5u
+ PD=5.5u
M$7936 \$165 9 9 9 sg13_hv_pmos L=5u W=5u AS=1.25p AD=2.55p PS=5.5u PD=11.02u
M$7937 9 9 \$159 9 sg13_hv_pmos L=5u W=5u AS=2.55p AD=1.25p PS=11.02u PD=5.5u
M$7938 \$159 \$165 \$166 9 sg13_hv_pmos L=5u W=5u AS=1.25p AD=1.25p PS=5.5u
+ PD=5.5u
M$7939 \$166 9 9 9 sg13_hv_pmos L=5u W=5u AS=1.25p AD=2.55p PS=5.5u PD=11.02u
M$7940 9 9 \$160 9 sg13_hv_pmos L=5u W=5u AS=2.55p AD=1.25p PS=11.02u PD=5.5u
M$7941 \$160 \$166 \$167 9 sg13_hv_pmos L=5u W=5u AS=1.25p AD=1.25p PS=5.5u
+ PD=5.5u
M$7942 \$167 9 9 9 sg13_hv_pmos L=5u W=5u AS=1.25p AD=2.55p PS=5.5u PD=11.02u
M$7943 9 9 \$161 9 sg13_hv_pmos L=5u W=5u AS=2.55p AD=1.25p PS=11.02u PD=5.5u
M$7944 \$161 \$167 \$168 9 sg13_hv_pmos L=5u W=5u AS=1.25p AD=1.25p PS=5.5u
+ PD=5.5u
M$7945 \$168 9 9 9 sg13_hv_pmos L=5u W=5u AS=1.25p AD=2.55p PS=5.5u PD=11.02u
M$7947 9 \$168 \$184 9 sg13_hv_pmos L=0.45u W=2u AS=0.5p AD=0.5p PS=3u PD=3u
M$7950 9 \$184 \$86 9 sg13_hv_pmos L=0.45u W=4u AS=1p AD=1p PS=6u PD=6u
M$7954 1 \$194 \$195 1 sg13_hv_pmos L=0.45u W=2u AS=0.5p AD=0.5p PS=3u PD=3u
M$7957 1 \$195 \$93 1 sg13_hv_pmos L=0.45u W=4u AS=1p AD=1p PS=6u PD=6u
M$7974 9 9 \$162 9 sg13_hv_pmos L=5u W=5u AS=2.55p AD=1.25p PS=11.02u PD=5.5u
M$7975 \$162 \$168 \$170 9 sg13_hv_pmos L=5u W=5u AS=1.25p AD=1.25p PS=5.5u
+ PD=5.5u
M$7976 \$170 9 9 9 sg13_hv_pmos L=5u W=5u AS=1.25p AD=2.55p PS=5.5u PD=11.02u
M$7977 9 9 \$163 9 sg13_hv_pmos L=5u W=5u AS=2.55p AD=1.25p PS=11.02u PD=5.5u
M$7978 \$163 6 \$169 9 sg13_hv_pmos L=5u W=5u AS=1.25p AD=1.25p PS=5.5u PD=5.5u
M$7979 \$169 9 9 9 sg13_hv_pmos L=5u W=5u AS=1.25p AD=2.55p PS=5.5u PD=11.02u
M$7980 A \$93 19|VDD 19|VDD sg13_hv_pmos L=0.4u W=2u AS=1.12p AD=1.12p PS=5.24u
+ PD=5.24u
M$7982 A$1 \$86 19|VDD 19|VDD sg13_hv_pmos L=0.4u W=2u AS=1.12p AD=1.12p
+ PS=5.24u PD=5.24u
M$7984 1 1 \$250 1 sg13_hv_pmos L=5u W=5u AS=2.55p AD=1.25p PS=11.02u PD=5.5u
M$7985 \$250 5 \$236 1 sg13_hv_pmos L=5u W=5u AS=1.25p AD=1.25p PS=5.5u PD=5.5u
M$7986 \$236 1 1 1 sg13_hv_pmos L=5u W=5u AS=1.25p AD=2.55p PS=5.5u PD=11.02u
M$7987 1 1 \$251 1 sg13_hv_pmos L=5u W=5u AS=2.55p AD=1.25p PS=11.02u PD=5.5u
M$7988 \$251 \$199 \$238 1 sg13_hv_pmos L=5u W=5u AS=1.25p AD=1.25p PS=5.5u
+ PD=5.5u
M$7989 \$238 1 1 1 sg13_hv_pmos L=5u W=5u AS=1.25p AD=2.55p PS=5.5u PD=11.02u
M$7990 1 1 \$252 1 sg13_hv_pmos L=5u W=5u AS=2.55p AD=1.25p PS=11.02u PD=5.5u
M$7991 \$252 \$238 \$239 1 sg13_hv_pmos L=5u W=5u AS=1.25p AD=1.25p PS=5.5u
+ PD=5.5u
M$7992 \$239 1 1 1 sg13_hv_pmos L=5u W=5u AS=1.25p AD=2.55p PS=5.5u PD=11.02u
M$7993 1 1 \$253 1 sg13_hv_pmos L=5u W=5u AS=2.55p AD=1.25p PS=11.02u PD=5.5u
M$7994 \$253 \$239 \$240 1 sg13_hv_pmos L=5u W=5u AS=1.25p AD=1.25p PS=5.5u
+ PD=5.5u
M$7995 \$240 1 1 1 sg13_hv_pmos L=5u W=5u AS=1.25p AD=2.55p PS=5.5u PD=11.02u
M$7996 1 1 \$254 1 sg13_hv_pmos L=5u W=5u AS=2.55p AD=1.25p PS=11.02u PD=5.5u
M$7997 \$254 \$240 \$194 1 sg13_hv_pmos L=5u W=5u AS=1.25p AD=1.25p PS=5.5u
+ PD=5.5u
M$7998 \$194 1 1 1 sg13_hv_pmos L=5u W=5u AS=1.25p AD=2.55p PS=5.5u PD=11.02u
M$7999 1 1 \$255 1 sg13_hv_pmos L=5u W=5u AS=2.55p AD=1.25p PS=11.02u PD=5.5u
M$8000 \$255 \$194 \$199 1 sg13_hv_pmos L=5u W=5u AS=1.25p AD=1.25p PS=5.5u
+ PD=5.5u
M$8001 \$199 1 1 1 sg13_hv_pmos L=5u W=5u AS=1.25p AD=2.55p PS=5.5u PD=11.02u
M$8002 1 1 \$256 1 sg13_hv_pmos L=5u W=5u AS=2.55p AD=1.25p PS=11.02u PD=5.5u
M$8003 \$256 5 \$237 1 sg13_hv_pmos L=5u W=5u AS=1.25p AD=1.25p PS=5.5u PD=5.5u
M$8004 \$237 1 1 1 sg13_hv_pmos L=5u W=5u AS=1.25p AD=2.55p PS=5.5u PD=11.02u
M$8005 1 1 1 1 sg13_hv_pmos L=4u W=49u AS=17.71p AD=15.89p PS=105.42u PD=94.78u
M$8006 1 \$224 \$224 1 sg13_hv_pmos L=4u W=8u AS=2p AD=2p PS=12u PD=12u
M$8013 1 \$225 \$225 1 sg13_hv_pmos L=4u W=8u AS=2p AD=2p PS=12u PD=12u
M$8020 1 \$226 \$226 1 sg13_hv_pmos L=4u W=8u AS=2p AD=2p PS=12u PD=12u
M$8027 1 \$227 \$227 1 sg13_hv_pmos L=4u W=8u AS=2p AD=2p PS=12u PD=12u
M$8034 1 \$228 \$228 1 sg13_hv_pmos L=4u W=8u AS=2p AD=2p PS=12u PD=12u
M$8041 1 \$229 \$229 1 sg13_hv_pmos L=4u W=8u AS=2p AD=2p PS=12u PD=12u
M$8048 1 \$230 \$230 1 sg13_hv_pmos L=4u W=8u AS=2p AD=2p PS=12u PD=12u
M$8055 1 \$224 \$250 1 sg13_hv_pmos L=4u W=5u AS=1.25p AD=1.25p PS=7.5u PD=7.5u
M$8060 \$250 1 1 1 sg13_hv_pmos L=4u W=1u AS=0.25p AD=0.51p PS=1.5u PD=3.02u
M$8062 1 \$225 \$251 1 sg13_hv_pmos L=4u W=5u AS=1.25p AD=1.25p PS=7.5u PD=7.5u
M$8067 \$251 1 1 1 sg13_hv_pmos L=4u W=1u AS=0.25p AD=0.51p PS=1.5u PD=3.02u
M$8069 1 \$226 \$252 1 sg13_hv_pmos L=4u W=5u AS=1.25p AD=1.25p PS=7.5u PD=7.5u
M$8074 \$252 1 1 1 sg13_hv_pmos L=4u W=1u AS=0.25p AD=0.51p PS=1.5u PD=3.02u
M$8076 1 \$227 \$253 1 sg13_hv_pmos L=4u W=5u AS=1.25p AD=1.25p PS=7.5u PD=7.5u
M$8081 \$253 1 1 1 sg13_hv_pmos L=4u W=1u AS=0.25p AD=0.51p PS=1.5u PD=3.02u
M$8083 1 \$228 \$254 1 sg13_hv_pmos L=4u W=5u AS=1.25p AD=1.25p PS=7.5u PD=7.5u
M$8088 \$254 1 1 1 sg13_hv_pmos L=4u W=1u AS=0.25p AD=0.51p PS=1.5u PD=3.02u
M$8090 1 \$229 \$255 1 sg13_hv_pmos L=4u W=5u AS=1.25p AD=1.25p PS=7.5u PD=7.5u
M$8095 \$255 1 1 1 sg13_hv_pmos L=4u W=1u AS=0.25p AD=0.51p PS=1.5u PD=3.02u
M$8097 1 \$230 \$256 1 sg13_hv_pmos L=4u W=5u AS=1.25p AD=1.25p PS=7.5u PD=7.5u
M$8102 \$256 1 1 1 sg13_hv_pmos L=4u W=1u AS=0.25p AD=0.51p PS=1.5u PD=3.02u
M$8152 1 1 1 1 sg13_hv_pmos L=7u W=33.6u AS=26.2374p AD=26.2374p PS=183.54u
+ PD=183.54u
M$8153 1 1 \$204 1 sg13_hv_pmos L=7u W=4.8u AS=2.3868p AD=2.3868p PS=16.92u
+ PD=16.92u
M$8161 1 2 \$205 1 sg13_hv_pmos L=7u W=3.6u AS=1.7901p AD=1.7901p PS=12.69u
+ PD=12.69u
M$8169 1 2 \$206 1 sg13_hv_pmos L=7u W=3.6u AS=1.7901p AD=1.7901p PS=12.69u
+ PD=12.69u
M$8177 1 2 \$207 1 sg13_hv_pmos L=7u W=3.6u AS=1.7901p AD=1.7901p PS=12.69u
+ PD=12.69u
M$8185 1 2 \$208 1 sg13_hv_pmos L=7u W=3.6u AS=1.7901p AD=1.7901p PS=12.69u
+ PD=12.69u
M$8193 1 2 \$209 1 sg13_hv_pmos L=7u W=3.6u AS=1.7901p AD=1.7901p PS=12.69u
+ PD=12.69u
M$8201 1 1 \$210 1 sg13_hv_pmos L=7u W=4.8u AS=2.3868p AD=2.3868p PS=16.92u
+ PD=16.92u
M$8213 1 1 \$205 1 sg13_hv_pmos L=7u W=0.8u AS=0.3978p AD=0.3978p PS=2.82u
+ PD=2.82u
M$8214 \$205 5 1 1 sg13_hv_pmos L=7u W=0.4u AS=0.1989p AD=0.1989p PS=1.41u
+ PD=1.41u
M$8217 1 1 \$206 1 sg13_hv_pmos L=7u W=0.8u AS=0.3978p AD=0.3978p PS=2.82u
+ PD=2.82u
M$8218 \$206 5 1 1 sg13_hv_pmos L=7u W=0.4u AS=0.1989p AD=0.1989p PS=1.41u
+ PD=1.41u
M$8221 1 1 \$207 1 sg13_hv_pmos L=7u W=0.8u AS=0.3978p AD=0.3978p PS=2.82u
+ PD=2.82u
M$8222 \$207 3 1 1 sg13_hv_pmos L=7u W=0.4u AS=0.1989p AD=0.1989p PS=1.41u
+ PD=1.41u
M$8225 1 1 \$208 1 sg13_hv_pmos L=7u W=0.8u AS=0.3978p AD=0.3978p PS=2.82u
+ PD=2.82u
M$8226 \$208 3 1 1 sg13_hv_pmos L=7u W=0.4u AS=0.1989p AD=0.1989p PS=1.41u
+ PD=1.41u
M$8229 1 1 \$209 1 sg13_hv_pmos L=7u W=0.8u AS=0.3978p AD=0.3978p PS=2.82u
+ PD=2.82u
M$8230 \$209 5 1 1 sg13_hv_pmos L=7u W=0.4u AS=0.1989p AD=0.1989p PS=1.41u
+ PD=1.41u
M$8320 27 \$414 28 28 sg13_hv_pmos L=0.4u W=120960u AS=44217.6p AD=44217.6p
+ PS=134283.52u PD=134283.52u
M$11722 \$414 \$563 23 23 sg13_hv_pmos L=0.4u W=2500u AS=638p AD=638p
+ PS=2677.6u PD=2677.6u
M$11772 23 23 23 23 sg13_hv_pmos L=0.4u W=280u AS=75.2p AD=75.2p PS=315.04u
+ PD=315.04u
M$11775 23 23 \$563 23 sg13_hv_pmos L=0.4u W=20u AS=5p AD=5p PS=21u PD=21u
M$11776 \$563 \$567 23 23 sg13_hv_pmos L=0.4u W=300u AS=75p AD=75p PS=315u
+ PD=315u
M$11808 23 23 \$567 23 sg13_hv_pmos L=0.4u W=10u AS=2.5p AD=2.5p PS=10.5u
+ PD=10.5u
M$11809 \$567 \$568 23 23 sg13_hv_pmos L=0.4u W=10u AS=2.5p AD=2.5p PS=10.5u
+ PD=10.5u
M$11818 23 23 \$568 23 sg13_hv_pmos L=0.4u W=10u AS=2.5p AD=2.5p PS=10.5u
+ PD=10.5u
M$11819 \$568 \$567 23 23 sg13_hv_pmos L=0.4u W=10u AS=2.5p AD=2.5p PS=10.5u
+ PD=10.5u
M$11822 \$562 \$564 23 23 sg13_hv_pmos L=0.4u W=2500u AS=638p AD=638p
+ PS=2677.6u PD=2677.6u
M$11875 23 23 \$564 23 sg13_hv_pmos L=0.4u W=20u AS=5p AD=5p PS=21u PD=21u
M$11876 \$564 \$569 23 23 sg13_hv_pmos L=0.4u W=300u AS=75p AD=75p PS=315u
+ PD=315u
M$11908 23 23 \$569 23 sg13_hv_pmos L=0.4u W=10u AS=2.5p AD=2.5p PS=10.5u
+ PD=10.5u
M$11909 \$569 \$570 23 23 sg13_hv_pmos L=0.4u W=10u AS=2.5p AD=2.5p PS=10.5u
+ PD=10.5u
M$11918 23 23 \$570 23 sg13_hv_pmos L=0.4u W=10u AS=2.5p AD=2.5p PS=10.5u
+ PD=10.5u
M$11919 \$570 \$569 23 23 sg13_hv_pmos L=0.4u W=10u AS=2.5p AD=2.5p PS=10.5u
+ PD=10.5u
M$19504 23 23 23 23 sg13_hv_pmos L=0.45u W=32u AS=9.04p AD=9.04p PS=54.08u
+ PD=54.08u
M$19505 23 \$623 21 23 sg13_hv_pmos L=0.45u W=64u AS=16p AD=16p PS=96u PD=96u
M$19538 23 \$627 \$623 23 sg13_hv_pmos L=0.45u W=32u AS=8p AD=8p PS=48u PD=48u
M$19555 23 \$634 \$627 23 sg13_hv_pmos L=0.45u W=16u AS=4p AD=4p PS=24u PD=24u
M$19564 23 \$635 \$634 23 sg13_hv_pmos L=0.45u W=8u AS=2p AD=2p PS=12u PD=12u
M$19569 23 \$637 \$635 23 sg13_hv_pmos L=0.45u W=4u AS=1p AD=1p PS=6u PD=6u
M$19572 23 \$562 \$637 23 sg13_hv_pmos L=0.45u W=2u AS=0.5p AD=0.5p PS=3u PD=3u
M$21162 23 \$651 \$652 23 sg13_hv_pmos L=0.45u W=4u AS=1p AD=1p PS=6u PD=6u
M$21165 23 \$652 \$653 23 sg13_hv_pmos L=0.45u W=8u AS=2p AD=2p PS=12u PD=12u
M$21170 23 \$653 \$654 23 sg13_hv_pmos L=0.45u W=16u AS=4p AD=4p PS=24u PD=24u
M$21179 23 \$654 \$655 23 sg13_hv_pmos L=0.45u W=32u AS=8p AD=8p PS=48u PD=48u
M$21196 23 \$655 22 23 sg13_hv_pmos L=0.45u W=64u AS=16p AD=16p PS=96u PD=96u
M$21230 23 \$414 \$651 23 sg13_hv_pmos L=0.45u W=2u AS=0.5p AD=0.5p PS=3u PD=3u
D$21300 15|25|VSS 24 8 diodevdd_2kv m=1
D$21301 15|25|VSS 24 9 diodevdd_2kv m=1
D$21302 15|25|VSS 24 10|A1|VINS_OL diodevdd_2kv m=1
D$21303 15|25|VSS 24 11|A1|VINR_OL diodevdd_2kv m=1
D$21304 15|25|VSS 24 12|S|VSEL_OL diodevdd_2kv m=1
D$21305 15|25|VSS 24 13|S|VSEL_DT diodevdd_2kv m=1
D$21306 15|25|VSS 24 14|VINR_BUFF|X diodevdd_2kv m=1
D$21307 15|25|VSS 24 7 diodevdd_2kv m=1
D$21308 15|25|VSS 24 15|25|VSS diodevdd_2kv m=2
D$21309 15|25|VSS 24 6 diodevdd_2kv m=1
D$21310 15|25|VSS 24 16|PD_BUFF|X diodevdd_2kv m=1
D$21311 15|25|VSS 24 5 diodevdd_2kv m=1
D$21312 15|25|VSS 24 17|NOC_N_BUFF|X diodevdd_2kv m=1
D$21313 15|25|VSS 24 4 diodevdd_2kv m=1
D$21314 15|25|VSS 24 18|NOC_P_BUFF|X diodevdd_2kv m=1
D$21315 15|25|VSS 24 3 diodevdd_2kv m=1
D$21316 15|25|VSS 24 19|VDD diodevdd_2kv m=1
D$21317 15|25|VSS 24 2 diodevdd_2kv m=1
D$21318 15|25|VSS 24 20 diodevdd_2kv m=1
D$21319 15|25|VSS 24 1 diodevdd_2kv m=1
D$21320 15|25|VSS 24 21 diodevdd_2kv m=1
D$21321 15|25|VSS 24 28 diodevdd_2kv m=1
D$21322 15|25|VSS 24 27 diodevdd_2kv m=1
D$21323 15|25|VSS 24 26 diodevdd_2kv m=1
D$21325 15|25|VSS 24 24 diodevdd_2kv m=1
D$21326 15|25|VSS 24 23 diodevdd_2kv m=1
D$21327 15|25|VSS 24 22 diodevdd_2kv m=1
D$21328 24 15|25|VSS 8 diodevss_2kv m=1
D$21329 24 15|25|VSS 9 diodevss_2kv m=1
D$21330 24 15|25|VSS 10|A1|VINS_OL diodevss_2kv m=1
D$21331 24 15|25|VSS 11|A1|VINR_OL diodevss_2kv m=1
D$21332 24 15|25|VSS 12|S|VSEL_OL diodevss_2kv m=1
D$21333 24 15|25|VSS 13|S|VSEL_DT diodevss_2kv m=1
D$21334 24 15|25|VSS 14|VINR_BUFF|X diodevss_2kv m=1
D$21335 24 15|25|VSS 7 diodevss_2kv m=1
D$21336 24 15|25|VSS 15|25|VSS diodevss_2kv m=2
D$21337 24 15|25|VSS 6 diodevss_2kv m=1
D$21338 24 15|25|VSS 16|PD_BUFF|X diodevss_2kv m=1
D$21339 24 15|25|VSS 5 diodevss_2kv m=1
D$21340 24 15|25|VSS 17|NOC_N_BUFF|X diodevss_2kv m=1
D$21341 24 15|25|VSS 4 diodevss_2kv m=1
D$21342 24 15|25|VSS 18|NOC_P_BUFF|X diodevss_2kv m=1
D$21343 24 15|25|VSS 3 diodevss_2kv m=1
D$21344 24 15|25|VSS 19|VDD diodevss_2kv m=1
D$21345 24 15|25|VSS 2 diodevss_2kv m=1
D$21346 24 15|25|VSS 20 diodevss_2kv m=1
D$21347 24 15|25|VSS 1 diodevss_2kv m=1
D$21348 24 15|25|VSS 21 diodevss_2kv m=1
D$21349 24 15|25|VSS 28 diodevss_2kv m=1
D$21350 24 15|25|VSS 27 diodevss_2kv m=1
D$21351 24 15|25|VSS 26 diodevss_2kv m=1
D$21353 24 15|25|VSS 24 diodevss_2kv m=1
D$21354 24 15|25|VSS 23 diodevss_2kv m=1
D$21355 24 15|25|VSS 22 diodevss_2kv m=1
.ENDS top
