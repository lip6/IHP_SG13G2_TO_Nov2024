* testlib


* Device subcircuits
*
.subckt rsil n1 n2 l=1e-6 w=1e-6
.param rsil_res={l*7.0/w}
Rres n1 n2 r={rsil_res} rsil l=l w=w
.ends rsil

.subckt rppd n1 n2 l=1e-6 w=1e-6
.param rppd_res={l*260.0/w}
Rres n1 n2 r={rppd_res} rppd l=l w=w
.ends rppd

.subckt dantenna an cat params: w=0.48e-6 l=0.48e-6
Ddio an cat dantenna a=(w*l) p=(2*(w + l))
.ends dantenna

.subckt dpantenna an cat params: w=0.48e-6 l=0.48e-6
Ddio an cat dpantenna a=(w*l) p=(2*(w + l))
.ends dpantenna

.subckt sg13_lv_nmos s g d b params: l=0.13e-6 w=0.15e-6
Mtrans s g d b sg13_lv_nmos l=l w=w
.ends sg13_lv_nmos

.subckt sg13_lv_pmos s g d b params: l=0.13e-6 w=0.15e-6
Mtrans s g d b sg13_lv_pmos l=l w=w
.ends sg13_lv_pmos

.subckt sg13_hv_nmos s g d b params: l=0.45e-6 w=0.3e-6
Mtrans s g d b sg13_hv_nmos l=l w=w
.ends sg13_hv_nmos

.subckt sg13_hv_pmos s g d b params: l=0.45e-6 w=0.3e-6
Mtrans s g d b sg13_hv_pmos l=l w=w
.ends sg13_hv_pmos

* Library cells
*
.subckt BondPad PAD
.ends BondPad

.subckt SP6TVar0Cell wl bl bl_n vdd vss
Xpu1 vdd bit_n bit vdd sg13_lv_pmos l=1.3e-07 w=3e-07
Xpd1 bit bit_n vss vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpu2 vdd bit bit_n vdd sg13_lv_pmos l=1.3e-07 w=3e-07
Xpd2 bit_n bit vss vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg1 bit wl bl vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg2 bit_n wl bl_n vss sg13_lv_nmos l=1.3e-07 w=3e-07
.ends SP6TVar0Cell

.subckt SP6TVar0Array_2X1 vss vdd wl[0] wl[1] bl[0] bl_n[0]
Xinst0x0 wl[0] bl[0] bl_n[0] vdd vss SP6TVar0Cell
Xinst1x0 wl[1] bl[0] bl_n[0] vdd vss SP6TVar0Cell
.ends SP6TVar0Array_2X1

.subckt SP6TVar0Array_2X2 vss vdd wl[0] wl[1] bl[0] bl_n[0] bl[1] bl_n[1]
Xinst0x0 vss vdd wl[0] wl[1] bl[0] bl_n[0] SP6TVar0Array_2X1
Xinst0x1 vss vdd wl[0] wl[1] bl[1] bl_n[1] SP6TVar0Array_2X1
.ends SP6TVar0Array_2X2

.subckt SP6TVar0Array_4X2 vss vdd wl[0] wl[1] wl[2] wl[3] bl[0] bl_n[0] bl[1] bl_n[1]
Xinst0x0 vss vdd wl[0] wl[1] bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar0Array_2X2
Xinst1x0 vss vdd wl[2] wl[3] bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar0Array_2X2
.ends SP6TVar0Array_4X2

.subckt SP6TVar0Array_4X4 vss vdd wl[0] wl[1] wl[2] wl[3] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar0Array_4X2
Xinst0x1 vss vdd wl[0] wl[1] wl[2] wl[3] bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar0Array_4X2
.ends SP6TVar0Array_4X4

.subckt SP6TVar0Array_8X4 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar0Array_4X4
Xinst1x0 vss vdd wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar0Array_4X4
.ends SP6TVar0Array_8X4

.subckt SP6TVar0Array_8X8 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar0Array_8X4
Xinst0x1 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7] SP6TVar0Array_8X4
.ends SP6TVar0Array_8X8

.subckt SP6TVar0BulkConn vdd vss bl bl_n
.ends SP6TVar0BulkConn

.subckt SP6TVar0BulkConnRow_2 vss vdd bl[0] bl_n[0] bl[1] bl_n[1]
Xinst0 vdd vss bl[0] bl_n[0] SP6TVar0BulkConn
Xinst1 vdd vss bl[1] bl_n[1] SP6TVar0BulkConn
.ends SP6TVar0BulkConnRow_2

.subckt SP6TVar0BulkConnRow_4 vss vdd bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3]
Xinst0 vss vdd bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar0BulkConnRow_2
Xinst1 vss vdd bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar0BulkConnRow_2
.ends SP6TVar0BulkConnRow_4

.subckt SP6TVar0BulkConnRow_8 vss vdd bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7]
Xinst0 vss vdd bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar0BulkConnRow_4
Xinst1 vss vdd bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7] SP6TVar0BulkConnRow_4
.ends SP6TVar0BulkConnRow_8

.subckt SP6TVar0Array_16X8BC vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7] SP6TVar0Array_8X8
Xinst1x0 vss vdd wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7] SP6TVar0Array_8X8
Xbottombcrow vss vdd bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7] SP6TVar0BulkConnRow_8
Xtopbcrow vss vdd bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7] SP6TVar0BulkConnRow_8
.ends SP6TVar0Array_16X8BC

.subckt zero_x1 vdd vss zero
Xnpass vss one zero vss sg13_lv_nmos l=1.3e-07 w=1.51e-06
Xppass one zero vdd vdd sg13_lv_pmos l=1.3e-07 w=1.5e-06
.ends zero_x1

.subckt SP6TVar0TestArray_16X8 vss vdd bl bl_n wl
Xarray vss vdd zero zero zero zero zero zero zero zero wl zero zero zero zero zero zero zero bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl bl_n bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7] SP6TVar0Array_16X8BC
Xzero vdd vss zero zero_x1
.ends SP6TVar0TestArray_16X8

.subckt SP6TVar0Array_4X1 vss vdd wl[0] wl[1] wl[2] wl[3] bl[0] bl_n[0]
Xinst0x0 vss vdd wl[0] wl[1] bl[0] bl_n[0] SP6TVar0Array_2X1
Xinst1x0 vss vdd wl[2] wl[3] bl[0] bl_n[0] SP6TVar0Array_2X1
.ends SP6TVar0Array_4X1

.subckt SP6TVar0Array_8X1 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] bl[0] bl_n[0] SP6TVar0Array_4X1
Xinst1x0 vss vdd wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] SP6TVar0Array_4X1
.ends SP6TVar0Array_8X1

.subckt SP6TVar0Array_16X1BC vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] bl[0] bl_n[0]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] SP6TVar0Array_8X1
Xinst1x0 vss vdd wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] bl[0] bl_n[0] SP6TVar0Array_8X1
Xbottombcrow vdd vss bl[0] bl_n[0] SP6TVar0BulkConn
Xtopbcrow vdd vss bl[0] bl_n[0] SP6TVar0BulkConn
.ends SP6TVar0Array_16X1BC

.subckt SP6TVar0Array_8X2 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar0Array_4X2
Xinst1x0 vss vdd wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar0Array_4X2
.ends SP6TVar0Array_8X2

.subckt SP6TVar0Array_16X2BC vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] bl[0] bl_n[0] bl[1] bl_n[1]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar0Array_8X2
Xinst1x0 vss vdd wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar0Array_8X2
Xbottombcrow vss vdd bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar0BulkConnRow_2
Xtopbcrow vss vdd bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar0BulkConnRow_2
.ends SP6TVar0Array_16X2BC

.subckt SP6TVar0Array_16X4BC vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar0Array_8X4
Xinst1x0 vss vdd wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar0Array_8X4
Xbottombcrow vss vdd bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar0BulkConnRow_4
Xtopbcrow vss vdd bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar0BulkConnRow_4
.ends SP6TVar0Array_16X4BC

.subckt SP6TVar0Array_6X1 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] bl[0] bl_n[0]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] bl[0] bl_n[0] SP6TVar0Array_4X1
Xinst1x0 vss vdd wl[4] wl[5] bl[0] bl_n[0] SP6TVar0Array_2X1
.ends SP6TVar0Array_6X1

.subckt SP6TVar0CellConnectOut wl bl bl_n vdd vss bit bit_n
Xpu1 vdd bit_n bit vdd sg13_lv_pmos l=1.3e-07 w=3e-07
Xpd1 bit bit_n vss vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpu2 vdd bit bit_n vdd sg13_lv_pmos l=1.3e-07 w=3e-07
Xpd2 bit_n bit vss vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg1 bit wl bl vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg2 bit_n wl bl_n vss sg13_lv_nmos l=1.3e-07 w=3e-07
.ends SP6TVar0CellConnectOut

.subckt SP6TVar0TestArray_16X8C vss vdd bl bl_n bit bit_n wl
Xarray_0 vss vdd zero zero zero zero zero zero zero zero wl zero zero zero zero zero zero zero array_0_bl[0] array_0_bl_n[0] SP6TVar0Array_16X1BC
Xarray_1 vss vdd zero zero zero zero zero zero zero zero wl zero zero zero zero zero zero zero array_1_bl[0] array_1_bl_n[0] array_1_bl[1] array_1_bl_n[1] SP6TVar0Array_16X2BC
Xarray_2 vss vdd zero zero zero zero zero zero zero zero wl zero zero zero zero zero zero zero array_2_bl[0] array_2_bl_n[0] array_2_bl[1] array_2_bl_n[1] array_2_bl[2] array_2_bl_n[2] array_2_bl[3] array_2_bl_n[3] SP6TVar0Array_16X4BC
Xcolbc_0 vdd vss bl bl_n SP6TVar0BulkConn
Xcolbc_1 vdd vss bl bl_n SP6TVar0BulkConn
Xcolarray_0 vss vdd zero zero zero zero zero zero zero zero bl bl_n SP6TVar0Array_8X1
Xcolarray_1 vss vdd zero zero zero zero zero zero bl bl_n SP6TVar0Array_6X1
Xbc_noconn zero bl bl_n vdd vss SP6TVar0Cell
Xbc_conn wl bl bl_n vdd vss bit bit_n SP6TVar0CellConnectOut
Xzero vdd vss zero zero_x1
.ends SP6TVar0TestArray_16X8C

.subckt PadFrame_SP00 PAD0x0 PAD0x1 PAD0x2 PAD0x3 PAD0x4 PAD0x5 PAD0x6 PAD0x7 PAD0x8 PAD0x9 PAD1x0 PAD1x1 PAD1x2 PAD1x3 PAD1x4 PAD1x5 PAD1x6 PAD1x7 PAD1x8 PAD1x9
XPAD0x0 PAD0x0 BondPad
XPAD0x1 PAD0x1 BondPad
XPAD0x2 PAD0x2 BondPad
XPAD0x3 PAD0x3 BondPad
XPAD0x4 PAD0x4 BondPad
XPAD0x5 PAD0x5 BondPad
XPAD0x6 PAD0x6 BondPad
XPAD0x7 PAD0x7 BondPad
XPAD0x8 PAD0x8 BondPad
XPAD0x9 PAD0x9 BondPad
XPAD1x0 PAD1x0 BondPad
XPAD1x1 PAD1x1 BondPad
XPAD1x2 PAD1x2 BondPad
XPAD1x3 PAD1x3 BondPad
XPAD1x4 PAD1x4 BondPad
XPAD1x5 PAD1x5 BondPad
XPAD1x6 PAD1x6 BondPad
XPAD1x7 PAD1x7 BondPad
XPAD1x8 PAD1x8 BondPad
XPAD1x9 PAD1x9 BondPad
.ends PadFrame_SP00

.subckt SP6TVar0 vss noco_vdd noco_wl noco_bl noco_bl_n co_vdd co_bl co_bl_n co_bit co_bit_n co_wl
Xframe noco_vdd noco_wl NoConn_PAD0x2 co_vdd co_bl_n co_bit co_bit_n NoConn_PAD0x7 NoConn_PAD0x8 NoConn_PAD0x9 vss noco_bl noco_bl_n vss co_bl co_wl NoConn_PAD1x6 NoConn_PAD1x7 NoConn_PAD1x8 NoConn_PAD1x9 PadFrame_SP00
Xtestarray_noco vss noco_vdd noco_bl noco_bl_n noco_wl SP6TVar0TestArray_16X8
Xtestarray_co vss co_vdd co_bl co_bl_n co_bit co_bit_n co_wl SP6TVar0TestArray_16X8C
.ends SP6TVar0

.subckt DP8TVar0Cell wl1 wl2 bl1 bl1_n bl2 bl2_n vdd vss
Xpu1 vdd bit_n bit vdd sg13_lv_pmos l=1.3e-07 w=3e-07
Xpd1 bit bit_n vss vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpu2 vdd bit bit_n vdd sg13_lv_pmos l=1.3e-07 w=3e-07
Xpd2 bit_n bit vss vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg1 bit wl1 bl1 vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg1n bit_n wl1 bl1_n vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg2 bit wl2 bl2 vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg2n bit_n wl2 bl2_n vss sg13_lv_nmos l=1.3e-07 w=3e-07
.ends DP8TVar0Cell

.subckt DP8TVar0Array_2X1 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0]
Xinst0x0 wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] vdd vss DP8TVar0Cell
Xinst1x0 wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0] vdd vss DP8TVar0Cell
.ends DP8TVar0Array_2X1

.subckt DP8TVar0Array_2X2 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0] DP8TVar0Array_2X1
Xinst0x1 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TVar0Array_2X1
.ends DP8TVar0Array_2X2

.subckt DP8TVar0Array_4X2 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TVar0Array_2X2
Xinst1x0 vss vdd wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TVar0Array_2X2
.ends DP8TVar0Array_4X2

.subckt DP8TVar0Array_4X4 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TVar0Array_4X2
Xinst0x1 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar0Array_4X2
.ends DP8TVar0Array_4X4

.subckt DP8TVar0Array_8X4 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar0Array_4X4
Xinst1x0 vss vdd wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar0Array_4X4
.ends DP8TVar0Array_8X4

.subckt DP8TVar0Array_8X8 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar0Array_8X4
Xinst0x1 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar0Array_8X4
.ends DP8TVar0Array_8X8

.subckt DP8TVar0BulkConn vdd vss bl1 bl2 bl1_n bl2_n
.ends DP8TVar0BulkConn

.subckt DP8TVar0BulkConnRow_2 vss vdd bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1]
Xinst0 vdd vss bl1[0] bl2[0] bl1_n[0] bl2_n[0] DP8TVar0BulkConn
Xinst1 vdd vss bl1[1] bl2[1] bl1_n[1] bl2_n[1] DP8TVar0BulkConn
.ends DP8TVar0BulkConnRow_2

.subckt DP8TVar0BulkConnRow_4 vss vdd bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3]
Xinst0 vss vdd bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TVar0BulkConnRow_2
Xinst1 vss vdd bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar0BulkConnRow_2
.ends DP8TVar0BulkConnRow_4

.subckt DP8TVar0BulkConnRow_8 vss vdd bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0 vss vdd bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar0BulkConnRow_4
Xinst1 vss vdd bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar0BulkConnRow_4
.ends DP8TVar0BulkConnRow_8

.subckt DP8TVar0Array_16X8BC vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] wl1[8] wl2[8] wl1[9] wl2[9] wl1[10] wl2[10] wl1[11] wl2[11] wl1[12] wl2[12] wl1[13] wl2[13] wl1[14] wl2[14] wl1[15] wl2[15] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar0Array_8X8
Xinst1x0 vss vdd wl1[8] wl2[8] wl1[9] wl2[9] wl1[10] wl2[10] wl1[11] wl2[11] wl1[12] wl2[12] wl1[13] wl2[13] wl1[14] wl2[14] wl1[15] wl2[15] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar0Array_8X8
Xbottombcrow vss vdd bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar0BulkConnRow_8
Xtopbcrow vss vdd bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar0BulkConnRow_8
.ends DP8TVar0Array_16X8BC

.subckt DP8TVar0TestArray_16X8 vss vdd wl1 wl2 bl1 bl1_n bl2 bl2_n
Xarray vss vdd zero zero zero zero zero zero zero zero zero zero zero zero zero zero zero zero wl1 wl2 zero zero zero zero zero zero zero zero zero zero zero zero zero zero bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1 bl1_n bl2 bl2_n bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar0Array_16X8BC
Xzero vdd vss zero zero_x1
.ends DP8TVar0TestArray_16X8

.subckt DP8TVar0Array_4X8 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar0Array_4X4
Xinst0x1 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar0Array_4X4
.ends DP8TVar0Array_4X8

.subckt DP8TVar0Array_2X4 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TVar0Array_2X2
Xinst0x1 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar0Array_2X2
.ends DP8TVar0Array_2X4

.subckt DP8TVar0Array_2X8 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar0Array_2X4
Xinst0x1 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar0Array_2X4
.ends DP8TVar0Array_2X8

.subckt DP8TVar0Array_1X2 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1]
Xinst0x0 wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] vdd vss DP8TVar0Cell
Xinst0x1 wl1[0] wl2[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] vdd vss DP8TVar0Cell
.ends DP8TVar0Array_1X2

.subckt DP8TVar0Array_1X4 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3]
Xinst0x0 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TVar0Array_1X2
Xinst0x1 vss vdd wl1[0] wl2[0] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar0Array_1X2
.ends DP8TVar0Array_1X4

.subckt DP8TVar0Array_1X8 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar0Array_1X4
Xinst0x1 vss vdd wl1[0] wl2[0] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar0Array_1X4
.ends DP8TVar0Array_1X8

.subckt DP8TVar0Array_7X8 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar0Array_4X8
Xinst1x0 vss vdd wl1[4] wl2[4] wl1[5] wl2[5] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar0Array_2X8
Xinst2x0 vss vdd wl1[6] wl2[6] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar0Array_1X8
.ends DP8TVar0Array_7X8

.subckt DP8TVar0CellShWL1 wl1 wl2 bl1 bl1_n bl2 bl2_n vdd vss
Xpu1 vdd bit_n bit vdd sg13_lv_pmos l=1.3e-07 w=3e-07
Xpd1 bit bit_n vss vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpu2 vdd bit bit_n vdd sg13_lv_pmos l=1.3e-07 w=3e-07
Xpd2 bit_n bit vss vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg1 bit wl1 bl1 vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg1n bit_n wl1 bl1_n vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg2 bit wl1 bl2 vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg2n bit_n wl1 bl2_n vss sg13_lv_nmos l=1.3e-07 w=3e-07
.ends DP8TVar0CellShWL1

.subckt DP8TVar0ArrayShWL1_1X2 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1]
Xinst0x0 wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] vdd vss DP8TVar0CellShWL1
Xinst0x1 wl1[0] wl2[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] vdd vss DP8TVar0CellShWL1
.ends DP8TVar0ArrayShWL1_1X2

.subckt DP8TVar0ArrayShWL1_1X4 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3]
Xinst0x0 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TVar0ArrayShWL1_1X2
Xinst0x1 vss vdd wl1[0] wl2[0] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar0ArrayShWL1_1X2
.ends DP8TVar0ArrayShWL1_1X4

.subckt DP8TVar0ArrayShWL1_1X8 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar0ArrayShWL1_1X4
Xinst0x1 vss vdd wl1[0] wl2[0] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar0ArrayShWL1_1X4
.ends DP8TVar0ArrayShWL1_1X8

.subckt DP8TVar0CellConnectOut wl1 wl2 bl1 bl1_n bl2 bl2_n vdd vss bit bit_n
Xpu1 vdd bit_n bit vdd sg13_lv_pmos l=1.3e-07 w=3e-07
Xpd1 bit bit_n vss vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpu2 vdd bit bit_n vdd sg13_lv_pmos l=1.3e-07 w=3e-07
Xpd2 bit_n bit vss vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg1 bit wl1 bl1 vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg1n bit_n wl1 bl1_n vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg2 bit wl2 bl2 vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg2n bit_n wl2 bl2_n vss sg13_lv_nmos l=1.3e-07 w=3e-07
.ends DP8TVar0CellConnectOut

.subckt DP8TVar0CellShWL2 wl1 wl2 bl1 bl1_n bl2 bl2_n vdd vss
Xpu1 vdd bit_n bit vdd sg13_lv_pmos l=1.3e-07 w=3e-07
Xpd1 bit bit_n vss vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpu2 vdd bit bit_n vdd sg13_lv_pmos l=1.3e-07 w=3e-07
Xpd2 bit_n bit vss vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg1 bit wl2 bl1 vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg1n bit_n wl2 bl1_n vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg2 bit wl2 bl2 vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg2n bit_n wl2 bl2_n vss sg13_lv_nmos l=1.3e-07 w=3e-07
.ends DP8TVar0CellShWL2

.subckt DP8TVar0ArrayShWL2_1X2 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1]
Xinst0x0 wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] vdd vss DP8TVar0CellShWL2
Xinst0x1 wl1[0] wl2[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] vdd vss DP8TVar0CellShWL2
.ends DP8TVar0ArrayShWL2_1X2

.subckt DP8TVar0ArrayShWL2_1X4 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3]
Xinst0x0 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TVar0ArrayShWL2_1X2
Xinst0x1 vss vdd wl1[0] wl2[0] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar0ArrayShWL2_1X2
.ends DP8TVar0ArrayShWL2_1X4

.subckt DP8TVar0ArrayShWL2_1X8 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar0ArrayShWL2_1X4
Xinst0x1 vss vdd wl1[0] wl2[0] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar0ArrayShWL2_1X4
.ends DP8TVar0ArrayShWL2_1X8

.subckt DP8TVar0Array_6X8 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar0Array_4X8
Xinst1x0 vss vdd wl1[4] wl2[4] wl1[5] wl2[5] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar0Array_2X8
.ends DP8TVar0Array_6X8

.subckt DP8TVar0TestArray_16X8C vss vdd wl1 wl2 bl1 bl1_n bl2 bl2_n bit bit_n
Xbcconn_bot vss vdd bcconn_bot_bl1[0] bcconn_bot_bl1_n[0] bcconn_bot_bl2[0] bcconn_bot_bl2_n[0] bcconn_bot_bl1[1] bcconn_bot_bl1_n[1] bcconn_bot_bl2[1] bcconn_bot_bl2_n[1] bcconn_bot_bl1[2] bcconn_bot_bl1_n[2] bcconn_bot_bl2[2] bcconn_bot_bl2_n[2] bcconn_bot_bl1[3] bcconn_bot_bl1_n[3] bcconn_bot_bl2[3] bcconn_bot_bl2_n[3] bl1 bl1_n bl2 bl2_n bcconn_bot_bl1[5] bcconn_bot_bl1_n[5] bcconn_bot_bl2[5] bcconn_bot_bl2_n[5] bcconn_bot_bl1[6] bcconn_bot_bl1_n[6] bcconn_bot_bl2[6] bcconn_bot_bl2_n[6] bcconn_bot_bl1[7] bcconn_bot_bl1_n[7] bcconn_bot_bl2[7] bcconn_bot_bl2_n[7] DP8TVar0BulkConnRow_8
Xbcconn_top vss vdd bcconn_top_bl1[0] bcconn_top_bl1_n[0] bcconn_top_bl2[0] bcconn_top_bl2_n[0] bcconn_top_bl1[1] bcconn_top_bl1_n[1] bcconn_top_bl2[1] bcconn_top_bl2_n[1] bcconn_top_bl1[2] bcconn_top_bl1_n[2] bcconn_top_bl2[2] bcconn_top_bl2_n[2] bcconn_top_bl1[3] bcconn_top_bl1_n[3] bcconn_top_bl2[3] bcconn_top_bl2_n[3] bl1 bl1_n bl2 bl2_n bcconn_top_bl1[5] bcconn_top_bl1_n[5] bcconn_top_bl2[5] bcconn_top_bl2_n[5] bcconn_top_bl1[6] bcconn_top_bl1_n[6] bcconn_top_bl2[6] bcconn_top_bl2_n[6] bcconn_top_bl1[7] bcconn_top_bl1_n[7] bcconn_top_bl2[7] bcconn_top_bl2_n[7] DP8TVar0BulkConnRow_8
Xarray_bot vss vdd zero zero zero zero zero zero zero zero zero zero zero zero zero zero array_bot_bl1[0] array_bot_bl1_n[0] array_bot_bl2[0] array_bot_bl2_n[0] array_bot_bl1[1] array_bot_bl1_n[1] array_bot_bl2[1] array_bot_bl2_n[1] array_bot_bl1[2] array_bot_bl1_n[2] array_bot_bl2[2] array_bot_bl2_n[2] array_bot_bl1[3] array_bot_bl1_n[3] array_bot_bl2[3] array_bot_bl2_n[3] bl1 bl1_n bl2 bl2_n array_bot_bl1[5] array_bot_bl1_n[5] array_bot_bl2[5] array_bot_bl2_n[5] array_bot_bl1[6] array_bot_bl1_n[6] array_bot_bl2[6] array_bot_bl2_n[6] array_bot_bl1[7] array_bot_bl1_n[7] array_bot_bl2[7] array_bot_bl2_n[7] DP8TVar0Array_7X8
Xshwl1_row vss vdd zero bit shwl1_row_bl1[0] shwl1_row_bl1_n[0] shwl1_row_bl2[0] shwl1_row_bl2_n[0] shwl1_row_bl1[1] shwl1_row_bl1_n[1] shwl1_row_bl2[1] shwl1_row_bl2_n[1] shwl1_row_bl1[2] shwl1_row_bl1_n[2] shwl1_row_bl2[2] shwl1_row_bl2_n[2] shwl1_row_bl1[3] shwl1_row_bl1_n[3] shwl1_row_bl2[3] shwl1_row_bl2_n[3] bl1 bl1_n bl2 bl2_n shwl1_row_bl1[5] shwl1_row_bl1_n[5] shwl1_row_bl2[5] shwl1_row_bl2_n[5] shwl1_row_bl1[6] shwl1_row_bl1_n[6] shwl1_row_bl2[6] shwl1_row_bl2_n[6] shwl1_row_bl1[7] shwl1_row_bl1_n[7] shwl1_row_bl2[7] shwl1_row_bl2_n[7] DP8TVar0ArrayShWL1_1X8
Xcell_cols_left vss vdd wl1 wl2 cell_cols_left_bl1[0] cell_cols_left_bl1_n[0] cell_cols_left_bl2[0] cell_cols_left_bl2_n[0] cell_cols_left_bl1[1] cell_cols_left_bl1_n[1] cell_cols_left_bl2[1] cell_cols_left_bl2_n[1] cell_cols_left_bl1[2] cell_cols_left_bl1_n[2] cell_cols_left_bl2[2] cell_cols_left_bl2_n[2] cell_cols_left_bl1[3] cell_cols_left_bl1_n[3] cell_cols_left_bl2[3] cell_cols_left_bl2_n[3] DP8TVar0Array_1X4
Xconncell wl1 wl2 bl1 bl1_n bl2 bl2_n vdd vss bit bit_n DP8TVar0CellConnectOut
Xfillcell wl1 wl2 fillcell_bl1 fillcell_bl1_n fillcell_bl2 fillcell_bl2_n vdd vss DP8TVar0Cell
Xcell_cols_right vss vdd wl1 wl2 cell_cols_right_bl1[0] cell_cols_right_bl1_n[0] cell_cols_right_bl2[0] cell_cols_right_bl2_n[0] cell_cols_right_bl1[1] cell_cols_right_bl1_n[1] cell_cols_right_bl2[1] cell_cols_right_bl2_n[1] DP8TVar0Array_1X2
Xshwl2_row vss vdd bit_n zero shwl2_row_bl1[0] shwl2_row_bl1_n[0] shwl2_row_bl2[0] shwl2_row_bl2_n[0] shwl2_row_bl1[1] shwl2_row_bl1_n[1] shwl2_row_bl2[1] shwl2_row_bl2_n[1] shwl2_row_bl1[2] shwl2_row_bl1_n[2] shwl2_row_bl2[2] shwl2_row_bl2_n[2] shwl2_row_bl1[3] shwl2_row_bl1_n[3] shwl2_row_bl2[3] shwl2_row_bl2_n[3] bl1 bl1_n bl2 bl2_n shwl2_row_bl1[5] shwl2_row_bl1_n[5] shwl2_row_bl2[5] shwl2_row_bl2_n[5] shwl2_row_bl1[6] shwl2_row_bl1_n[6] shwl2_row_bl2[6] shwl2_row_bl2_n[6] shwl2_row_bl1[7] shwl2_row_bl1_n[7] shwl2_row_bl2[7] shwl2_row_bl2_n[7] DP8TVar0ArrayShWL2_1X8
Xarray_top vss vdd zero zero zero zero zero zero zero zero zero zero zero zero array_top_bl1[0] array_top_bl1_n[0] array_top_bl2[0] array_top_bl2_n[0] array_top_bl1[1] array_top_bl1_n[1] array_top_bl2[1] array_top_bl2_n[1] array_top_bl1[2] array_top_bl1_n[2] array_top_bl2[2] array_top_bl2_n[2] array_top_bl1[3] array_top_bl1_n[3] array_top_bl2[3] array_top_bl2_n[3] bl1 bl1_n bl2 bl2_n array_top_bl1[5] array_top_bl1_n[5] array_top_bl2[5] array_top_bl2_n[5] array_top_bl1[6] array_top_bl1_n[6] array_top_bl2[6] array_top_bl2_n[6] array_top_bl1[7] array_top_bl1_n[7] array_top_bl2[7] array_top_bl2_n[7] DP8TVar0Array_6X8
Xzero vdd vss zero zero_x1
.ends DP8TVar0TestArray_16X8C

.subckt PadFrame_DP00 PAD0x0 PAD0x1 PAD0x2 PAD0x3 PAD0x4 PAD0x5 PAD0x6 PAD0x7 PAD0x8 PAD0x9 PAD1x0 PAD1x1 PAD1x2 PAD1x3 PAD1x4 PAD1x5 PAD1x6 PAD1x7 PAD1x8 PAD1x9
XPAD0x0 PAD0x0 BondPad
XPAD0x1 PAD0x1 BondPad
XPAD0x2 PAD0x2 BondPad
XPAD0x3 PAD0x3 BondPad
XPAD0x4 PAD0x4 BondPad
XPAD0x5 PAD0x5 BondPad
XPAD0x6 PAD0x6 BondPad
XPAD0x7 PAD0x7 BondPad
XPAD0x8 PAD0x8 BondPad
XPAD0x9 PAD0x9 BondPad
XPAD1x0 PAD1x0 BondPad
XPAD1x1 PAD1x1 BondPad
XPAD1x2 PAD1x2 BondPad
XPAD1x3 PAD1x3 BondPad
XPAD1x4 PAD1x4 BondPad
XPAD1x5 PAD1x5 BondPad
XPAD1x6 PAD1x6 BondPad
XPAD1x7 PAD1x7 BondPad
XPAD1x8 PAD1x8 BondPad
XPAD1x9 PAD1x9 BondPad
.ends PadFrame_DP00

.subckt DP8TVar0 vss noco_vdd noco_wl1 noco_wl2 noco_bl1 noco_bl1_n noco_bl2 noco_bl2_n co_vdd co_bit co_bit_n co_wl1 co_wl2 co_bl1 co_bl1_n co_bl2_n co_bl2
Xframe noco_vdd noco_wl1 noco_wl2 noco_bl2 co_vdd co_bit co_bit_n co_wl1 co_wl2 NoConn_PAD0x9 vss noco_bl1 noco_bl1_n noco_bl2_n vss co_bl1 co_bl1_n co_bl2_n co_bl2 NoConn_PAD1x9 PadFrame_DP00
Xtestarray_noco vss noco_vdd noco_wl1 noco_wl2 noco_bl1 noco_bl1_n noco_bl2 noco_bl2_n DP8TVar0TestArray_16X8
Xtestarray_co vss co_vdd co_wl1 co_wl2 co_bl1 co_bl1_n co_bl2 co_bl2_n co_bit co_bit_n DP8TVar0TestArray_16X8C
.ends DP8TVar0

.subckt SP6TVar1Cell wl bl bl_n vdd vss
Xpu1 vdd bit_n bit vdd sg13_lv_pmos l=1.3e-07 w=2e-07
Xpd1 bit bit_n vss vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpu2 vdd bit bit_n vdd sg13_lv_pmos l=1.3e-07 w=2e-07
Xpd2 bit_n bit vss vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg1 bit wl bl vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg2 bit_n wl bl_n vss sg13_lv_nmos l=1.3e-07 w=3e-07
.ends SP6TVar1Cell

.subckt SP6TVar1Array_2X1 vss vdd wl[0] wl[1] bl[0] bl_n[0]
Xinst0x0 wl[0] bl[0] bl_n[0] vdd vss SP6TVar1Cell
Xinst1x0 wl[1] bl[0] bl_n[0] vdd vss SP6TVar1Cell
.ends SP6TVar1Array_2X1

.subckt SP6TVar1Array_2X2 vss vdd wl[0] wl[1] bl[0] bl_n[0] bl[1] bl_n[1]
Xinst0x0 vss vdd wl[0] wl[1] bl[0] bl_n[0] SP6TVar1Array_2X1
Xinst0x1 vss vdd wl[0] wl[1] bl[1] bl_n[1] SP6TVar1Array_2X1
.ends SP6TVar1Array_2X2

.subckt SP6TVar1Array_4X2 vss vdd wl[0] wl[1] wl[2] wl[3] bl[0] bl_n[0] bl[1] bl_n[1]
Xinst0x0 vss vdd wl[0] wl[1] bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar1Array_2X2
Xinst1x0 vss vdd wl[2] wl[3] bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar1Array_2X2
.ends SP6TVar1Array_4X2

.subckt SP6TVar1Array_4X4 vss vdd wl[0] wl[1] wl[2] wl[3] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar1Array_4X2
Xinst0x1 vss vdd wl[0] wl[1] wl[2] wl[3] bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar1Array_4X2
.ends SP6TVar1Array_4X4

.subckt SP6TVar1Array_8X4 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar1Array_4X4
Xinst1x0 vss vdd wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar1Array_4X4
.ends SP6TVar1Array_8X4

.subckt SP6TVar1Array_8X8 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar1Array_8X4
Xinst0x1 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7] SP6TVar1Array_8X4
.ends SP6TVar1Array_8X8

.subckt SP6TVar1BulkConn vdd vss bl bl_n
.ends SP6TVar1BulkConn

.subckt SP6TVar1BulkConnRow_2 vss vdd bl[0] bl_n[0] bl[1] bl_n[1]
Xinst0 vdd vss bl[0] bl_n[0] SP6TVar1BulkConn
Xinst1 vdd vss bl[1] bl_n[1] SP6TVar1BulkConn
.ends SP6TVar1BulkConnRow_2

.subckt SP6TVar1BulkConnRow_4 vss vdd bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3]
Xinst0 vss vdd bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar1BulkConnRow_2
Xinst1 vss vdd bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar1BulkConnRow_2
.ends SP6TVar1BulkConnRow_4

.subckt SP6TVar1BulkConnRow_8 vss vdd bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7]
Xinst0 vss vdd bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar1BulkConnRow_4
Xinst1 vss vdd bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7] SP6TVar1BulkConnRow_4
.ends SP6TVar1BulkConnRow_8

.subckt SP6TVar1Array_16X8BC vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7] SP6TVar1Array_8X8
Xinst1x0 vss vdd wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7] SP6TVar1Array_8X8
Xbottombcrow vss vdd bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7] SP6TVar1BulkConnRow_8
Xtopbcrow vss vdd bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7] SP6TVar1BulkConnRow_8
.ends SP6TVar1Array_16X8BC

.subckt SP6TVar1TestArray_16X8 vss vdd bl bl_n wl
Xarray vss vdd zero zero zero zero zero zero zero zero wl zero zero zero zero zero zero zero bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl bl_n bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7] SP6TVar1Array_16X8BC
Xzero vdd vss zero zero_x1
.ends SP6TVar1TestArray_16X8

.subckt SP6TVar1Array_4X1 vss vdd wl[0] wl[1] wl[2] wl[3] bl[0] bl_n[0]
Xinst0x0 vss vdd wl[0] wl[1] bl[0] bl_n[0] SP6TVar1Array_2X1
Xinst1x0 vss vdd wl[2] wl[3] bl[0] bl_n[0] SP6TVar1Array_2X1
.ends SP6TVar1Array_4X1

.subckt SP6TVar1Array_8X1 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] bl[0] bl_n[0] SP6TVar1Array_4X1
Xinst1x0 vss vdd wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] SP6TVar1Array_4X1
.ends SP6TVar1Array_8X1

.subckt SP6TVar1Array_16X1BC vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] bl[0] bl_n[0]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] SP6TVar1Array_8X1
Xinst1x0 vss vdd wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] bl[0] bl_n[0] SP6TVar1Array_8X1
Xbottombcrow vdd vss bl[0] bl_n[0] SP6TVar1BulkConn
Xtopbcrow vdd vss bl[0] bl_n[0] SP6TVar1BulkConn
.ends SP6TVar1Array_16X1BC

.subckt SP6TVar1Array_8X2 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar1Array_4X2
Xinst1x0 vss vdd wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar1Array_4X2
.ends SP6TVar1Array_8X2

.subckt SP6TVar1Array_16X2BC vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] bl[0] bl_n[0] bl[1] bl_n[1]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar1Array_8X2
Xinst1x0 vss vdd wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar1Array_8X2
Xbottombcrow vss vdd bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar1BulkConnRow_2
Xtopbcrow vss vdd bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar1BulkConnRow_2
.ends SP6TVar1Array_16X2BC

.subckt SP6TVar1Array_16X4BC vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar1Array_8X4
Xinst1x0 vss vdd wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar1Array_8X4
Xbottombcrow vss vdd bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar1BulkConnRow_4
Xtopbcrow vss vdd bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar1BulkConnRow_4
.ends SP6TVar1Array_16X4BC

.subckt SP6TVar1Array_6X1 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] bl[0] bl_n[0]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] bl[0] bl_n[0] SP6TVar1Array_4X1
Xinst1x0 vss vdd wl[4] wl[5] bl[0] bl_n[0] SP6TVar1Array_2X1
.ends SP6TVar1Array_6X1

.subckt SP6TVar1CellConnectOut wl bl bl_n vdd vss bit bit_n
Xpu1 vdd bit_n bit vdd sg13_lv_pmos l=1.3e-07 w=2e-07
Xpd1 bit bit_n vss vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpu2 vdd bit bit_n vdd sg13_lv_pmos l=1.3e-07 w=2e-07
Xpd2 bit_n bit vss vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg1 bit wl bl vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg2 bit_n wl bl_n vss sg13_lv_nmos l=1.3e-07 w=3e-07
.ends SP6TVar1CellConnectOut

.subckt SP6TVar1TestArray_16X8C vss vdd bl bl_n bit bit_n wl
Xarray_0 vss vdd zero zero zero zero zero zero zero zero wl zero zero zero zero zero zero zero array_0_bl[0] array_0_bl_n[0] SP6TVar1Array_16X1BC
Xarray_1 vss vdd zero zero zero zero zero zero zero zero wl zero zero zero zero zero zero zero array_1_bl[0] array_1_bl_n[0] array_1_bl[1] array_1_bl_n[1] SP6TVar1Array_16X2BC
Xarray_2 vss vdd zero zero zero zero zero zero zero zero wl zero zero zero zero zero zero zero array_2_bl[0] array_2_bl_n[0] array_2_bl[1] array_2_bl_n[1] array_2_bl[2] array_2_bl_n[2] array_2_bl[3] array_2_bl_n[3] SP6TVar1Array_16X4BC
Xcolbc_0 vdd vss bl bl_n SP6TVar1BulkConn
Xcolbc_1 vdd vss bl bl_n SP6TVar1BulkConn
Xcolarray_0 vss vdd zero zero zero zero zero zero zero zero bl bl_n SP6TVar1Array_8X1
Xcolarray_1 vss vdd zero zero zero zero zero zero bl bl_n SP6TVar1Array_6X1
Xbc_noconn zero bl bl_n vdd vss SP6TVar1Cell
Xbc_conn wl bl bl_n vdd vss bit bit_n SP6TVar1CellConnectOut
Xzero vdd vss zero zero_x1
.ends SP6TVar1TestArray_16X8C

.subckt PadFrame_SP01 PAD0x0 PAD0x1 PAD0x2 PAD0x3 PAD0x4 PAD0x5 PAD0x6 PAD0x7 PAD0x8 PAD0x9 PAD1x0 PAD1x1 PAD1x2 PAD1x3 PAD1x4 PAD1x5 PAD1x6 PAD1x7 PAD1x8 PAD1x9
XPAD0x0 PAD0x0 BondPad
XPAD0x1 PAD0x1 BondPad
XPAD0x2 PAD0x2 BondPad
XPAD0x3 PAD0x3 BondPad
XPAD0x4 PAD0x4 BondPad
XPAD0x5 PAD0x5 BondPad
XPAD0x6 PAD0x6 BondPad
XPAD0x7 PAD0x7 BondPad
XPAD0x8 PAD0x8 BondPad
XPAD0x9 PAD0x9 BondPad
XPAD1x0 PAD1x0 BondPad
XPAD1x1 PAD1x1 BondPad
XPAD1x2 PAD1x2 BondPad
XPAD1x3 PAD1x3 BondPad
XPAD1x4 PAD1x4 BondPad
XPAD1x5 PAD1x5 BondPad
XPAD1x6 PAD1x6 BondPad
XPAD1x7 PAD1x7 BondPad
XPAD1x8 PAD1x8 BondPad
XPAD1x9 PAD1x9 BondPad
.ends PadFrame_SP01

.subckt SP6TVar1 vss noco_vdd noco_wl noco_bl noco_bl_n co_vdd co_bl co_bl_n co_bit co_bit_n co_wl
Xframe noco_vdd noco_wl NoConn_PAD0x2 co_vdd co_bl_n co_bit co_bit_n NoConn_PAD0x7 NoConn_PAD0x8 NoConn_PAD0x9 vss noco_bl noco_bl_n vss co_bl co_wl NoConn_PAD1x6 NoConn_PAD1x7 NoConn_PAD1x8 NoConn_PAD1x9 PadFrame_SP01
Xtestarray_noco vss noco_vdd noco_bl noco_bl_n noco_wl SP6TVar1TestArray_16X8
Xtestarray_co vss co_vdd co_bl co_bl_n co_bit co_bit_n co_wl SP6TVar1TestArray_16X8C
.ends SP6TVar1

.subckt DP8TVar1Cell wl1 wl2 bl1 bl1_n bl2 bl2_n vdd vss
Xpu1 vdd bit_n bit vdd sg13_lv_pmos l=1.3e-07 w=2e-07
Xpd1 bit bit_n vss vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpu2 vdd bit bit_n vdd sg13_lv_pmos l=1.3e-07 w=2e-07
Xpd2 bit_n bit vss vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg1 bit wl1 bl1 vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg1n bit_n wl1 bl1_n vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg2 bit wl2 bl2 vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg2n bit_n wl2 bl2_n vss sg13_lv_nmos l=1.3e-07 w=3e-07
.ends DP8TVar1Cell

.subckt DP8TVar1Array_2X1 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0]
Xinst0x0 wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] vdd vss DP8TVar1Cell
Xinst1x0 wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0] vdd vss DP8TVar1Cell
.ends DP8TVar1Array_2X1

.subckt DP8TVar1Array_2X2 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0] DP8TVar1Array_2X1
Xinst0x1 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TVar1Array_2X1
.ends DP8TVar1Array_2X2

.subckt DP8TVar1Array_4X2 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TVar1Array_2X2
Xinst1x0 vss vdd wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TVar1Array_2X2
.ends DP8TVar1Array_4X2

.subckt DP8TVar1Array_4X4 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TVar1Array_4X2
Xinst0x1 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar1Array_4X2
.ends DP8TVar1Array_4X4

.subckt DP8TVar1Array_8X4 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar1Array_4X4
Xinst1x0 vss vdd wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar1Array_4X4
.ends DP8TVar1Array_8X4

.subckt DP8TVar1Array_8X8 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar1Array_8X4
Xinst0x1 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar1Array_8X4
.ends DP8TVar1Array_8X8

.subckt DP8TVar1BulkConn vdd vss bl1 bl2 bl1_n bl2_n
.ends DP8TVar1BulkConn

.subckt DP8TVar1BulkConnRow_2 vss vdd bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1]
Xinst0 vdd vss bl1[0] bl2[0] bl1_n[0] bl2_n[0] DP8TVar1BulkConn
Xinst1 vdd vss bl1[1] bl2[1] bl1_n[1] bl2_n[1] DP8TVar1BulkConn
.ends DP8TVar1BulkConnRow_2

.subckt DP8TVar1BulkConnRow_4 vss vdd bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3]
Xinst0 vss vdd bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TVar1BulkConnRow_2
Xinst1 vss vdd bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar1BulkConnRow_2
.ends DP8TVar1BulkConnRow_4

.subckt DP8TVar1BulkConnRow_8 vss vdd bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0 vss vdd bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar1BulkConnRow_4
Xinst1 vss vdd bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar1BulkConnRow_4
.ends DP8TVar1BulkConnRow_8

.subckt DP8TVar1Array_16X8BC vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] wl1[8] wl2[8] wl1[9] wl2[9] wl1[10] wl2[10] wl1[11] wl2[11] wl1[12] wl2[12] wl1[13] wl2[13] wl1[14] wl2[14] wl1[15] wl2[15] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar1Array_8X8
Xinst1x0 vss vdd wl1[8] wl2[8] wl1[9] wl2[9] wl1[10] wl2[10] wl1[11] wl2[11] wl1[12] wl2[12] wl1[13] wl2[13] wl1[14] wl2[14] wl1[15] wl2[15] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar1Array_8X8
Xbottombcrow vss vdd bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar1BulkConnRow_8
Xtopbcrow vss vdd bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar1BulkConnRow_8
.ends DP8TVar1Array_16X8BC

.subckt DP8TVar1TestArray_16X8 vss vdd wl1 wl2 bl1 bl1_n bl2 bl2_n
Xarray vss vdd zero zero zero zero zero zero zero zero zero zero zero zero zero zero zero zero wl1 wl2 zero zero zero zero zero zero zero zero zero zero zero zero zero zero bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1 bl1_n bl2 bl2_n bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar1Array_16X8BC
Xzero vdd vss zero zero_x1
.ends DP8TVar1TestArray_16X8

.subckt DP8TVar1Array_4X8 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar1Array_4X4
Xinst0x1 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar1Array_4X4
.ends DP8TVar1Array_4X8

.subckt DP8TVar1Array_2X4 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TVar1Array_2X2
Xinst0x1 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar1Array_2X2
.ends DP8TVar1Array_2X4

.subckt DP8TVar1Array_2X8 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar1Array_2X4
Xinst0x1 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar1Array_2X4
.ends DP8TVar1Array_2X8

.subckt DP8TVar1Array_1X2 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1]
Xinst0x0 wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] vdd vss DP8TVar1Cell
Xinst0x1 wl1[0] wl2[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] vdd vss DP8TVar1Cell
.ends DP8TVar1Array_1X2

.subckt DP8TVar1Array_1X4 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3]
Xinst0x0 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TVar1Array_1X2
Xinst0x1 vss vdd wl1[0] wl2[0] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar1Array_1X2
.ends DP8TVar1Array_1X4

.subckt DP8TVar1Array_1X8 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar1Array_1X4
Xinst0x1 vss vdd wl1[0] wl2[0] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar1Array_1X4
.ends DP8TVar1Array_1X8

.subckt DP8TVar1Array_7X8 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar1Array_4X8
Xinst1x0 vss vdd wl1[4] wl2[4] wl1[5] wl2[5] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar1Array_2X8
Xinst2x0 vss vdd wl1[6] wl2[6] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar1Array_1X8
.ends DP8TVar1Array_7X8

.subckt DP8TVar1CellShWL1 wl1 wl2 bl1 bl1_n bl2 bl2_n vdd vss
Xpu1 vdd bit_n bit vdd sg13_lv_pmos l=1.3e-07 w=2e-07
Xpd1 bit bit_n vss vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpu2 vdd bit bit_n vdd sg13_lv_pmos l=1.3e-07 w=2e-07
Xpd2 bit_n bit vss vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg1 bit wl1 bl1 vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg1n bit_n wl1 bl1_n vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg2 bit wl1 bl2 vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg2n bit_n wl1 bl2_n vss sg13_lv_nmos l=1.3e-07 w=3e-07
.ends DP8TVar1CellShWL1

.subckt DP8TVar1ArrayShWL1_1X2 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1]
Xinst0x0 wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] vdd vss DP8TVar1CellShWL1
Xinst0x1 wl1[0] wl2[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] vdd vss DP8TVar1CellShWL1
.ends DP8TVar1ArrayShWL1_1X2

.subckt DP8TVar1ArrayShWL1_1X4 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3]
Xinst0x0 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TVar1ArrayShWL1_1X2
Xinst0x1 vss vdd wl1[0] wl2[0] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar1ArrayShWL1_1X2
.ends DP8TVar1ArrayShWL1_1X4

.subckt DP8TVar1ArrayShWL1_1X8 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar1ArrayShWL1_1X4
Xinst0x1 vss vdd wl1[0] wl2[0] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar1ArrayShWL1_1X4
.ends DP8TVar1ArrayShWL1_1X8

.subckt DP8TVar1CellConnectOut wl1 wl2 bl1 bl1_n bl2 bl2_n vdd vss bit bit_n
Xpu1 vdd bit_n bit vdd sg13_lv_pmos l=1.3e-07 w=2e-07
Xpd1 bit bit_n vss vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpu2 vdd bit bit_n vdd sg13_lv_pmos l=1.3e-07 w=2e-07
Xpd2 bit_n bit vss vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg1 bit wl1 bl1 vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg1n bit_n wl1 bl1_n vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg2 bit wl2 bl2 vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg2n bit_n wl2 bl2_n vss sg13_lv_nmos l=1.3e-07 w=3e-07
.ends DP8TVar1CellConnectOut

.subckt DP8TVar1CellShWL2 wl1 wl2 bl1 bl1_n bl2 bl2_n vdd vss
Xpu1 vdd bit_n bit vdd sg13_lv_pmos l=1.3e-07 w=2e-07
Xpd1 bit bit_n vss vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpu2 vdd bit bit_n vdd sg13_lv_pmos l=1.3e-07 w=2e-07
Xpd2 bit_n bit vss vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg1 bit wl2 bl1 vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg1n bit_n wl2 bl1_n vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg2 bit wl2 bl2 vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg2n bit_n wl2 bl2_n vss sg13_lv_nmos l=1.3e-07 w=3e-07
.ends DP8TVar1CellShWL2

.subckt DP8TVar1ArrayShWL2_1X2 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1]
Xinst0x0 wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] vdd vss DP8TVar1CellShWL2
Xinst0x1 wl1[0] wl2[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] vdd vss DP8TVar1CellShWL2
.ends DP8TVar1ArrayShWL2_1X2

.subckt DP8TVar1ArrayShWL2_1X4 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3]
Xinst0x0 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TVar1ArrayShWL2_1X2
Xinst0x1 vss vdd wl1[0] wl2[0] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar1ArrayShWL2_1X2
.ends DP8TVar1ArrayShWL2_1X4

.subckt DP8TVar1ArrayShWL2_1X8 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar1ArrayShWL2_1X4
Xinst0x1 vss vdd wl1[0] wl2[0] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar1ArrayShWL2_1X4
.ends DP8TVar1ArrayShWL2_1X8

.subckt DP8TVar1Array_6X8 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar1Array_4X8
Xinst1x0 vss vdd wl1[4] wl2[4] wl1[5] wl2[5] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar1Array_2X8
.ends DP8TVar1Array_6X8

.subckt DP8TVar1TestArray_16X8C vss vdd wl1 wl2 bl1 bl1_n bl2 bl2_n bit bit_n
Xbcconn_bot vss vdd bcconn_bot_bl1[0] bcconn_bot_bl1_n[0] bcconn_bot_bl2[0] bcconn_bot_bl2_n[0] bcconn_bot_bl1[1] bcconn_bot_bl1_n[1] bcconn_bot_bl2[1] bcconn_bot_bl2_n[1] bcconn_bot_bl1[2] bcconn_bot_bl1_n[2] bcconn_bot_bl2[2] bcconn_bot_bl2_n[2] bcconn_bot_bl1[3] bcconn_bot_bl1_n[3] bcconn_bot_bl2[3] bcconn_bot_bl2_n[3] bl1 bl1_n bl2 bl2_n bcconn_bot_bl1[5] bcconn_bot_bl1_n[5] bcconn_bot_bl2[5] bcconn_bot_bl2_n[5] bcconn_bot_bl1[6] bcconn_bot_bl1_n[6] bcconn_bot_bl2[6] bcconn_bot_bl2_n[6] bcconn_bot_bl1[7] bcconn_bot_bl1_n[7] bcconn_bot_bl2[7] bcconn_bot_bl2_n[7] DP8TVar1BulkConnRow_8
Xbcconn_top vss vdd bcconn_top_bl1[0] bcconn_top_bl1_n[0] bcconn_top_bl2[0] bcconn_top_bl2_n[0] bcconn_top_bl1[1] bcconn_top_bl1_n[1] bcconn_top_bl2[1] bcconn_top_bl2_n[1] bcconn_top_bl1[2] bcconn_top_bl1_n[2] bcconn_top_bl2[2] bcconn_top_bl2_n[2] bcconn_top_bl1[3] bcconn_top_bl1_n[3] bcconn_top_bl2[3] bcconn_top_bl2_n[3] bl1 bl1_n bl2 bl2_n bcconn_top_bl1[5] bcconn_top_bl1_n[5] bcconn_top_bl2[5] bcconn_top_bl2_n[5] bcconn_top_bl1[6] bcconn_top_bl1_n[6] bcconn_top_bl2[6] bcconn_top_bl2_n[6] bcconn_top_bl1[7] bcconn_top_bl1_n[7] bcconn_top_bl2[7] bcconn_top_bl2_n[7] DP8TVar1BulkConnRow_8
Xarray_bot vss vdd zero zero zero zero zero zero zero zero zero zero zero zero zero zero array_bot_bl1[0] array_bot_bl1_n[0] array_bot_bl2[0] array_bot_bl2_n[0] array_bot_bl1[1] array_bot_bl1_n[1] array_bot_bl2[1] array_bot_bl2_n[1] array_bot_bl1[2] array_bot_bl1_n[2] array_bot_bl2[2] array_bot_bl2_n[2] array_bot_bl1[3] array_bot_bl1_n[3] array_bot_bl2[3] array_bot_bl2_n[3] bl1 bl1_n bl2 bl2_n array_bot_bl1[5] array_bot_bl1_n[5] array_bot_bl2[5] array_bot_bl2_n[5] array_bot_bl1[6] array_bot_bl1_n[6] array_bot_bl2[6] array_bot_bl2_n[6] array_bot_bl1[7] array_bot_bl1_n[7] array_bot_bl2[7] array_bot_bl2_n[7] DP8TVar1Array_7X8
Xshwl1_row vss vdd zero bit shwl1_row_bl1[0] shwl1_row_bl1_n[0] shwl1_row_bl2[0] shwl1_row_bl2_n[0] shwl1_row_bl1[1] shwl1_row_bl1_n[1] shwl1_row_bl2[1] shwl1_row_bl2_n[1] shwl1_row_bl1[2] shwl1_row_bl1_n[2] shwl1_row_bl2[2] shwl1_row_bl2_n[2] shwl1_row_bl1[3] shwl1_row_bl1_n[3] shwl1_row_bl2[3] shwl1_row_bl2_n[3] bl1 bl1_n bl2 bl2_n shwl1_row_bl1[5] shwl1_row_bl1_n[5] shwl1_row_bl2[5] shwl1_row_bl2_n[5] shwl1_row_bl1[6] shwl1_row_bl1_n[6] shwl1_row_bl2[6] shwl1_row_bl2_n[6] shwl1_row_bl1[7] shwl1_row_bl1_n[7] shwl1_row_bl2[7] shwl1_row_bl2_n[7] DP8TVar1ArrayShWL1_1X8
Xcell_cols_left vss vdd wl1 wl2 cell_cols_left_bl1[0] cell_cols_left_bl1_n[0] cell_cols_left_bl2[0] cell_cols_left_bl2_n[0] cell_cols_left_bl1[1] cell_cols_left_bl1_n[1] cell_cols_left_bl2[1] cell_cols_left_bl2_n[1] cell_cols_left_bl1[2] cell_cols_left_bl1_n[2] cell_cols_left_bl2[2] cell_cols_left_bl2_n[2] cell_cols_left_bl1[3] cell_cols_left_bl1_n[3] cell_cols_left_bl2[3] cell_cols_left_bl2_n[3] DP8TVar1Array_1X4
Xconncell wl1 wl2 bl1 bl1_n bl2 bl2_n vdd vss bit bit_n DP8TVar1CellConnectOut
Xfillcell wl1 wl2 fillcell_bl1 fillcell_bl1_n fillcell_bl2 fillcell_bl2_n vdd vss DP8TVar1Cell
Xcell_cols_right vss vdd wl1 wl2 cell_cols_right_bl1[0] cell_cols_right_bl1_n[0] cell_cols_right_bl2[0] cell_cols_right_bl2_n[0] cell_cols_right_bl1[1] cell_cols_right_bl1_n[1] cell_cols_right_bl2[1] cell_cols_right_bl2_n[1] DP8TVar1Array_1X2
Xshwl2_row vss vdd bit_n zero shwl2_row_bl1[0] shwl2_row_bl1_n[0] shwl2_row_bl2[0] shwl2_row_bl2_n[0] shwl2_row_bl1[1] shwl2_row_bl1_n[1] shwl2_row_bl2[1] shwl2_row_bl2_n[1] shwl2_row_bl1[2] shwl2_row_bl1_n[2] shwl2_row_bl2[2] shwl2_row_bl2_n[2] shwl2_row_bl1[3] shwl2_row_bl1_n[3] shwl2_row_bl2[3] shwl2_row_bl2_n[3] bl1 bl1_n bl2 bl2_n shwl2_row_bl1[5] shwl2_row_bl1_n[5] shwl2_row_bl2[5] shwl2_row_bl2_n[5] shwl2_row_bl1[6] shwl2_row_bl1_n[6] shwl2_row_bl2[6] shwl2_row_bl2_n[6] shwl2_row_bl1[7] shwl2_row_bl1_n[7] shwl2_row_bl2[7] shwl2_row_bl2_n[7] DP8TVar1ArrayShWL2_1X8
Xarray_top vss vdd zero zero zero zero zero zero zero zero zero zero zero zero array_top_bl1[0] array_top_bl1_n[0] array_top_bl2[0] array_top_bl2_n[0] array_top_bl1[1] array_top_bl1_n[1] array_top_bl2[1] array_top_bl2_n[1] array_top_bl1[2] array_top_bl1_n[2] array_top_bl2[2] array_top_bl2_n[2] array_top_bl1[3] array_top_bl1_n[3] array_top_bl2[3] array_top_bl2_n[3] bl1 bl1_n bl2 bl2_n array_top_bl1[5] array_top_bl1_n[5] array_top_bl2[5] array_top_bl2_n[5] array_top_bl1[6] array_top_bl1_n[6] array_top_bl2[6] array_top_bl2_n[6] array_top_bl1[7] array_top_bl1_n[7] array_top_bl2[7] array_top_bl2_n[7] DP8TVar1Array_6X8
Xzero vdd vss zero zero_x1
.ends DP8TVar1TestArray_16X8C

.subckt PadFrame_DP01 PAD0x0 PAD0x1 PAD0x2 PAD0x3 PAD0x4 PAD0x5 PAD0x6 PAD0x7 PAD0x8 PAD0x9 PAD1x0 PAD1x1 PAD1x2 PAD1x3 PAD1x4 PAD1x5 PAD1x6 PAD1x7 PAD1x8 PAD1x9
XPAD0x0 PAD0x0 BondPad
XPAD0x1 PAD0x1 BondPad
XPAD0x2 PAD0x2 BondPad
XPAD0x3 PAD0x3 BondPad
XPAD0x4 PAD0x4 BondPad
XPAD0x5 PAD0x5 BondPad
XPAD0x6 PAD0x6 BondPad
XPAD0x7 PAD0x7 BondPad
XPAD0x8 PAD0x8 BondPad
XPAD0x9 PAD0x9 BondPad
XPAD1x0 PAD1x0 BondPad
XPAD1x1 PAD1x1 BondPad
XPAD1x2 PAD1x2 BondPad
XPAD1x3 PAD1x3 BondPad
XPAD1x4 PAD1x4 BondPad
XPAD1x5 PAD1x5 BondPad
XPAD1x6 PAD1x6 BondPad
XPAD1x7 PAD1x7 BondPad
XPAD1x8 PAD1x8 BondPad
XPAD1x9 PAD1x9 BondPad
.ends PadFrame_DP01

.subckt DP8TVar1 vss noco_vdd noco_wl1 noco_wl2 noco_bl1 noco_bl1_n noco_bl2 noco_bl2_n co_vdd co_bit co_bit_n co_wl1 co_wl2 co_bl1 co_bl1_n co_bl2_n co_bl2
Xframe noco_vdd noco_wl1 noco_wl2 noco_bl2 co_vdd co_bit co_bit_n co_wl1 co_wl2 NoConn_PAD0x9 vss noco_bl1 noco_bl1_n noco_bl2_n vss co_bl1 co_bl1_n co_bl2_n co_bl2 NoConn_PAD1x9 PadFrame_DP01
Xtestarray_noco vss noco_vdd noco_wl1 noco_wl2 noco_bl1 noco_bl1_n noco_bl2 noco_bl2_n DP8TVar1TestArray_16X8
Xtestarray_co vss co_vdd co_wl1 co_wl2 co_bl1 co_bl1_n co_bl2 co_bl2_n co_bit co_bit_n DP8TVar1TestArray_16X8C
.ends DP8TVar1

.subckt SP6TVar2Cell wl bl bl_n vdd vss
Xpu1 vdd bit_n bit vdd sg13_lv_pmos l=1.3e-07 w=1.5e-07
Xpd1 bit bit_n vss vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpu2 vdd bit bit_n vdd sg13_lv_pmos l=1.3e-07 w=1.5e-07
Xpd2 bit_n bit vss vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg1 bit wl bl vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg2 bit_n wl bl_n vss sg13_lv_nmos l=1.3e-07 w=3e-07
.ends SP6TVar2Cell

.subckt SP6TVar2Array_2X1 vss vdd wl[0] wl[1] bl[0] bl_n[0]
Xinst0x0 wl[0] bl[0] bl_n[0] vdd vss SP6TVar2Cell
Xinst1x0 wl[1] bl[0] bl_n[0] vdd vss SP6TVar2Cell
.ends SP6TVar2Array_2X1

.subckt SP6TVar2Array_2X2 vss vdd wl[0] wl[1] bl[0] bl_n[0] bl[1] bl_n[1]
Xinst0x0 vss vdd wl[0] wl[1] bl[0] bl_n[0] SP6TVar2Array_2X1
Xinst0x1 vss vdd wl[0] wl[1] bl[1] bl_n[1] SP6TVar2Array_2X1
.ends SP6TVar2Array_2X2

.subckt SP6TVar2Array_4X2 vss vdd wl[0] wl[1] wl[2] wl[3] bl[0] bl_n[0] bl[1] bl_n[1]
Xinst0x0 vss vdd wl[0] wl[1] bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar2Array_2X2
Xinst1x0 vss vdd wl[2] wl[3] bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar2Array_2X2
.ends SP6TVar2Array_4X2

.subckt SP6TVar2Array_4X4 vss vdd wl[0] wl[1] wl[2] wl[3] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar2Array_4X2
Xinst0x1 vss vdd wl[0] wl[1] wl[2] wl[3] bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar2Array_4X2
.ends SP6TVar2Array_4X4

.subckt SP6TVar2Array_8X4 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar2Array_4X4
Xinst1x0 vss vdd wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar2Array_4X4
.ends SP6TVar2Array_8X4

.subckt SP6TVar2Array_8X8 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar2Array_8X4
Xinst0x1 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7] SP6TVar2Array_8X4
.ends SP6TVar2Array_8X8

.subckt SP6TVar2BulkConn vdd vss bl bl_n
.ends SP6TVar2BulkConn

.subckt SP6TVar2BulkConnRow_2 vss vdd bl[0] bl_n[0] bl[1] bl_n[1]
Xinst0 vdd vss bl[0] bl_n[0] SP6TVar2BulkConn
Xinst1 vdd vss bl[1] bl_n[1] SP6TVar2BulkConn
.ends SP6TVar2BulkConnRow_2

.subckt SP6TVar2BulkConnRow_4 vss vdd bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3]
Xinst0 vss vdd bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar2BulkConnRow_2
Xinst1 vss vdd bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar2BulkConnRow_2
.ends SP6TVar2BulkConnRow_4

.subckt SP6TVar2BulkConnRow_8 vss vdd bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7]
Xinst0 vss vdd bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar2BulkConnRow_4
Xinst1 vss vdd bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7] SP6TVar2BulkConnRow_4
.ends SP6TVar2BulkConnRow_8

.subckt SP6TVar2Array_16X8BC vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7] SP6TVar2Array_8X8
Xinst1x0 vss vdd wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7] SP6TVar2Array_8X8
Xbottombcrow vss vdd bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7] SP6TVar2BulkConnRow_8
Xtopbcrow vss vdd bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7] SP6TVar2BulkConnRow_8
.ends SP6TVar2Array_16X8BC

.subckt SP6TVar2TestArray_16X8 vss vdd bl bl_n wl
Xarray vss vdd zero zero zero zero zero zero zero zero wl zero zero zero zero zero zero zero bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl bl_n bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7] SP6TVar2Array_16X8BC
Xzero vdd vss zero zero_x1
.ends SP6TVar2TestArray_16X8

.subckt SP6TVar2Array_4X1 vss vdd wl[0] wl[1] wl[2] wl[3] bl[0] bl_n[0]
Xinst0x0 vss vdd wl[0] wl[1] bl[0] bl_n[0] SP6TVar2Array_2X1
Xinst1x0 vss vdd wl[2] wl[3] bl[0] bl_n[0] SP6TVar2Array_2X1
.ends SP6TVar2Array_4X1

.subckt SP6TVar2Array_8X1 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] bl[0] bl_n[0] SP6TVar2Array_4X1
Xinst1x0 vss vdd wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] SP6TVar2Array_4X1
.ends SP6TVar2Array_8X1

.subckt SP6TVar2Array_16X1BC vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] bl[0] bl_n[0]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] SP6TVar2Array_8X1
Xinst1x0 vss vdd wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] bl[0] bl_n[0] SP6TVar2Array_8X1
Xbottombcrow vdd vss bl[0] bl_n[0] SP6TVar2BulkConn
Xtopbcrow vdd vss bl[0] bl_n[0] SP6TVar2BulkConn
.ends SP6TVar2Array_16X1BC

.subckt SP6TVar2Array_8X2 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar2Array_4X2
Xinst1x0 vss vdd wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar2Array_4X2
.ends SP6TVar2Array_8X2

.subckt SP6TVar2Array_16X2BC vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] bl[0] bl_n[0] bl[1] bl_n[1]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar2Array_8X2
Xinst1x0 vss vdd wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar2Array_8X2
Xbottombcrow vss vdd bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar2BulkConnRow_2
Xtopbcrow vss vdd bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar2BulkConnRow_2
.ends SP6TVar2Array_16X2BC

.subckt SP6TVar2Array_16X4BC vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar2Array_8X4
Xinst1x0 vss vdd wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar2Array_8X4
Xbottombcrow vss vdd bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar2BulkConnRow_4
Xtopbcrow vss vdd bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar2BulkConnRow_4
.ends SP6TVar2Array_16X4BC

.subckt SP6TVar2Array_6X1 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] bl[0] bl_n[0]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] bl[0] bl_n[0] SP6TVar2Array_4X1
Xinst1x0 vss vdd wl[4] wl[5] bl[0] bl_n[0] SP6TVar2Array_2X1
.ends SP6TVar2Array_6X1

.subckt SP6TVar2CellConnectOut wl bl bl_n vdd vss bit bit_n
Xpu1 vdd bit_n bit vdd sg13_lv_pmos l=1.3e-07 w=1.5e-07
Xpd1 bit bit_n vss vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpu2 vdd bit bit_n vdd sg13_lv_pmos l=1.3e-07 w=1.5e-07
Xpd2 bit_n bit vss vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg1 bit wl bl vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg2 bit_n wl bl_n vss sg13_lv_nmos l=1.3e-07 w=3e-07
.ends SP6TVar2CellConnectOut

.subckt SP6TVar2TestArray_16X8C vss vdd bl bl_n bit bit_n wl
Xarray_0 vss vdd zero zero zero zero zero zero zero zero wl zero zero zero zero zero zero zero array_0_bl[0] array_0_bl_n[0] SP6TVar2Array_16X1BC
Xarray_1 vss vdd zero zero zero zero zero zero zero zero wl zero zero zero zero zero zero zero array_1_bl[0] array_1_bl_n[0] array_1_bl[1] array_1_bl_n[1] SP6TVar2Array_16X2BC
Xarray_2 vss vdd zero zero zero zero zero zero zero zero wl zero zero zero zero zero zero zero array_2_bl[0] array_2_bl_n[0] array_2_bl[1] array_2_bl_n[1] array_2_bl[2] array_2_bl_n[2] array_2_bl[3] array_2_bl_n[3] SP6TVar2Array_16X4BC
Xcolbc_0 vdd vss bl bl_n SP6TVar2BulkConn
Xcolbc_1 vdd vss bl bl_n SP6TVar2BulkConn
Xcolarray_0 vss vdd zero zero zero zero zero zero zero zero bl bl_n SP6TVar2Array_8X1
Xcolarray_1 vss vdd zero zero zero zero zero zero bl bl_n SP6TVar2Array_6X1
Xbc_noconn zero bl bl_n vdd vss SP6TVar2Cell
Xbc_conn wl bl bl_n vdd vss bit bit_n SP6TVar2CellConnectOut
Xzero vdd vss zero zero_x1
.ends SP6TVar2TestArray_16X8C

.subckt PadFrame_SP02 PAD0x0 PAD0x1 PAD0x2 PAD0x3 PAD0x4 PAD0x5 PAD0x6 PAD0x7 PAD0x8 PAD0x9 PAD1x0 PAD1x1 PAD1x2 PAD1x3 PAD1x4 PAD1x5 PAD1x6 PAD1x7 PAD1x8 PAD1x9
XPAD0x0 PAD0x0 BondPad
XPAD0x1 PAD0x1 BondPad
XPAD0x2 PAD0x2 BondPad
XPAD0x3 PAD0x3 BondPad
XPAD0x4 PAD0x4 BondPad
XPAD0x5 PAD0x5 BondPad
XPAD0x6 PAD0x6 BondPad
XPAD0x7 PAD0x7 BondPad
XPAD0x8 PAD0x8 BondPad
XPAD0x9 PAD0x9 BondPad
XPAD1x0 PAD1x0 BondPad
XPAD1x1 PAD1x1 BondPad
XPAD1x2 PAD1x2 BondPad
XPAD1x3 PAD1x3 BondPad
XPAD1x4 PAD1x4 BondPad
XPAD1x5 PAD1x5 BondPad
XPAD1x6 PAD1x6 BondPad
XPAD1x7 PAD1x7 BondPad
XPAD1x8 PAD1x8 BondPad
XPAD1x9 PAD1x9 BondPad
.ends PadFrame_SP02

.subckt SP6TVar2 vss noco_vdd noco_wl noco_bl noco_bl_n co_vdd co_bl co_bl_n co_bit co_bit_n co_wl
Xframe noco_vdd noco_wl NoConn_PAD0x2 co_vdd co_bl_n co_bit co_bit_n NoConn_PAD0x7 NoConn_PAD0x8 NoConn_PAD0x9 vss noco_bl noco_bl_n vss co_bl co_wl NoConn_PAD1x6 NoConn_PAD1x7 NoConn_PAD1x8 NoConn_PAD1x9 PadFrame_SP02
Xtestarray_noco vss noco_vdd noco_bl noco_bl_n noco_wl SP6TVar2TestArray_16X8
Xtestarray_co vss co_vdd co_bl co_bl_n co_bit co_bit_n co_wl SP6TVar2TestArray_16X8C
.ends SP6TVar2

.subckt DP8TVar2Cell wl1 wl2 bl1 bl1_n bl2 bl2_n vdd vss
Xpu1 vdd bit_n bit vdd sg13_lv_pmos l=1.3e-07 w=1.5e-07
Xpd1 bit bit_n vss vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpu2 vdd bit bit_n vdd sg13_lv_pmos l=1.3e-07 w=1.5e-07
Xpd2 bit_n bit vss vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg1 bit wl1 bl1 vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg1n bit_n wl1 bl1_n vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg2 bit wl2 bl2 vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg2n bit_n wl2 bl2_n vss sg13_lv_nmos l=1.3e-07 w=3e-07
.ends DP8TVar2Cell

.subckt DP8TVar2Array_2X1 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0]
Xinst0x0 wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] vdd vss DP8TVar2Cell
Xinst1x0 wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0] vdd vss DP8TVar2Cell
.ends DP8TVar2Array_2X1

.subckt DP8TVar2Array_2X2 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0] DP8TVar2Array_2X1
Xinst0x1 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TVar2Array_2X1
.ends DP8TVar2Array_2X2

.subckt DP8TVar2Array_4X2 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TVar2Array_2X2
Xinst1x0 vss vdd wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TVar2Array_2X2
.ends DP8TVar2Array_4X2

.subckt DP8TVar2Array_4X4 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TVar2Array_4X2
Xinst0x1 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar2Array_4X2
.ends DP8TVar2Array_4X4

.subckt DP8TVar2Array_8X4 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar2Array_4X4
Xinst1x0 vss vdd wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar2Array_4X4
.ends DP8TVar2Array_8X4

.subckt DP8TVar2Array_8X8 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar2Array_8X4
Xinst0x1 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar2Array_8X4
.ends DP8TVar2Array_8X8

.subckt DP8TVar2BulkConn vdd vss bl1 bl2 bl1_n bl2_n
.ends DP8TVar2BulkConn

.subckt DP8TVar2BulkConnRow_2 vss vdd bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1]
Xinst0 vdd vss bl1[0] bl2[0] bl1_n[0] bl2_n[0] DP8TVar2BulkConn
Xinst1 vdd vss bl1[1] bl2[1] bl1_n[1] bl2_n[1] DP8TVar2BulkConn
.ends DP8TVar2BulkConnRow_2

.subckt DP8TVar2BulkConnRow_4 vss vdd bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3]
Xinst0 vss vdd bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TVar2BulkConnRow_2
Xinst1 vss vdd bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar2BulkConnRow_2
.ends DP8TVar2BulkConnRow_4

.subckt DP8TVar2BulkConnRow_8 vss vdd bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0 vss vdd bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar2BulkConnRow_4
Xinst1 vss vdd bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar2BulkConnRow_4
.ends DP8TVar2BulkConnRow_8

.subckt DP8TVar2Array_16X8BC vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] wl1[8] wl2[8] wl1[9] wl2[9] wl1[10] wl2[10] wl1[11] wl2[11] wl1[12] wl2[12] wl1[13] wl2[13] wl1[14] wl2[14] wl1[15] wl2[15] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar2Array_8X8
Xinst1x0 vss vdd wl1[8] wl2[8] wl1[9] wl2[9] wl1[10] wl2[10] wl1[11] wl2[11] wl1[12] wl2[12] wl1[13] wl2[13] wl1[14] wl2[14] wl1[15] wl2[15] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar2Array_8X8
Xbottombcrow vss vdd bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar2BulkConnRow_8
Xtopbcrow vss vdd bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar2BulkConnRow_8
.ends DP8TVar2Array_16X8BC

.subckt DP8TVar2TestArray_16X8 vss vdd wl1 wl2 bl1 bl1_n bl2 bl2_n
Xarray vss vdd zero zero zero zero zero zero zero zero zero zero zero zero zero zero zero zero wl1 wl2 zero zero zero zero zero zero zero zero zero zero zero zero zero zero bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1 bl1_n bl2 bl2_n bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar2Array_16X8BC
Xzero vdd vss zero zero_x1
.ends DP8TVar2TestArray_16X8

.subckt DP8TVar2Array_4X8 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar2Array_4X4
Xinst0x1 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar2Array_4X4
.ends DP8TVar2Array_4X8

.subckt DP8TVar2Array_2X4 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TVar2Array_2X2
Xinst0x1 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar2Array_2X2
.ends DP8TVar2Array_2X4

.subckt DP8TVar2Array_2X8 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar2Array_2X4
Xinst0x1 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar2Array_2X4
.ends DP8TVar2Array_2X8

.subckt DP8TVar2Array_1X2 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1]
Xinst0x0 wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] vdd vss DP8TVar2Cell
Xinst0x1 wl1[0] wl2[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] vdd vss DP8TVar2Cell
.ends DP8TVar2Array_1X2

.subckt DP8TVar2Array_1X4 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3]
Xinst0x0 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TVar2Array_1X2
Xinst0x1 vss vdd wl1[0] wl2[0] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar2Array_1X2
.ends DP8TVar2Array_1X4

.subckt DP8TVar2Array_1X8 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar2Array_1X4
Xinst0x1 vss vdd wl1[0] wl2[0] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar2Array_1X4
.ends DP8TVar2Array_1X8

.subckt DP8TVar2Array_7X8 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar2Array_4X8
Xinst1x0 vss vdd wl1[4] wl2[4] wl1[5] wl2[5] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar2Array_2X8
Xinst2x0 vss vdd wl1[6] wl2[6] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar2Array_1X8
.ends DP8TVar2Array_7X8

.subckt DP8TVar2CellShWL1 wl1 wl2 bl1 bl1_n bl2 bl2_n vdd vss
Xpu1 vdd bit_n bit vdd sg13_lv_pmos l=1.3e-07 w=1.5e-07
Xpd1 bit bit_n vss vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpu2 vdd bit bit_n vdd sg13_lv_pmos l=1.3e-07 w=1.5e-07
Xpd2 bit_n bit vss vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg1 bit wl1 bl1 vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg1n bit_n wl1 bl1_n vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg2 bit wl1 bl2 vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg2n bit_n wl1 bl2_n vss sg13_lv_nmos l=1.3e-07 w=3e-07
.ends DP8TVar2CellShWL1

.subckt DP8TVar2ArrayShWL1_1X2 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1]
Xinst0x0 wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] vdd vss DP8TVar2CellShWL1
Xinst0x1 wl1[0] wl2[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] vdd vss DP8TVar2CellShWL1
.ends DP8TVar2ArrayShWL1_1X2

.subckt DP8TVar2ArrayShWL1_1X4 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3]
Xinst0x0 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TVar2ArrayShWL1_1X2
Xinst0x1 vss vdd wl1[0] wl2[0] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar2ArrayShWL1_1X2
.ends DP8TVar2ArrayShWL1_1X4

.subckt DP8TVar2ArrayShWL1_1X8 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar2ArrayShWL1_1X4
Xinst0x1 vss vdd wl1[0] wl2[0] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar2ArrayShWL1_1X4
.ends DP8TVar2ArrayShWL1_1X8

.subckt DP8TVar2CellConnectOut wl1 wl2 bl1 bl1_n bl2 bl2_n vdd vss bit bit_n
Xpu1 vdd bit_n bit vdd sg13_lv_pmos l=1.3e-07 w=1.5e-07
Xpd1 bit bit_n vss vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpu2 vdd bit bit_n vdd sg13_lv_pmos l=1.3e-07 w=1.5e-07
Xpd2 bit_n bit vss vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg1 bit wl1 bl1 vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg1n bit_n wl1 bl1_n vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg2 bit wl2 bl2 vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg2n bit_n wl2 bl2_n vss sg13_lv_nmos l=1.3e-07 w=3e-07
.ends DP8TVar2CellConnectOut

.subckt DP8TVar2CellShWL2 wl1 wl2 bl1 bl1_n bl2 bl2_n vdd vss
Xpu1 vdd bit_n bit vdd sg13_lv_pmos l=1.3e-07 w=1.5e-07
Xpd1 bit bit_n vss vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpu2 vdd bit bit_n vdd sg13_lv_pmos l=1.3e-07 w=1.5e-07
Xpd2 bit_n bit vss vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg1 bit wl2 bl1 vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg1n bit_n wl2 bl1_n vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg2 bit wl2 bl2 vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg2n bit_n wl2 bl2_n vss sg13_lv_nmos l=1.3e-07 w=3e-07
.ends DP8TVar2CellShWL2

.subckt DP8TVar2ArrayShWL2_1X2 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1]
Xinst0x0 wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] vdd vss DP8TVar2CellShWL2
Xinst0x1 wl1[0] wl2[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] vdd vss DP8TVar2CellShWL2
.ends DP8TVar2ArrayShWL2_1X2

.subckt DP8TVar2ArrayShWL2_1X4 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3]
Xinst0x0 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TVar2ArrayShWL2_1X2
Xinst0x1 vss vdd wl1[0] wl2[0] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar2ArrayShWL2_1X2
.ends DP8TVar2ArrayShWL2_1X4

.subckt DP8TVar2ArrayShWL2_1X8 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar2ArrayShWL2_1X4
Xinst0x1 vss vdd wl1[0] wl2[0] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar2ArrayShWL2_1X4
.ends DP8TVar2ArrayShWL2_1X8

.subckt DP8TVar2Array_6X8 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar2Array_4X8
Xinst1x0 vss vdd wl1[4] wl2[4] wl1[5] wl2[5] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar2Array_2X8
.ends DP8TVar2Array_6X8

.subckt DP8TVar2TestArray_16X8C vss vdd wl1 wl2 bl1 bl1_n bl2 bl2_n bit bit_n
Xbcconn_bot vss vdd bcconn_bot_bl1[0] bcconn_bot_bl1_n[0] bcconn_bot_bl2[0] bcconn_bot_bl2_n[0] bcconn_bot_bl1[1] bcconn_bot_bl1_n[1] bcconn_bot_bl2[1] bcconn_bot_bl2_n[1] bcconn_bot_bl1[2] bcconn_bot_bl1_n[2] bcconn_bot_bl2[2] bcconn_bot_bl2_n[2] bcconn_bot_bl1[3] bcconn_bot_bl1_n[3] bcconn_bot_bl2[3] bcconn_bot_bl2_n[3] bl1 bl1_n bl2 bl2_n bcconn_bot_bl1[5] bcconn_bot_bl1_n[5] bcconn_bot_bl2[5] bcconn_bot_bl2_n[5] bcconn_bot_bl1[6] bcconn_bot_bl1_n[6] bcconn_bot_bl2[6] bcconn_bot_bl2_n[6] bcconn_bot_bl1[7] bcconn_bot_bl1_n[7] bcconn_bot_bl2[7] bcconn_bot_bl2_n[7] DP8TVar2BulkConnRow_8
Xbcconn_top vss vdd bcconn_top_bl1[0] bcconn_top_bl1_n[0] bcconn_top_bl2[0] bcconn_top_bl2_n[0] bcconn_top_bl1[1] bcconn_top_bl1_n[1] bcconn_top_bl2[1] bcconn_top_bl2_n[1] bcconn_top_bl1[2] bcconn_top_bl1_n[2] bcconn_top_bl2[2] bcconn_top_bl2_n[2] bcconn_top_bl1[3] bcconn_top_bl1_n[3] bcconn_top_bl2[3] bcconn_top_bl2_n[3] bl1 bl1_n bl2 bl2_n bcconn_top_bl1[5] bcconn_top_bl1_n[5] bcconn_top_bl2[5] bcconn_top_bl2_n[5] bcconn_top_bl1[6] bcconn_top_bl1_n[6] bcconn_top_bl2[6] bcconn_top_bl2_n[6] bcconn_top_bl1[7] bcconn_top_bl1_n[7] bcconn_top_bl2[7] bcconn_top_bl2_n[7] DP8TVar2BulkConnRow_8
Xarray_bot vss vdd zero zero zero zero zero zero zero zero zero zero zero zero zero zero array_bot_bl1[0] array_bot_bl1_n[0] array_bot_bl2[0] array_bot_bl2_n[0] array_bot_bl1[1] array_bot_bl1_n[1] array_bot_bl2[1] array_bot_bl2_n[1] array_bot_bl1[2] array_bot_bl1_n[2] array_bot_bl2[2] array_bot_bl2_n[2] array_bot_bl1[3] array_bot_bl1_n[3] array_bot_bl2[3] array_bot_bl2_n[3] bl1 bl1_n bl2 bl2_n array_bot_bl1[5] array_bot_bl1_n[5] array_bot_bl2[5] array_bot_bl2_n[5] array_bot_bl1[6] array_bot_bl1_n[6] array_bot_bl2[6] array_bot_bl2_n[6] array_bot_bl1[7] array_bot_bl1_n[7] array_bot_bl2[7] array_bot_bl2_n[7] DP8TVar2Array_7X8
Xshwl1_row vss vdd zero bit shwl1_row_bl1[0] shwl1_row_bl1_n[0] shwl1_row_bl2[0] shwl1_row_bl2_n[0] shwl1_row_bl1[1] shwl1_row_bl1_n[1] shwl1_row_bl2[1] shwl1_row_bl2_n[1] shwl1_row_bl1[2] shwl1_row_bl1_n[2] shwl1_row_bl2[2] shwl1_row_bl2_n[2] shwl1_row_bl1[3] shwl1_row_bl1_n[3] shwl1_row_bl2[3] shwl1_row_bl2_n[3] bl1 bl1_n bl2 bl2_n shwl1_row_bl1[5] shwl1_row_bl1_n[5] shwl1_row_bl2[5] shwl1_row_bl2_n[5] shwl1_row_bl1[6] shwl1_row_bl1_n[6] shwl1_row_bl2[6] shwl1_row_bl2_n[6] shwl1_row_bl1[7] shwl1_row_bl1_n[7] shwl1_row_bl2[7] shwl1_row_bl2_n[7] DP8TVar2ArrayShWL1_1X8
Xcell_cols_left vss vdd wl1 wl2 cell_cols_left_bl1[0] cell_cols_left_bl1_n[0] cell_cols_left_bl2[0] cell_cols_left_bl2_n[0] cell_cols_left_bl1[1] cell_cols_left_bl1_n[1] cell_cols_left_bl2[1] cell_cols_left_bl2_n[1] cell_cols_left_bl1[2] cell_cols_left_bl1_n[2] cell_cols_left_bl2[2] cell_cols_left_bl2_n[2] cell_cols_left_bl1[3] cell_cols_left_bl1_n[3] cell_cols_left_bl2[3] cell_cols_left_bl2_n[3] DP8TVar2Array_1X4
Xconncell wl1 wl2 bl1 bl1_n bl2 bl2_n vdd vss bit bit_n DP8TVar2CellConnectOut
Xfillcell wl1 wl2 fillcell_bl1 fillcell_bl1_n fillcell_bl2 fillcell_bl2_n vdd vss DP8TVar2Cell
Xcell_cols_right vss vdd wl1 wl2 cell_cols_right_bl1[0] cell_cols_right_bl1_n[0] cell_cols_right_bl2[0] cell_cols_right_bl2_n[0] cell_cols_right_bl1[1] cell_cols_right_bl1_n[1] cell_cols_right_bl2[1] cell_cols_right_bl2_n[1] DP8TVar2Array_1X2
Xshwl2_row vss vdd bit_n zero shwl2_row_bl1[0] shwl2_row_bl1_n[0] shwl2_row_bl2[0] shwl2_row_bl2_n[0] shwl2_row_bl1[1] shwl2_row_bl1_n[1] shwl2_row_bl2[1] shwl2_row_bl2_n[1] shwl2_row_bl1[2] shwl2_row_bl1_n[2] shwl2_row_bl2[2] shwl2_row_bl2_n[2] shwl2_row_bl1[3] shwl2_row_bl1_n[3] shwl2_row_bl2[3] shwl2_row_bl2_n[3] bl1 bl1_n bl2 bl2_n shwl2_row_bl1[5] shwl2_row_bl1_n[5] shwl2_row_bl2[5] shwl2_row_bl2_n[5] shwl2_row_bl1[6] shwl2_row_bl1_n[6] shwl2_row_bl2[6] shwl2_row_bl2_n[6] shwl2_row_bl1[7] shwl2_row_bl1_n[7] shwl2_row_bl2[7] shwl2_row_bl2_n[7] DP8TVar2ArrayShWL2_1X8
Xarray_top vss vdd zero zero zero zero zero zero zero zero zero zero zero zero array_top_bl1[0] array_top_bl1_n[0] array_top_bl2[0] array_top_bl2_n[0] array_top_bl1[1] array_top_bl1_n[1] array_top_bl2[1] array_top_bl2_n[1] array_top_bl1[2] array_top_bl1_n[2] array_top_bl2[2] array_top_bl2_n[2] array_top_bl1[3] array_top_bl1_n[3] array_top_bl2[3] array_top_bl2_n[3] bl1 bl1_n bl2 bl2_n array_top_bl1[5] array_top_bl1_n[5] array_top_bl2[5] array_top_bl2_n[5] array_top_bl1[6] array_top_bl1_n[6] array_top_bl2[6] array_top_bl2_n[6] array_top_bl1[7] array_top_bl1_n[7] array_top_bl2[7] array_top_bl2_n[7] DP8TVar2Array_6X8
Xzero vdd vss zero zero_x1
.ends DP8TVar2TestArray_16X8C

.subckt PadFrame_DP02 PAD0x0 PAD0x1 PAD0x2 PAD0x3 PAD0x4 PAD0x5 PAD0x6 PAD0x7 PAD0x8 PAD0x9 PAD1x0 PAD1x1 PAD1x2 PAD1x3 PAD1x4 PAD1x5 PAD1x6 PAD1x7 PAD1x8 PAD1x9
XPAD0x0 PAD0x0 BondPad
XPAD0x1 PAD0x1 BondPad
XPAD0x2 PAD0x2 BondPad
XPAD0x3 PAD0x3 BondPad
XPAD0x4 PAD0x4 BondPad
XPAD0x5 PAD0x5 BondPad
XPAD0x6 PAD0x6 BondPad
XPAD0x7 PAD0x7 BondPad
XPAD0x8 PAD0x8 BondPad
XPAD0x9 PAD0x9 BondPad
XPAD1x0 PAD1x0 BondPad
XPAD1x1 PAD1x1 BondPad
XPAD1x2 PAD1x2 BondPad
XPAD1x3 PAD1x3 BondPad
XPAD1x4 PAD1x4 BondPad
XPAD1x5 PAD1x5 BondPad
XPAD1x6 PAD1x6 BondPad
XPAD1x7 PAD1x7 BondPad
XPAD1x8 PAD1x8 BondPad
XPAD1x9 PAD1x9 BondPad
.ends PadFrame_DP02

.subckt DP8TVar2 vss noco_vdd noco_wl1 noco_wl2 noco_bl1 noco_bl1_n noco_bl2 noco_bl2_n co_vdd co_bit co_bit_n co_wl1 co_wl2 co_bl1 co_bl1_n co_bl2_n co_bl2
Xframe noco_vdd noco_wl1 noco_wl2 noco_bl2 co_vdd co_bit co_bit_n co_wl1 co_wl2 NoConn_PAD0x9 vss noco_bl1 noco_bl1_n noco_bl2_n vss co_bl1 co_bl1_n co_bl2_n co_bl2 NoConn_PAD1x9 PadFrame_DP02
Xtestarray_noco vss noco_vdd noco_wl1 noco_wl2 noco_bl1 noco_bl1_n noco_bl2 noco_bl2_n DP8TVar2TestArray_16X8
Xtestarray_co vss co_vdd co_wl1 co_wl2 co_bl1 co_bl1_n co_bl2 co_bl2_n co_bit co_bit_n DP8TVar2TestArray_16X8C
.ends DP8TVar2

.subckt SP6TVar3Cell wl bl bl_n vdd vss
Xpu1 vdd bit_n bit vdd sg13_lv_pmos l=1.3e-07 w=2e-07
Xpd1 bit bit_n vss vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpu2 vdd bit bit_n vdd sg13_lv_pmos l=1.3e-07 w=2e-07
Xpd2 bit_n bit vss vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg1 bit wl bl vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg2 bit_n wl bl_n vss sg13_lv_nmos l=1.3e-07 w=2e-07
.ends SP6TVar3Cell

.subckt SP6TVar3Array_2X1 vss vdd wl[0] wl[1] bl[0] bl_n[0]
Xinst0x0 wl[0] bl[0] bl_n[0] vdd vss SP6TVar3Cell
Xinst1x0 wl[1] bl[0] bl_n[0] vdd vss SP6TVar3Cell
.ends SP6TVar3Array_2X1

.subckt SP6TVar3Array_2X2 vss vdd wl[0] wl[1] bl[0] bl_n[0] bl[1] bl_n[1]
Xinst0x0 vss vdd wl[0] wl[1] bl[0] bl_n[0] SP6TVar3Array_2X1
Xinst0x1 vss vdd wl[0] wl[1] bl[1] bl_n[1] SP6TVar3Array_2X1
.ends SP6TVar3Array_2X2

.subckt SP6TVar3Array_4X2 vss vdd wl[0] wl[1] wl[2] wl[3] bl[0] bl_n[0] bl[1] bl_n[1]
Xinst0x0 vss vdd wl[0] wl[1] bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar3Array_2X2
Xinst1x0 vss vdd wl[2] wl[3] bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar3Array_2X2
.ends SP6TVar3Array_4X2

.subckt SP6TVar3Array_4X4 vss vdd wl[0] wl[1] wl[2] wl[3] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar3Array_4X2
Xinst0x1 vss vdd wl[0] wl[1] wl[2] wl[3] bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar3Array_4X2
.ends SP6TVar3Array_4X4

.subckt SP6TVar3Array_8X4 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar3Array_4X4
Xinst1x0 vss vdd wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar3Array_4X4
.ends SP6TVar3Array_8X4

.subckt SP6TVar3Array_8X8 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar3Array_8X4
Xinst0x1 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7] SP6TVar3Array_8X4
.ends SP6TVar3Array_8X8

.subckt SP6TVar3BulkConn vdd vss bl bl_n
.ends SP6TVar3BulkConn

.subckt SP6TVar3BulkConnRow_2 vss vdd bl[0] bl_n[0] bl[1] bl_n[1]
Xinst0 vdd vss bl[0] bl_n[0] SP6TVar3BulkConn
Xinst1 vdd vss bl[1] bl_n[1] SP6TVar3BulkConn
.ends SP6TVar3BulkConnRow_2

.subckt SP6TVar3BulkConnRow_4 vss vdd bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3]
Xinst0 vss vdd bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar3BulkConnRow_2
Xinst1 vss vdd bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar3BulkConnRow_2
.ends SP6TVar3BulkConnRow_4

.subckt SP6TVar3BulkConnRow_8 vss vdd bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7]
Xinst0 vss vdd bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar3BulkConnRow_4
Xinst1 vss vdd bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7] SP6TVar3BulkConnRow_4
.ends SP6TVar3BulkConnRow_8

.subckt SP6TVar3Array_16X8BC vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7] SP6TVar3Array_8X8
Xinst1x0 vss vdd wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7] SP6TVar3Array_8X8
Xbottombcrow vss vdd bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7] SP6TVar3BulkConnRow_8
Xtopbcrow vss vdd bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7] SP6TVar3BulkConnRow_8
.ends SP6TVar3Array_16X8BC

.subckt SP6TVar3TestArray_16X8 vss vdd bl bl_n wl
Xarray vss vdd zero zero zero zero zero zero zero zero wl zero zero zero zero zero zero zero bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl bl_n bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7] SP6TVar3Array_16X8BC
Xzero vdd vss zero zero_x1
.ends SP6TVar3TestArray_16X8

.subckt SP6TVar3Array_4X1 vss vdd wl[0] wl[1] wl[2] wl[3] bl[0] bl_n[0]
Xinst0x0 vss vdd wl[0] wl[1] bl[0] bl_n[0] SP6TVar3Array_2X1
Xinst1x0 vss vdd wl[2] wl[3] bl[0] bl_n[0] SP6TVar3Array_2X1
.ends SP6TVar3Array_4X1

.subckt SP6TVar3Array_8X1 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] bl[0] bl_n[0] SP6TVar3Array_4X1
Xinst1x0 vss vdd wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] SP6TVar3Array_4X1
.ends SP6TVar3Array_8X1

.subckt SP6TVar3Array_16X1BC vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] bl[0] bl_n[0]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] SP6TVar3Array_8X1
Xinst1x0 vss vdd wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] bl[0] bl_n[0] SP6TVar3Array_8X1
Xbottombcrow vdd vss bl[0] bl_n[0] SP6TVar3BulkConn
Xtopbcrow vdd vss bl[0] bl_n[0] SP6TVar3BulkConn
.ends SP6TVar3Array_16X1BC

.subckt SP6TVar3Array_8X2 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar3Array_4X2
Xinst1x0 vss vdd wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar3Array_4X2
.ends SP6TVar3Array_8X2

.subckt SP6TVar3Array_16X2BC vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] bl[0] bl_n[0] bl[1] bl_n[1]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar3Array_8X2
Xinst1x0 vss vdd wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar3Array_8X2
Xbottombcrow vss vdd bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar3BulkConnRow_2
Xtopbcrow vss vdd bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar3BulkConnRow_2
.ends SP6TVar3Array_16X2BC

.subckt SP6TVar3Array_16X4BC vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar3Array_8X4
Xinst1x0 vss vdd wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar3Array_8X4
Xbottombcrow vss vdd bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar3BulkConnRow_4
Xtopbcrow vss vdd bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar3BulkConnRow_4
.ends SP6TVar3Array_16X4BC

.subckt SP6TVar3Array_6X1 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] bl[0] bl_n[0]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] bl[0] bl_n[0] SP6TVar3Array_4X1
Xinst1x0 vss vdd wl[4] wl[5] bl[0] bl_n[0] SP6TVar3Array_2X1
.ends SP6TVar3Array_6X1

.subckt SP6TVar3CellConnectOut wl bl bl_n vdd vss bit bit_n
Xpu1 vdd bit_n bit vdd sg13_lv_pmos l=1.3e-07 w=2e-07
Xpd1 bit bit_n vss vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpu2 vdd bit bit_n vdd sg13_lv_pmos l=1.3e-07 w=2e-07
Xpd2 bit_n bit vss vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg1 bit wl bl vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg2 bit_n wl bl_n vss sg13_lv_nmos l=1.3e-07 w=2e-07
.ends SP6TVar3CellConnectOut

.subckt SP6TVar3TestArray_16X8C vss vdd bl bl_n bit bit_n wl
Xarray_0 vss vdd zero zero zero zero zero zero zero zero wl zero zero zero zero zero zero zero array_0_bl[0] array_0_bl_n[0] SP6TVar3Array_16X1BC
Xarray_1 vss vdd zero zero zero zero zero zero zero zero wl zero zero zero zero zero zero zero array_1_bl[0] array_1_bl_n[0] array_1_bl[1] array_1_bl_n[1] SP6TVar3Array_16X2BC
Xarray_2 vss vdd zero zero zero zero zero zero zero zero wl zero zero zero zero zero zero zero array_2_bl[0] array_2_bl_n[0] array_2_bl[1] array_2_bl_n[1] array_2_bl[2] array_2_bl_n[2] array_2_bl[3] array_2_bl_n[3] SP6TVar3Array_16X4BC
Xcolbc_0 vdd vss bl bl_n SP6TVar3BulkConn
Xcolbc_1 vdd vss bl bl_n SP6TVar3BulkConn
Xcolarray_0 vss vdd zero zero zero zero zero zero zero zero bl bl_n SP6TVar3Array_8X1
Xcolarray_1 vss vdd zero zero zero zero zero zero bl bl_n SP6TVar3Array_6X1
Xbc_noconn zero bl bl_n vdd vss SP6TVar3Cell
Xbc_conn wl bl bl_n vdd vss bit bit_n SP6TVar3CellConnectOut
Xzero vdd vss zero zero_x1
.ends SP6TVar3TestArray_16X8C

.subckt PadFrame_SP03 PAD0x0 PAD0x1 PAD0x2 PAD0x3 PAD0x4 PAD0x5 PAD0x6 PAD0x7 PAD0x8 PAD0x9 PAD1x0 PAD1x1 PAD1x2 PAD1x3 PAD1x4 PAD1x5 PAD1x6 PAD1x7 PAD1x8 PAD1x9
XPAD0x0 PAD0x0 BondPad
XPAD0x1 PAD0x1 BondPad
XPAD0x2 PAD0x2 BondPad
XPAD0x3 PAD0x3 BondPad
XPAD0x4 PAD0x4 BondPad
XPAD0x5 PAD0x5 BondPad
XPAD0x6 PAD0x6 BondPad
XPAD0x7 PAD0x7 BondPad
XPAD0x8 PAD0x8 BondPad
XPAD0x9 PAD0x9 BondPad
XPAD1x0 PAD1x0 BondPad
XPAD1x1 PAD1x1 BondPad
XPAD1x2 PAD1x2 BondPad
XPAD1x3 PAD1x3 BondPad
XPAD1x4 PAD1x4 BondPad
XPAD1x5 PAD1x5 BondPad
XPAD1x6 PAD1x6 BondPad
XPAD1x7 PAD1x7 BondPad
XPAD1x8 PAD1x8 BondPad
XPAD1x9 PAD1x9 BondPad
.ends PadFrame_SP03

.subckt SP6TVar3 vss noco_vdd noco_wl noco_bl noco_bl_n co_vdd co_bl co_bl_n co_bit co_bit_n co_wl
Xframe noco_vdd noco_wl NoConn_PAD0x2 co_vdd co_bl_n co_bit co_bit_n NoConn_PAD0x7 NoConn_PAD0x8 NoConn_PAD0x9 vss noco_bl noco_bl_n vss co_bl co_wl NoConn_PAD1x6 NoConn_PAD1x7 NoConn_PAD1x8 NoConn_PAD1x9 PadFrame_SP03
Xtestarray_noco vss noco_vdd noco_bl noco_bl_n noco_wl SP6TVar3TestArray_16X8
Xtestarray_co vss co_vdd co_bl co_bl_n co_bit co_bit_n co_wl SP6TVar3TestArray_16X8C
.ends SP6TVar3

.subckt DP8TVar3Cell wl1 wl2 bl1 bl1_n bl2 bl2_n vdd vss
Xpu1 vdd bit_n bit vdd sg13_lv_pmos l=1.3e-07 w=2e-07
Xpd1 bit bit_n vss vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpu2 vdd bit bit_n vdd sg13_lv_pmos l=1.3e-07 w=2e-07
Xpd2 bit_n bit vss vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg1 bit wl1 bl1 vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg1n bit_n wl1 bl1_n vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg2 bit wl2 bl2 vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg2n bit_n wl2 bl2_n vss sg13_lv_nmos l=1.3e-07 w=2e-07
.ends DP8TVar3Cell

.subckt DP8TVar3Array_2X1 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0]
Xinst0x0 wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] vdd vss DP8TVar3Cell
Xinst1x0 wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0] vdd vss DP8TVar3Cell
.ends DP8TVar3Array_2X1

.subckt DP8TVar3Array_2X2 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0] DP8TVar3Array_2X1
Xinst0x1 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TVar3Array_2X1
.ends DP8TVar3Array_2X2

.subckt DP8TVar3Array_4X2 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TVar3Array_2X2
Xinst1x0 vss vdd wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TVar3Array_2X2
.ends DP8TVar3Array_4X2

.subckt DP8TVar3Array_4X4 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TVar3Array_4X2
Xinst0x1 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar3Array_4X2
.ends DP8TVar3Array_4X4

.subckt DP8TVar3Array_8X4 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar3Array_4X4
Xinst1x0 vss vdd wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar3Array_4X4
.ends DP8TVar3Array_8X4

.subckt DP8TVar3Array_8X8 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar3Array_8X4
Xinst0x1 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar3Array_8X4
.ends DP8TVar3Array_8X8

.subckt DP8TVar3BulkConn vdd vss bl1 bl2 bl1_n bl2_n
.ends DP8TVar3BulkConn

.subckt DP8TVar3BulkConnRow_2 vss vdd bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1]
Xinst0 vdd vss bl1[0] bl2[0] bl1_n[0] bl2_n[0] DP8TVar3BulkConn
Xinst1 vdd vss bl1[1] bl2[1] bl1_n[1] bl2_n[1] DP8TVar3BulkConn
.ends DP8TVar3BulkConnRow_2

.subckt DP8TVar3BulkConnRow_4 vss vdd bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3]
Xinst0 vss vdd bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TVar3BulkConnRow_2
Xinst1 vss vdd bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar3BulkConnRow_2
.ends DP8TVar3BulkConnRow_4

.subckt DP8TVar3BulkConnRow_8 vss vdd bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0 vss vdd bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar3BulkConnRow_4
Xinst1 vss vdd bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar3BulkConnRow_4
.ends DP8TVar3BulkConnRow_8

.subckt DP8TVar3Array_16X8BC vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] wl1[8] wl2[8] wl1[9] wl2[9] wl1[10] wl2[10] wl1[11] wl2[11] wl1[12] wl2[12] wl1[13] wl2[13] wl1[14] wl2[14] wl1[15] wl2[15] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar3Array_8X8
Xinst1x0 vss vdd wl1[8] wl2[8] wl1[9] wl2[9] wl1[10] wl2[10] wl1[11] wl2[11] wl1[12] wl2[12] wl1[13] wl2[13] wl1[14] wl2[14] wl1[15] wl2[15] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar3Array_8X8
Xbottombcrow vss vdd bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar3BulkConnRow_8
Xtopbcrow vss vdd bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar3BulkConnRow_8
.ends DP8TVar3Array_16X8BC

.subckt DP8TVar3TestArray_16X8 vss vdd wl1 wl2 bl1 bl1_n bl2 bl2_n
Xarray vss vdd zero zero zero zero zero zero zero zero zero zero zero zero zero zero zero zero wl1 wl2 zero zero zero zero zero zero zero zero zero zero zero zero zero zero bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1 bl1_n bl2 bl2_n bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar3Array_16X8BC
Xzero vdd vss zero zero_x1
.ends DP8TVar3TestArray_16X8

.subckt DP8TVar3Array_4X8 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar3Array_4X4
Xinst0x1 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar3Array_4X4
.ends DP8TVar3Array_4X8

.subckt DP8TVar3Array_2X4 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TVar3Array_2X2
Xinst0x1 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar3Array_2X2
.ends DP8TVar3Array_2X4

.subckt DP8TVar3Array_2X8 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar3Array_2X4
Xinst0x1 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar3Array_2X4
.ends DP8TVar3Array_2X8

.subckt DP8TVar3Array_1X2 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1]
Xinst0x0 wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] vdd vss DP8TVar3Cell
Xinst0x1 wl1[0] wl2[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] vdd vss DP8TVar3Cell
.ends DP8TVar3Array_1X2

.subckt DP8TVar3Array_1X4 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3]
Xinst0x0 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TVar3Array_1X2
Xinst0x1 vss vdd wl1[0] wl2[0] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar3Array_1X2
.ends DP8TVar3Array_1X4

.subckt DP8TVar3Array_1X8 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar3Array_1X4
Xinst0x1 vss vdd wl1[0] wl2[0] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar3Array_1X4
.ends DP8TVar3Array_1X8

.subckt DP8TVar3Array_7X8 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar3Array_4X8
Xinst1x0 vss vdd wl1[4] wl2[4] wl1[5] wl2[5] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar3Array_2X8
Xinst2x0 vss vdd wl1[6] wl2[6] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar3Array_1X8
.ends DP8TVar3Array_7X8

.subckt DP8TVar3CellShWL1 wl1 wl2 bl1 bl1_n bl2 bl2_n vdd vss
Xpu1 vdd bit_n bit vdd sg13_lv_pmos l=1.3e-07 w=2e-07
Xpd1 bit bit_n vss vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpu2 vdd bit bit_n vdd sg13_lv_pmos l=1.3e-07 w=2e-07
Xpd2 bit_n bit vss vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg1 bit wl1 bl1 vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg1n bit_n wl1 bl1_n vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg2 bit wl1 bl2 vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg2n bit_n wl1 bl2_n vss sg13_lv_nmos l=1.3e-07 w=2e-07
.ends DP8TVar3CellShWL1

.subckt DP8TVar3ArrayShWL1_1X2 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1]
Xinst0x0 wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] vdd vss DP8TVar3CellShWL1
Xinst0x1 wl1[0] wl2[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] vdd vss DP8TVar3CellShWL1
.ends DP8TVar3ArrayShWL1_1X2

.subckt DP8TVar3ArrayShWL1_1X4 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3]
Xinst0x0 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TVar3ArrayShWL1_1X2
Xinst0x1 vss vdd wl1[0] wl2[0] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar3ArrayShWL1_1X2
.ends DP8TVar3ArrayShWL1_1X4

.subckt DP8TVar3ArrayShWL1_1X8 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar3ArrayShWL1_1X4
Xinst0x1 vss vdd wl1[0] wl2[0] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar3ArrayShWL1_1X4
.ends DP8TVar3ArrayShWL1_1X8

.subckt DP8TVar3CellConnectOut wl1 wl2 bl1 bl1_n bl2 bl2_n vdd vss bit bit_n
Xpu1 vdd bit_n bit vdd sg13_lv_pmos l=1.3e-07 w=2e-07
Xpd1 bit bit_n vss vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpu2 vdd bit bit_n vdd sg13_lv_pmos l=1.3e-07 w=2e-07
Xpd2 bit_n bit vss vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg1 bit wl1 bl1 vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg1n bit_n wl1 bl1_n vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg2 bit wl2 bl2 vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg2n bit_n wl2 bl2_n vss sg13_lv_nmos l=1.3e-07 w=2e-07
.ends DP8TVar3CellConnectOut

.subckt DP8TVar3CellShWL2 wl1 wl2 bl1 bl1_n bl2 bl2_n vdd vss
Xpu1 vdd bit_n bit vdd sg13_lv_pmos l=1.3e-07 w=2e-07
Xpd1 bit bit_n vss vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpu2 vdd bit bit_n vdd sg13_lv_pmos l=1.3e-07 w=2e-07
Xpd2 bit_n bit vss vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg1 bit wl2 bl1 vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg1n bit_n wl2 bl1_n vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg2 bit wl2 bl2 vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg2n bit_n wl2 bl2_n vss sg13_lv_nmos l=1.3e-07 w=2e-07
.ends DP8TVar3CellShWL2

.subckt DP8TVar3ArrayShWL2_1X2 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1]
Xinst0x0 wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] vdd vss DP8TVar3CellShWL2
Xinst0x1 wl1[0] wl2[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] vdd vss DP8TVar3CellShWL2
.ends DP8TVar3ArrayShWL2_1X2

.subckt DP8TVar3ArrayShWL2_1X4 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3]
Xinst0x0 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TVar3ArrayShWL2_1X2
Xinst0x1 vss vdd wl1[0] wl2[0] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar3ArrayShWL2_1X2
.ends DP8TVar3ArrayShWL2_1X4

.subckt DP8TVar3ArrayShWL2_1X8 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar3ArrayShWL2_1X4
Xinst0x1 vss vdd wl1[0] wl2[0] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar3ArrayShWL2_1X4
.ends DP8TVar3ArrayShWL2_1X8

.subckt DP8TVar3Array_6X8 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar3Array_4X8
Xinst1x0 vss vdd wl1[4] wl2[4] wl1[5] wl2[5] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar3Array_2X8
.ends DP8TVar3Array_6X8

.subckt DP8TVar3TestArray_16X8C vss vdd wl1 wl2 bl1 bl1_n bl2 bl2_n bit bit_n
Xbcconn_bot vss vdd bcconn_bot_bl1[0] bcconn_bot_bl1_n[0] bcconn_bot_bl2[0] bcconn_bot_bl2_n[0] bcconn_bot_bl1[1] bcconn_bot_bl1_n[1] bcconn_bot_bl2[1] bcconn_bot_bl2_n[1] bcconn_bot_bl1[2] bcconn_bot_bl1_n[2] bcconn_bot_bl2[2] bcconn_bot_bl2_n[2] bcconn_bot_bl1[3] bcconn_bot_bl1_n[3] bcconn_bot_bl2[3] bcconn_bot_bl2_n[3] bl1 bl1_n bl2 bl2_n bcconn_bot_bl1[5] bcconn_bot_bl1_n[5] bcconn_bot_bl2[5] bcconn_bot_bl2_n[5] bcconn_bot_bl1[6] bcconn_bot_bl1_n[6] bcconn_bot_bl2[6] bcconn_bot_bl2_n[6] bcconn_bot_bl1[7] bcconn_bot_bl1_n[7] bcconn_bot_bl2[7] bcconn_bot_bl2_n[7] DP8TVar3BulkConnRow_8
Xbcconn_top vss vdd bcconn_top_bl1[0] bcconn_top_bl1_n[0] bcconn_top_bl2[0] bcconn_top_bl2_n[0] bcconn_top_bl1[1] bcconn_top_bl1_n[1] bcconn_top_bl2[1] bcconn_top_bl2_n[1] bcconn_top_bl1[2] bcconn_top_bl1_n[2] bcconn_top_bl2[2] bcconn_top_bl2_n[2] bcconn_top_bl1[3] bcconn_top_bl1_n[3] bcconn_top_bl2[3] bcconn_top_bl2_n[3] bl1 bl1_n bl2 bl2_n bcconn_top_bl1[5] bcconn_top_bl1_n[5] bcconn_top_bl2[5] bcconn_top_bl2_n[5] bcconn_top_bl1[6] bcconn_top_bl1_n[6] bcconn_top_bl2[6] bcconn_top_bl2_n[6] bcconn_top_bl1[7] bcconn_top_bl1_n[7] bcconn_top_bl2[7] bcconn_top_bl2_n[7] DP8TVar3BulkConnRow_8
Xarray_bot vss vdd zero zero zero zero zero zero zero zero zero zero zero zero zero zero array_bot_bl1[0] array_bot_bl1_n[0] array_bot_bl2[0] array_bot_bl2_n[0] array_bot_bl1[1] array_bot_bl1_n[1] array_bot_bl2[1] array_bot_bl2_n[1] array_bot_bl1[2] array_bot_bl1_n[2] array_bot_bl2[2] array_bot_bl2_n[2] array_bot_bl1[3] array_bot_bl1_n[3] array_bot_bl2[3] array_bot_bl2_n[3] bl1 bl1_n bl2 bl2_n array_bot_bl1[5] array_bot_bl1_n[5] array_bot_bl2[5] array_bot_bl2_n[5] array_bot_bl1[6] array_bot_bl1_n[6] array_bot_bl2[6] array_bot_bl2_n[6] array_bot_bl1[7] array_bot_bl1_n[7] array_bot_bl2[7] array_bot_bl2_n[7] DP8TVar3Array_7X8
Xshwl1_row vss vdd zero bit shwl1_row_bl1[0] shwl1_row_bl1_n[0] shwl1_row_bl2[0] shwl1_row_bl2_n[0] shwl1_row_bl1[1] shwl1_row_bl1_n[1] shwl1_row_bl2[1] shwl1_row_bl2_n[1] shwl1_row_bl1[2] shwl1_row_bl1_n[2] shwl1_row_bl2[2] shwl1_row_bl2_n[2] shwl1_row_bl1[3] shwl1_row_bl1_n[3] shwl1_row_bl2[3] shwl1_row_bl2_n[3] bl1 bl1_n bl2 bl2_n shwl1_row_bl1[5] shwl1_row_bl1_n[5] shwl1_row_bl2[5] shwl1_row_bl2_n[5] shwl1_row_bl1[6] shwl1_row_bl1_n[6] shwl1_row_bl2[6] shwl1_row_bl2_n[6] shwl1_row_bl1[7] shwl1_row_bl1_n[7] shwl1_row_bl2[7] shwl1_row_bl2_n[7] DP8TVar3ArrayShWL1_1X8
Xcell_cols_left vss vdd wl1 wl2 cell_cols_left_bl1[0] cell_cols_left_bl1_n[0] cell_cols_left_bl2[0] cell_cols_left_bl2_n[0] cell_cols_left_bl1[1] cell_cols_left_bl1_n[1] cell_cols_left_bl2[1] cell_cols_left_bl2_n[1] cell_cols_left_bl1[2] cell_cols_left_bl1_n[2] cell_cols_left_bl2[2] cell_cols_left_bl2_n[2] cell_cols_left_bl1[3] cell_cols_left_bl1_n[3] cell_cols_left_bl2[3] cell_cols_left_bl2_n[3] DP8TVar3Array_1X4
Xconncell wl1 wl2 bl1 bl1_n bl2 bl2_n vdd vss bit bit_n DP8TVar3CellConnectOut
Xfillcell wl1 wl2 fillcell_bl1 fillcell_bl1_n fillcell_bl2 fillcell_bl2_n vdd vss DP8TVar3Cell
Xcell_cols_right vss vdd wl1 wl2 cell_cols_right_bl1[0] cell_cols_right_bl1_n[0] cell_cols_right_bl2[0] cell_cols_right_bl2_n[0] cell_cols_right_bl1[1] cell_cols_right_bl1_n[1] cell_cols_right_bl2[1] cell_cols_right_bl2_n[1] DP8TVar3Array_1X2
Xshwl2_row vss vdd bit_n zero shwl2_row_bl1[0] shwl2_row_bl1_n[0] shwl2_row_bl2[0] shwl2_row_bl2_n[0] shwl2_row_bl1[1] shwl2_row_bl1_n[1] shwl2_row_bl2[1] shwl2_row_bl2_n[1] shwl2_row_bl1[2] shwl2_row_bl1_n[2] shwl2_row_bl2[2] shwl2_row_bl2_n[2] shwl2_row_bl1[3] shwl2_row_bl1_n[3] shwl2_row_bl2[3] shwl2_row_bl2_n[3] bl1 bl1_n bl2 bl2_n shwl2_row_bl1[5] shwl2_row_bl1_n[5] shwl2_row_bl2[5] shwl2_row_bl2_n[5] shwl2_row_bl1[6] shwl2_row_bl1_n[6] shwl2_row_bl2[6] shwl2_row_bl2_n[6] shwl2_row_bl1[7] shwl2_row_bl1_n[7] shwl2_row_bl2[7] shwl2_row_bl2_n[7] DP8TVar3ArrayShWL2_1X8
Xarray_top vss vdd zero zero zero zero zero zero zero zero zero zero zero zero array_top_bl1[0] array_top_bl1_n[0] array_top_bl2[0] array_top_bl2_n[0] array_top_bl1[1] array_top_bl1_n[1] array_top_bl2[1] array_top_bl2_n[1] array_top_bl1[2] array_top_bl1_n[2] array_top_bl2[2] array_top_bl2_n[2] array_top_bl1[3] array_top_bl1_n[3] array_top_bl2[3] array_top_bl2_n[3] bl1 bl1_n bl2 bl2_n array_top_bl1[5] array_top_bl1_n[5] array_top_bl2[5] array_top_bl2_n[5] array_top_bl1[6] array_top_bl1_n[6] array_top_bl2[6] array_top_bl2_n[6] array_top_bl1[7] array_top_bl1_n[7] array_top_bl2[7] array_top_bl2_n[7] DP8TVar3Array_6X8
Xzero vdd vss zero zero_x1
.ends DP8TVar3TestArray_16X8C

.subckt PadFrame_DP03 PAD0x0 PAD0x1 PAD0x2 PAD0x3 PAD0x4 PAD0x5 PAD0x6 PAD0x7 PAD0x8 PAD0x9 PAD1x0 PAD1x1 PAD1x2 PAD1x3 PAD1x4 PAD1x5 PAD1x6 PAD1x7 PAD1x8 PAD1x9
XPAD0x0 PAD0x0 BondPad
XPAD0x1 PAD0x1 BondPad
XPAD0x2 PAD0x2 BondPad
XPAD0x3 PAD0x3 BondPad
XPAD0x4 PAD0x4 BondPad
XPAD0x5 PAD0x5 BondPad
XPAD0x6 PAD0x6 BondPad
XPAD0x7 PAD0x7 BondPad
XPAD0x8 PAD0x8 BondPad
XPAD0x9 PAD0x9 BondPad
XPAD1x0 PAD1x0 BondPad
XPAD1x1 PAD1x1 BondPad
XPAD1x2 PAD1x2 BondPad
XPAD1x3 PAD1x3 BondPad
XPAD1x4 PAD1x4 BondPad
XPAD1x5 PAD1x5 BondPad
XPAD1x6 PAD1x6 BondPad
XPAD1x7 PAD1x7 BondPad
XPAD1x8 PAD1x8 BondPad
XPAD1x9 PAD1x9 BondPad
.ends PadFrame_DP03

.subckt DP8TVar3 vss noco_vdd noco_wl1 noco_wl2 noco_bl1 noco_bl1_n noco_bl2 noco_bl2_n co_vdd co_bit co_bit_n co_wl1 co_wl2 co_bl1 co_bl1_n co_bl2_n co_bl2
Xframe noco_vdd noco_wl1 noco_wl2 noco_bl2 co_vdd co_bit co_bit_n co_wl1 co_wl2 NoConn_PAD0x9 vss noco_bl1 noco_bl1_n noco_bl2_n vss co_bl1 co_bl1_n co_bl2_n co_bl2 NoConn_PAD1x9 PadFrame_DP03
Xtestarray_noco vss noco_vdd noco_wl1 noco_wl2 noco_bl1 noco_bl1_n noco_bl2 noco_bl2_n DP8TVar3TestArray_16X8
Xtestarray_co vss co_vdd co_wl1 co_wl2 co_bl1 co_bl1_n co_bl2 co_bl2_n co_bit co_bit_n DP8TVar3TestArray_16X8C
.ends DP8TVar3

.subckt SP6TVar4Cell wl bl bl_n vdd vss
Xpu1 vdd bit_n bit vdd sg13_lv_pmos l=1.3e-07 w=1.5e-07
Xpd1 bit bit_n vss vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpu2 vdd bit bit_n vdd sg13_lv_pmos l=1.3e-07 w=1.5e-07
Xpd2 bit_n bit vss vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg1 bit wl bl vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg2 bit_n wl bl_n vss sg13_lv_nmos l=1.3e-07 w=2e-07
.ends SP6TVar4Cell

.subckt SP6TVar4Array_2X1 vss vdd wl[0] wl[1] bl[0] bl_n[0]
Xinst0x0 wl[0] bl[0] bl_n[0] vdd vss SP6TVar4Cell
Xinst1x0 wl[1] bl[0] bl_n[0] vdd vss SP6TVar4Cell
.ends SP6TVar4Array_2X1

.subckt SP6TVar4Array_2X2 vss vdd wl[0] wl[1] bl[0] bl_n[0] bl[1] bl_n[1]
Xinst0x0 vss vdd wl[0] wl[1] bl[0] bl_n[0] SP6TVar4Array_2X1
Xinst0x1 vss vdd wl[0] wl[1] bl[1] bl_n[1] SP6TVar4Array_2X1
.ends SP6TVar4Array_2X2

.subckt SP6TVar4Array_4X2 vss vdd wl[0] wl[1] wl[2] wl[3] bl[0] bl_n[0] bl[1] bl_n[1]
Xinst0x0 vss vdd wl[0] wl[1] bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar4Array_2X2
Xinst1x0 vss vdd wl[2] wl[3] bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar4Array_2X2
.ends SP6TVar4Array_4X2

.subckt SP6TVar4Array_4X4 vss vdd wl[0] wl[1] wl[2] wl[3] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar4Array_4X2
Xinst0x1 vss vdd wl[0] wl[1] wl[2] wl[3] bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar4Array_4X2
.ends SP6TVar4Array_4X4

.subckt SP6TVar4Array_8X4 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar4Array_4X4
Xinst1x0 vss vdd wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar4Array_4X4
.ends SP6TVar4Array_8X4

.subckt SP6TVar4Array_8X8 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar4Array_8X4
Xinst0x1 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7] SP6TVar4Array_8X4
.ends SP6TVar4Array_8X8

.subckt SP6TVar4BulkConn vdd vss bl bl_n
.ends SP6TVar4BulkConn

.subckt SP6TVar4BulkConnRow_2 vss vdd bl[0] bl_n[0] bl[1] bl_n[1]
Xinst0 vdd vss bl[0] bl_n[0] SP6TVar4BulkConn
Xinst1 vdd vss bl[1] bl_n[1] SP6TVar4BulkConn
.ends SP6TVar4BulkConnRow_2

.subckt SP6TVar4BulkConnRow_4 vss vdd bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3]
Xinst0 vss vdd bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar4BulkConnRow_2
Xinst1 vss vdd bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar4BulkConnRow_2
.ends SP6TVar4BulkConnRow_4

.subckt SP6TVar4BulkConnRow_8 vss vdd bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7]
Xinst0 vss vdd bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar4BulkConnRow_4
Xinst1 vss vdd bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7] SP6TVar4BulkConnRow_4
.ends SP6TVar4BulkConnRow_8

.subckt SP6TVar4Array_16X8BC vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7] SP6TVar4Array_8X8
Xinst1x0 vss vdd wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7] SP6TVar4Array_8X8
Xbottombcrow vss vdd bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7] SP6TVar4BulkConnRow_8
Xtopbcrow vss vdd bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7] SP6TVar4BulkConnRow_8
.ends SP6TVar4Array_16X8BC

.subckt SP6TVar4TestArray_16X8 vss vdd bl bl_n wl
Xarray vss vdd zero zero zero zero zero zero zero zero wl zero zero zero zero zero zero zero bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl bl_n bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7] SP6TVar4Array_16X8BC
Xzero vdd vss zero zero_x1
.ends SP6TVar4TestArray_16X8

.subckt SP6TVar4Array_4X1 vss vdd wl[0] wl[1] wl[2] wl[3] bl[0] bl_n[0]
Xinst0x0 vss vdd wl[0] wl[1] bl[0] bl_n[0] SP6TVar4Array_2X1
Xinst1x0 vss vdd wl[2] wl[3] bl[0] bl_n[0] SP6TVar4Array_2X1
.ends SP6TVar4Array_4X1

.subckt SP6TVar4Array_8X1 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] bl[0] bl_n[0] SP6TVar4Array_4X1
Xinst1x0 vss vdd wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] SP6TVar4Array_4X1
.ends SP6TVar4Array_8X1

.subckt SP6TVar4Array_16X1BC vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] bl[0] bl_n[0]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] SP6TVar4Array_8X1
Xinst1x0 vss vdd wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] bl[0] bl_n[0] SP6TVar4Array_8X1
Xbottombcrow vdd vss bl[0] bl_n[0] SP6TVar4BulkConn
Xtopbcrow vdd vss bl[0] bl_n[0] SP6TVar4BulkConn
.ends SP6TVar4Array_16X1BC

.subckt SP6TVar4Array_8X2 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar4Array_4X2
Xinst1x0 vss vdd wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar4Array_4X2
.ends SP6TVar4Array_8X2

.subckt SP6TVar4Array_16X2BC vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] bl[0] bl_n[0] bl[1] bl_n[1]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar4Array_8X2
Xinst1x0 vss vdd wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar4Array_8X2
Xbottombcrow vss vdd bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar4BulkConnRow_2
Xtopbcrow vss vdd bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar4BulkConnRow_2
.ends SP6TVar4Array_16X2BC

.subckt SP6TVar4Array_16X4BC vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar4Array_8X4
Xinst1x0 vss vdd wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar4Array_8X4
Xbottombcrow vss vdd bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar4BulkConnRow_4
Xtopbcrow vss vdd bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar4BulkConnRow_4
.ends SP6TVar4Array_16X4BC

.subckt SP6TVar4Array_6X1 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] bl[0] bl_n[0]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] bl[0] bl_n[0] SP6TVar4Array_4X1
Xinst1x0 vss vdd wl[4] wl[5] bl[0] bl_n[0] SP6TVar4Array_2X1
.ends SP6TVar4Array_6X1

.subckt SP6TVar4CellConnectOut wl bl bl_n vdd vss bit bit_n
Xpu1 vdd bit_n bit vdd sg13_lv_pmos l=1.3e-07 w=1.5e-07
Xpd1 bit bit_n vss vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpu2 vdd bit bit_n vdd sg13_lv_pmos l=1.3e-07 w=1.5e-07
Xpd2 bit_n bit vss vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg1 bit wl bl vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg2 bit_n wl bl_n vss sg13_lv_nmos l=1.3e-07 w=2e-07
.ends SP6TVar4CellConnectOut

.subckt SP6TVar4TestArray_16X8C vss vdd bl bl_n bit bit_n wl
Xarray_0 vss vdd zero zero zero zero zero zero zero zero wl zero zero zero zero zero zero zero array_0_bl[0] array_0_bl_n[0] SP6TVar4Array_16X1BC
Xarray_1 vss vdd zero zero zero zero zero zero zero zero wl zero zero zero zero zero zero zero array_1_bl[0] array_1_bl_n[0] array_1_bl[1] array_1_bl_n[1] SP6TVar4Array_16X2BC
Xarray_2 vss vdd zero zero zero zero zero zero zero zero wl zero zero zero zero zero zero zero array_2_bl[0] array_2_bl_n[0] array_2_bl[1] array_2_bl_n[1] array_2_bl[2] array_2_bl_n[2] array_2_bl[3] array_2_bl_n[3] SP6TVar4Array_16X4BC
Xcolbc_0 vdd vss bl bl_n SP6TVar4BulkConn
Xcolbc_1 vdd vss bl bl_n SP6TVar4BulkConn
Xcolarray_0 vss vdd zero zero zero zero zero zero zero zero bl bl_n SP6TVar4Array_8X1
Xcolarray_1 vss vdd zero zero zero zero zero zero bl bl_n SP6TVar4Array_6X1
Xbc_noconn zero bl bl_n vdd vss SP6TVar4Cell
Xbc_conn wl bl bl_n vdd vss bit bit_n SP6TVar4CellConnectOut
Xzero vdd vss zero zero_x1
.ends SP6TVar4TestArray_16X8C

.subckt PadFrame_SP04 PAD0x0 PAD0x1 PAD0x2 PAD0x3 PAD0x4 PAD0x5 PAD0x6 PAD0x7 PAD0x8 PAD0x9 PAD1x0 PAD1x1 PAD1x2 PAD1x3 PAD1x4 PAD1x5 PAD1x6 PAD1x7 PAD1x8 PAD1x9
XPAD0x0 PAD0x0 BondPad
XPAD0x1 PAD0x1 BondPad
XPAD0x2 PAD0x2 BondPad
XPAD0x3 PAD0x3 BondPad
XPAD0x4 PAD0x4 BondPad
XPAD0x5 PAD0x5 BondPad
XPAD0x6 PAD0x6 BondPad
XPAD0x7 PAD0x7 BondPad
XPAD0x8 PAD0x8 BondPad
XPAD0x9 PAD0x9 BondPad
XPAD1x0 PAD1x0 BondPad
XPAD1x1 PAD1x1 BondPad
XPAD1x2 PAD1x2 BondPad
XPAD1x3 PAD1x3 BondPad
XPAD1x4 PAD1x4 BondPad
XPAD1x5 PAD1x5 BondPad
XPAD1x6 PAD1x6 BondPad
XPAD1x7 PAD1x7 BondPad
XPAD1x8 PAD1x8 BondPad
XPAD1x9 PAD1x9 BondPad
.ends PadFrame_SP04

.subckt SP6TVar4 vss noco_vdd noco_wl noco_bl noco_bl_n co_vdd co_bl co_bl_n co_bit co_bit_n co_wl
Xframe noco_vdd noco_wl NoConn_PAD0x2 co_vdd co_bl_n co_bit co_bit_n NoConn_PAD0x7 NoConn_PAD0x8 NoConn_PAD0x9 vss noco_bl noco_bl_n vss co_bl co_wl NoConn_PAD1x6 NoConn_PAD1x7 NoConn_PAD1x8 NoConn_PAD1x9 PadFrame_SP04
Xtestarray_noco vss noco_vdd noco_bl noco_bl_n noco_wl SP6TVar4TestArray_16X8
Xtestarray_co vss co_vdd co_bl co_bl_n co_bit co_bit_n co_wl SP6TVar4TestArray_16X8C
.ends SP6TVar4

.subckt DP8TVar4Cell wl1 wl2 bl1 bl1_n bl2 bl2_n vdd vss
Xpu1 vdd bit_n bit vdd sg13_lv_pmos l=1.3e-07 w=1.5e-07
Xpd1 bit bit_n vss vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpu2 vdd bit bit_n vdd sg13_lv_pmos l=1.3e-07 w=1.5e-07
Xpd2 bit_n bit vss vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg1 bit wl1 bl1 vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg1n bit_n wl1 bl1_n vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg2 bit wl2 bl2 vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg2n bit_n wl2 bl2_n vss sg13_lv_nmos l=1.3e-07 w=2e-07
.ends DP8TVar4Cell

.subckt DP8TVar4Array_2X1 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0]
Xinst0x0 wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] vdd vss DP8TVar4Cell
Xinst1x0 wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0] vdd vss DP8TVar4Cell
.ends DP8TVar4Array_2X1

.subckt DP8TVar4Array_2X2 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0] DP8TVar4Array_2X1
Xinst0x1 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TVar4Array_2X1
.ends DP8TVar4Array_2X2

.subckt DP8TVar4Array_4X2 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TVar4Array_2X2
Xinst1x0 vss vdd wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TVar4Array_2X2
.ends DP8TVar4Array_4X2

.subckt DP8TVar4Array_4X4 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TVar4Array_4X2
Xinst0x1 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar4Array_4X2
.ends DP8TVar4Array_4X4

.subckt DP8TVar4Array_8X4 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar4Array_4X4
Xinst1x0 vss vdd wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar4Array_4X4
.ends DP8TVar4Array_8X4

.subckt DP8TVar4Array_8X8 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar4Array_8X4
Xinst0x1 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar4Array_8X4
.ends DP8TVar4Array_8X8

.subckt DP8TVar4BulkConn vdd vss bl1 bl2 bl1_n bl2_n
.ends DP8TVar4BulkConn

.subckt DP8TVar4BulkConnRow_2 vss vdd bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1]
Xinst0 vdd vss bl1[0] bl2[0] bl1_n[0] bl2_n[0] DP8TVar4BulkConn
Xinst1 vdd vss bl1[1] bl2[1] bl1_n[1] bl2_n[1] DP8TVar4BulkConn
.ends DP8TVar4BulkConnRow_2

.subckt DP8TVar4BulkConnRow_4 vss vdd bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3]
Xinst0 vss vdd bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TVar4BulkConnRow_2
Xinst1 vss vdd bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar4BulkConnRow_2
.ends DP8TVar4BulkConnRow_4

.subckt DP8TVar4BulkConnRow_8 vss vdd bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0 vss vdd bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar4BulkConnRow_4
Xinst1 vss vdd bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar4BulkConnRow_4
.ends DP8TVar4BulkConnRow_8

.subckt DP8TVar4Array_16X8BC vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] wl1[8] wl2[8] wl1[9] wl2[9] wl1[10] wl2[10] wl1[11] wl2[11] wl1[12] wl2[12] wl1[13] wl2[13] wl1[14] wl2[14] wl1[15] wl2[15] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar4Array_8X8
Xinst1x0 vss vdd wl1[8] wl2[8] wl1[9] wl2[9] wl1[10] wl2[10] wl1[11] wl2[11] wl1[12] wl2[12] wl1[13] wl2[13] wl1[14] wl2[14] wl1[15] wl2[15] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar4Array_8X8
Xbottombcrow vss vdd bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar4BulkConnRow_8
Xtopbcrow vss vdd bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar4BulkConnRow_8
.ends DP8TVar4Array_16X8BC

.subckt DP8TVar4TestArray_16X8 vss vdd wl1 wl2 bl1 bl1_n bl2 bl2_n
Xarray vss vdd zero zero zero zero zero zero zero zero zero zero zero zero zero zero zero zero wl1 wl2 zero zero zero zero zero zero zero zero zero zero zero zero zero zero bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1 bl1_n bl2 bl2_n bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar4Array_16X8BC
Xzero vdd vss zero zero_x1
.ends DP8TVar4TestArray_16X8

.subckt DP8TVar4Array_4X8 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar4Array_4X4
Xinst0x1 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar4Array_4X4
.ends DP8TVar4Array_4X8

.subckt DP8TVar4Array_2X4 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TVar4Array_2X2
Xinst0x1 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar4Array_2X2
.ends DP8TVar4Array_2X4

.subckt DP8TVar4Array_2X8 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar4Array_2X4
Xinst0x1 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar4Array_2X4
.ends DP8TVar4Array_2X8

.subckt DP8TVar4Array_1X2 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1]
Xinst0x0 wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] vdd vss DP8TVar4Cell
Xinst0x1 wl1[0] wl2[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] vdd vss DP8TVar4Cell
.ends DP8TVar4Array_1X2

.subckt DP8TVar4Array_1X4 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3]
Xinst0x0 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TVar4Array_1X2
Xinst0x1 vss vdd wl1[0] wl2[0] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar4Array_1X2
.ends DP8TVar4Array_1X4

.subckt DP8TVar4Array_1X8 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar4Array_1X4
Xinst0x1 vss vdd wl1[0] wl2[0] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar4Array_1X4
.ends DP8TVar4Array_1X8

.subckt DP8TVar4Array_7X8 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar4Array_4X8
Xinst1x0 vss vdd wl1[4] wl2[4] wl1[5] wl2[5] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar4Array_2X8
Xinst2x0 vss vdd wl1[6] wl2[6] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar4Array_1X8
.ends DP8TVar4Array_7X8

.subckt DP8TVar4CellShWL1 wl1 wl2 bl1 bl1_n bl2 bl2_n vdd vss
Xpu1 vdd bit_n bit vdd sg13_lv_pmos l=1.3e-07 w=1.5e-07
Xpd1 bit bit_n vss vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpu2 vdd bit bit_n vdd sg13_lv_pmos l=1.3e-07 w=1.5e-07
Xpd2 bit_n bit vss vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg1 bit wl1 bl1 vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg1n bit_n wl1 bl1_n vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg2 bit wl1 bl2 vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg2n bit_n wl1 bl2_n vss sg13_lv_nmos l=1.3e-07 w=2e-07
.ends DP8TVar4CellShWL1

.subckt DP8TVar4ArrayShWL1_1X2 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1]
Xinst0x0 wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] vdd vss DP8TVar4CellShWL1
Xinst0x1 wl1[0] wl2[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] vdd vss DP8TVar4CellShWL1
.ends DP8TVar4ArrayShWL1_1X2

.subckt DP8TVar4ArrayShWL1_1X4 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3]
Xinst0x0 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TVar4ArrayShWL1_1X2
Xinst0x1 vss vdd wl1[0] wl2[0] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar4ArrayShWL1_1X2
.ends DP8TVar4ArrayShWL1_1X4

.subckt DP8TVar4ArrayShWL1_1X8 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar4ArrayShWL1_1X4
Xinst0x1 vss vdd wl1[0] wl2[0] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar4ArrayShWL1_1X4
.ends DP8TVar4ArrayShWL1_1X8

.subckt DP8TVar4CellConnectOut wl1 wl2 bl1 bl1_n bl2 bl2_n vdd vss bit bit_n
Xpu1 vdd bit_n bit vdd sg13_lv_pmos l=1.3e-07 w=1.5e-07
Xpd1 bit bit_n vss vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpu2 vdd bit bit_n vdd sg13_lv_pmos l=1.3e-07 w=1.5e-07
Xpd2 bit_n bit vss vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg1 bit wl1 bl1 vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg1n bit_n wl1 bl1_n vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg2 bit wl2 bl2 vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg2n bit_n wl2 bl2_n vss sg13_lv_nmos l=1.3e-07 w=2e-07
.ends DP8TVar4CellConnectOut

.subckt DP8TVar4CellShWL2 wl1 wl2 bl1 bl1_n bl2 bl2_n vdd vss
Xpu1 vdd bit_n bit vdd sg13_lv_pmos l=1.3e-07 w=1.5e-07
Xpd1 bit bit_n vss vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpu2 vdd bit bit_n vdd sg13_lv_pmos l=1.3e-07 w=1.5e-07
Xpd2 bit_n bit vss vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg1 bit wl2 bl1 vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg1n bit_n wl2 bl1_n vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg2 bit wl2 bl2 vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg2n bit_n wl2 bl2_n vss sg13_lv_nmos l=1.3e-07 w=2e-07
.ends DP8TVar4CellShWL2

.subckt DP8TVar4ArrayShWL2_1X2 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1]
Xinst0x0 wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] vdd vss DP8TVar4CellShWL2
Xinst0x1 wl1[0] wl2[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] vdd vss DP8TVar4CellShWL2
.ends DP8TVar4ArrayShWL2_1X2

.subckt DP8TVar4ArrayShWL2_1X4 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3]
Xinst0x0 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TVar4ArrayShWL2_1X2
Xinst0x1 vss vdd wl1[0] wl2[0] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar4ArrayShWL2_1X2
.ends DP8TVar4ArrayShWL2_1X4

.subckt DP8TVar4ArrayShWL2_1X8 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar4ArrayShWL2_1X4
Xinst0x1 vss vdd wl1[0] wl2[0] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar4ArrayShWL2_1X4
.ends DP8TVar4ArrayShWL2_1X8

.subckt DP8TVar4Array_6X8 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar4Array_4X8
Xinst1x0 vss vdd wl1[4] wl2[4] wl1[5] wl2[5] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar4Array_2X8
.ends DP8TVar4Array_6X8

.subckt DP8TVar4TestArray_16X8C vss vdd wl1 wl2 bl1 bl1_n bl2 bl2_n bit bit_n
Xbcconn_bot vss vdd bcconn_bot_bl1[0] bcconn_bot_bl1_n[0] bcconn_bot_bl2[0] bcconn_bot_bl2_n[0] bcconn_bot_bl1[1] bcconn_bot_bl1_n[1] bcconn_bot_bl2[1] bcconn_bot_bl2_n[1] bcconn_bot_bl1[2] bcconn_bot_bl1_n[2] bcconn_bot_bl2[2] bcconn_bot_bl2_n[2] bcconn_bot_bl1[3] bcconn_bot_bl1_n[3] bcconn_bot_bl2[3] bcconn_bot_bl2_n[3] bl1 bl1_n bl2 bl2_n bcconn_bot_bl1[5] bcconn_bot_bl1_n[5] bcconn_bot_bl2[5] bcconn_bot_bl2_n[5] bcconn_bot_bl1[6] bcconn_bot_bl1_n[6] bcconn_bot_bl2[6] bcconn_bot_bl2_n[6] bcconn_bot_bl1[7] bcconn_bot_bl1_n[7] bcconn_bot_bl2[7] bcconn_bot_bl2_n[7] DP8TVar4BulkConnRow_8
Xbcconn_top vss vdd bcconn_top_bl1[0] bcconn_top_bl1_n[0] bcconn_top_bl2[0] bcconn_top_bl2_n[0] bcconn_top_bl1[1] bcconn_top_bl1_n[1] bcconn_top_bl2[1] bcconn_top_bl2_n[1] bcconn_top_bl1[2] bcconn_top_bl1_n[2] bcconn_top_bl2[2] bcconn_top_bl2_n[2] bcconn_top_bl1[3] bcconn_top_bl1_n[3] bcconn_top_bl2[3] bcconn_top_bl2_n[3] bl1 bl1_n bl2 bl2_n bcconn_top_bl1[5] bcconn_top_bl1_n[5] bcconn_top_bl2[5] bcconn_top_bl2_n[5] bcconn_top_bl1[6] bcconn_top_bl1_n[6] bcconn_top_bl2[6] bcconn_top_bl2_n[6] bcconn_top_bl1[7] bcconn_top_bl1_n[7] bcconn_top_bl2[7] bcconn_top_bl2_n[7] DP8TVar4BulkConnRow_8
Xarray_bot vss vdd zero zero zero zero zero zero zero zero zero zero zero zero zero zero array_bot_bl1[0] array_bot_bl1_n[0] array_bot_bl2[0] array_bot_bl2_n[0] array_bot_bl1[1] array_bot_bl1_n[1] array_bot_bl2[1] array_bot_bl2_n[1] array_bot_bl1[2] array_bot_bl1_n[2] array_bot_bl2[2] array_bot_bl2_n[2] array_bot_bl1[3] array_bot_bl1_n[3] array_bot_bl2[3] array_bot_bl2_n[3] bl1 bl1_n bl2 bl2_n array_bot_bl1[5] array_bot_bl1_n[5] array_bot_bl2[5] array_bot_bl2_n[5] array_bot_bl1[6] array_bot_bl1_n[6] array_bot_bl2[6] array_bot_bl2_n[6] array_bot_bl1[7] array_bot_bl1_n[7] array_bot_bl2[7] array_bot_bl2_n[7] DP8TVar4Array_7X8
Xshwl1_row vss vdd zero bit shwl1_row_bl1[0] shwl1_row_bl1_n[0] shwl1_row_bl2[0] shwl1_row_bl2_n[0] shwl1_row_bl1[1] shwl1_row_bl1_n[1] shwl1_row_bl2[1] shwl1_row_bl2_n[1] shwl1_row_bl1[2] shwl1_row_bl1_n[2] shwl1_row_bl2[2] shwl1_row_bl2_n[2] shwl1_row_bl1[3] shwl1_row_bl1_n[3] shwl1_row_bl2[3] shwl1_row_bl2_n[3] bl1 bl1_n bl2 bl2_n shwl1_row_bl1[5] shwl1_row_bl1_n[5] shwl1_row_bl2[5] shwl1_row_bl2_n[5] shwl1_row_bl1[6] shwl1_row_bl1_n[6] shwl1_row_bl2[6] shwl1_row_bl2_n[6] shwl1_row_bl1[7] shwl1_row_bl1_n[7] shwl1_row_bl2[7] shwl1_row_bl2_n[7] DP8TVar4ArrayShWL1_1X8
Xcell_cols_left vss vdd wl1 wl2 cell_cols_left_bl1[0] cell_cols_left_bl1_n[0] cell_cols_left_bl2[0] cell_cols_left_bl2_n[0] cell_cols_left_bl1[1] cell_cols_left_bl1_n[1] cell_cols_left_bl2[1] cell_cols_left_bl2_n[1] cell_cols_left_bl1[2] cell_cols_left_bl1_n[2] cell_cols_left_bl2[2] cell_cols_left_bl2_n[2] cell_cols_left_bl1[3] cell_cols_left_bl1_n[3] cell_cols_left_bl2[3] cell_cols_left_bl2_n[3] DP8TVar4Array_1X4
Xconncell wl1 wl2 bl1 bl1_n bl2 bl2_n vdd vss bit bit_n DP8TVar4CellConnectOut
Xfillcell wl1 wl2 fillcell_bl1 fillcell_bl1_n fillcell_bl2 fillcell_bl2_n vdd vss DP8TVar4Cell
Xcell_cols_right vss vdd wl1 wl2 cell_cols_right_bl1[0] cell_cols_right_bl1_n[0] cell_cols_right_bl2[0] cell_cols_right_bl2_n[0] cell_cols_right_bl1[1] cell_cols_right_bl1_n[1] cell_cols_right_bl2[1] cell_cols_right_bl2_n[1] DP8TVar4Array_1X2
Xshwl2_row vss vdd bit_n zero shwl2_row_bl1[0] shwl2_row_bl1_n[0] shwl2_row_bl2[0] shwl2_row_bl2_n[0] shwl2_row_bl1[1] shwl2_row_bl1_n[1] shwl2_row_bl2[1] shwl2_row_bl2_n[1] shwl2_row_bl1[2] shwl2_row_bl1_n[2] shwl2_row_bl2[2] shwl2_row_bl2_n[2] shwl2_row_bl1[3] shwl2_row_bl1_n[3] shwl2_row_bl2[3] shwl2_row_bl2_n[3] bl1 bl1_n bl2 bl2_n shwl2_row_bl1[5] shwl2_row_bl1_n[5] shwl2_row_bl2[5] shwl2_row_bl2_n[5] shwl2_row_bl1[6] shwl2_row_bl1_n[6] shwl2_row_bl2[6] shwl2_row_bl2_n[6] shwl2_row_bl1[7] shwl2_row_bl1_n[7] shwl2_row_bl2[7] shwl2_row_bl2_n[7] DP8TVar4ArrayShWL2_1X8
Xarray_top vss vdd zero zero zero zero zero zero zero zero zero zero zero zero array_top_bl1[0] array_top_bl1_n[0] array_top_bl2[0] array_top_bl2_n[0] array_top_bl1[1] array_top_bl1_n[1] array_top_bl2[1] array_top_bl2_n[1] array_top_bl1[2] array_top_bl1_n[2] array_top_bl2[2] array_top_bl2_n[2] array_top_bl1[3] array_top_bl1_n[3] array_top_bl2[3] array_top_bl2_n[3] bl1 bl1_n bl2 bl2_n array_top_bl1[5] array_top_bl1_n[5] array_top_bl2[5] array_top_bl2_n[5] array_top_bl1[6] array_top_bl1_n[6] array_top_bl2[6] array_top_bl2_n[6] array_top_bl1[7] array_top_bl1_n[7] array_top_bl2[7] array_top_bl2_n[7] DP8TVar4Array_6X8
Xzero vdd vss zero zero_x1
.ends DP8TVar4TestArray_16X8C

.subckt PadFrame_DP04 PAD0x0 PAD0x1 PAD0x2 PAD0x3 PAD0x4 PAD0x5 PAD0x6 PAD0x7 PAD0x8 PAD0x9 PAD1x0 PAD1x1 PAD1x2 PAD1x3 PAD1x4 PAD1x5 PAD1x6 PAD1x7 PAD1x8 PAD1x9
XPAD0x0 PAD0x0 BondPad
XPAD0x1 PAD0x1 BondPad
XPAD0x2 PAD0x2 BondPad
XPAD0x3 PAD0x3 BondPad
XPAD0x4 PAD0x4 BondPad
XPAD0x5 PAD0x5 BondPad
XPAD0x6 PAD0x6 BondPad
XPAD0x7 PAD0x7 BondPad
XPAD0x8 PAD0x8 BondPad
XPAD0x9 PAD0x9 BondPad
XPAD1x0 PAD1x0 BondPad
XPAD1x1 PAD1x1 BondPad
XPAD1x2 PAD1x2 BondPad
XPAD1x3 PAD1x3 BondPad
XPAD1x4 PAD1x4 BondPad
XPAD1x5 PAD1x5 BondPad
XPAD1x6 PAD1x6 BondPad
XPAD1x7 PAD1x7 BondPad
XPAD1x8 PAD1x8 BondPad
XPAD1x9 PAD1x9 BondPad
.ends PadFrame_DP04

.subckt DP8TVar4 vss noco_vdd noco_wl1 noco_wl2 noco_bl1 noco_bl1_n noco_bl2 noco_bl2_n co_vdd co_bit co_bit_n co_wl1 co_wl2 co_bl1 co_bl1_n co_bl2_n co_bl2
Xframe noco_vdd noco_wl1 noco_wl2 noco_bl2 co_vdd co_bit co_bit_n co_wl1 co_wl2 NoConn_PAD0x9 vss noco_bl1 noco_bl1_n noco_bl2_n vss co_bl1 co_bl1_n co_bl2_n co_bl2 NoConn_PAD1x9 PadFrame_DP04
Xtestarray_noco vss noco_vdd noco_wl1 noco_wl2 noco_bl1 noco_bl1_n noco_bl2 noco_bl2_n DP8TVar4TestArray_16X8
Xtestarray_co vss co_vdd co_wl1 co_wl2 co_bl1 co_bl1_n co_bl2 co_bl2_n co_bit co_bit_n DP8TVar4TestArray_16X8C
.ends DP8TVar4

.subckt SP6TVar5Cell wl bl bl_n vdd vss
Xpu1 vdd bit_n bit vdd sg13_lv_pmos l=1.3e-07 w=2e-07
Xpd1 bit bit_n vss vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpu2 vdd bit bit_n vdd sg13_lv_pmos l=1.3e-07 w=2e-07
Xpd2 bit_n bit vss vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg1 bit wl bl vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg2 bit_n wl bl_n vss sg13_lv_nmos l=1.3e-07 w=2e-07
.ends SP6TVar5Cell

.subckt SP6TVar5Array_2X1 vss vdd wl[0] wl[1] bl[0] bl_n[0]
Xinst0x0 wl[0] bl[0] bl_n[0] vdd vss SP6TVar5Cell
Xinst1x0 wl[1] bl[0] bl_n[0] vdd vss SP6TVar5Cell
.ends SP6TVar5Array_2X1

.subckt SP6TVar5Array_2X2 vss vdd wl[0] wl[1] bl[0] bl_n[0] bl[1] bl_n[1]
Xinst0x0 vss vdd wl[0] wl[1] bl[0] bl_n[0] SP6TVar5Array_2X1
Xinst0x1 vss vdd wl[0] wl[1] bl[1] bl_n[1] SP6TVar5Array_2X1
.ends SP6TVar5Array_2X2

.subckt SP6TVar5Array_4X2 vss vdd wl[0] wl[1] wl[2] wl[3] bl[0] bl_n[0] bl[1] bl_n[1]
Xinst0x0 vss vdd wl[0] wl[1] bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar5Array_2X2
Xinst1x0 vss vdd wl[2] wl[3] bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar5Array_2X2
.ends SP6TVar5Array_4X2

.subckt SP6TVar5Array_4X4 vss vdd wl[0] wl[1] wl[2] wl[3] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar5Array_4X2
Xinst0x1 vss vdd wl[0] wl[1] wl[2] wl[3] bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar5Array_4X2
.ends SP6TVar5Array_4X4

.subckt SP6TVar5Array_8X4 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar5Array_4X4
Xinst1x0 vss vdd wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar5Array_4X4
.ends SP6TVar5Array_8X4

.subckt SP6TVar5Array_8X8 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar5Array_8X4
Xinst0x1 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7] SP6TVar5Array_8X4
.ends SP6TVar5Array_8X8

.subckt SP6TVar5BulkConn vdd vss bl bl_n
.ends SP6TVar5BulkConn

.subckt SP6TVar5BulkConnRow_2 vss vdd bl[0] bl_n[0] bl[1] bl_n[1]
Xinst0 vdd vss bl[0] bl_n[0] SP6TVar5BulkConn
Xinst1 vdd vss bl[1] bl_n[1] SP6TVar5BulkConn
.ends SP6TVar5BulkConnRow_2

.subckt SP6TVar5BulkConnRow_4 vss vdd bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3]
Xinst0 vss vdd bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar5BulkConnRow_2
Xinst1 vss vdd bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar5BulkConnRow_2
.ends SP6TVar5BulkConnRow_4

.subckt SP6TVar5BulkConnRow_8 vss vdd bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7]
Xinst0 vss vdd bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar5BulkConnRow_4
Xinst1 vss vdd bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7] SP6TVar5BulkConnRow_4
.ends SP6TVar5BulkConnRow_8

.subckt SP6TVar5Array_16X8BC vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7] SP6TVar5Array_8X8
Xinst1x0 vss vdd wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7] SP6TVar5Array_8X8
Xbottombcrow vss vdd bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7] SP6TVar5BulkConnRow_8
Xtopbcrow vss vdd bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7] SP6TVar5BulkConnRow_8
.ends SP6TVar5Array_16X8BC

.subckt SP6TVar5TestArray_16X8 vss vdd bl bl_n wl
Xarray vss vdd zero zero zero zero zero zero zero zero wl zero zero zero zero zero zero zero bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl bl_n bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7] SP6TVar5Array_16X8BC
Xzero vdd vss zero zero_x1
.ends SP6TVar5TestArray_16X8

.subckt SP6TVar5Array_4X1 vss vdd wl[0] wl[1] wl[2] wl[3] bl[0] bl_n[0]
Xinst0x0 vss vdd wl[0] wl[1] bl[0] bl_n[0] SP6TVar5Array_2X1
Xinst1x0 vss vdd wl[2] wl[3] bl[0] bl_n[0] SP6TVar5Array_2X1
.ends SP6TVar5Array_4X1

.subckt SP6TVar5Array_8X1 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] bl[0] bl_n[0] SP6TVar5Array_4X1
Xinst1x0 vss vdd wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] SP6TVar5Array_4X1
.ends SP6TVar5Array_8X1

.subckt SP6TVar5Array_16X1BC vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] bl[0] bl_n[0]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] SP6TVar5Array_8X1
Xinst1x0 vss vdd wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] bl[0] bl_n[0] SP6TVar5Array_8X1
Xbottombcrow vdd vss bl[0] bl_n[0] SP6TVar5BulkConn
Xtopbcrow vdd vss bl[0] bl_n[0] SP6TVar5BulkConn
.ends SP6TVar5Array_16X1BC

.subckt SP6TVar5Array_8X2 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar5Array_4X2
Xinst1x0 vss vdd wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar5Array_4X2
.ends SP6TVar5Array_8X2

.subckt SP6TVar5Array_16X2BC vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] bl[0] bl_n[0] bl[1] bl_n[1]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar5Array_8X2
Xinst1x0 vss vdd wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar5Array_8X2
Xbottombcrow vss vdd bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar5BulkConnRow_2
Xtopbcrow vss vdd bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar5BulkConnRow_2
.ends SP6TVar5Array_16X2BC

.subckt SP6TVar5Array_16X4BC vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar5Array_8X4
Xinst1x0 vss vdd wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar5Array_8X4
Xbottombcrow vss vdd bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar5BulkConnRow_4
Xtopbcrow vss vdd bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar5BulkConnRow_4
.ends SP6TVar5Array_16X4BC

.subckt SP6TVar5Array_6X1 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] bl[0] bl_n[0]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] bl[0] bl_n[0] SP6TVar5Array_4X1
Xinst1x0 vss vdd wl[4] wl[5] bl[0] bl_n[0] SP6TVar5Array_2X1
.ends SP6TVar5Array_6X1

.subckt SP6TVar5CellConnectOut wl bl bl_n vdd vss bit bit_n
Xpu1 vdd bit_n bit vdd sg13_lv_pmos l=1.3e-07 w=2e-07
Xpd1 bit bit_n vss vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpu2 vdd bit bit_n vdd sg13_lv_pmos l=1.3e-07 w=2e-07
Xpd2 bit_n bit vss vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg1 bit wl bl vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg2 bit_n wl bl_n vss sg13_lv_nmos l=1.3e-07 w=2e-07
.ends SP6TVar5CellConnectOut

.subckt SP6TVar5TestArray_16X8C vss vdd bl bl_n bit bit_n wl
Xarray_0 vss vdd zero zero zero zero zero zero zero zero wl zero zero zero zero zero zero zero array_0_bl[0] array_0_bl_n[0] SP6TVar5Array_16X1BC
Xarray_1 vss vdd zero zero zero zero zero zero zero zero wl zero zero zero zero zero zero zero array_1_bl[0] array_1_bl_n[0] array_1_bl[1] array_1_bl_n[1] SP6TVar5Array_16X2BC
Xarray_2 vss vdd zero zero zero zero zero zero zero zero wl zero zero zero zero zero zero zero array_2_bl[0] array_2_bl_n[0] array_2_bl[1] array_2_bl_n[1] array_2_bl[2] array_2_bl_n[2] array_2_bl[3] array_2_bl_n[3] SP6TVar5Array_16X4BC
Xcolbc_0 vdd vss bl bl_n SP6TVar5BulkConn
Xcolbc_1 vdd vss bl bl_n SP6TVar5BulkConn
Xcolarray_0 vss vdd zero zero zero zero zero zero zero zero bl bl_n SP6TVar5Array_8X1
Xcolarray_1 vss vdd zero zero zero zero zero zero bl bl_n SP6TVar5Array_6X1
Xbc_noconn zero bl bl_n vdd vss SP6TVar5Cell
Xbc_conn wl bl bl_n vdd vss bit bit_n SP6TVar5CellConnectOut
Xzero vdd vss zero zero_x1
.ends SP6TVar5TestArray_16X8C

.subckt PadFrame_SP05 PAD0x0 PAD0x1 PAD0x2 PAD0x3 PAD0x4 PAD0x5 PAD0x6 PAD0x7 PAD0x8 PAD0x9 PAD1x0 PAD1x1 PAD1x2 PAD1x3 PAD1x4 PAD1x5 PAD1x6 PAD1x7 PAD1x8 PAD1x9
XPAD0x0 PAD0x0 BondPad
XPAD0x1 PAD0x1 BondPad
XPAD0x2 PAD0x2 BondPad
XPAD0x3 PAD0x3 BondPad
XPAD0x4 PAD0x4 BondPad
XPAD0x5 PAD0x5 BondPad
XPAD0x6 PAD0x6 BondPad
XPAD0x7 PAD0x7 BondPad
XPAD0x8 PAD0x8 BondPad
XPAD0x9 PAD0x9 BondPad
XPAD1x0 PAD1x0 BondPad
XPAD1x1 PAD1x1 BondPad
XPAD1x2 PAD1x2 BondPad
XPAD1x3 PAD1x3 BondPad
XPAD1x4 PAD1x4 BondPad
XPAD1x5 PAD1x5 BondPad
XPAD1x6 PAD1x6 BondPad
XPAD1x7 PAD1x7 BondPad
XPAD1x8 PAD1x8 BondPad
XPAD1x9 PAD1x9 BondPad
.ends PadFrame_SP05

.subckt SP6TVar5 vss noco_vdd noco_wl noco_bl noco_bl_n co_vdd co_bl co_bl_n co_bit co_bit_n co_wl
Xframe noco_vdd noco_wl NoConn_PAD0x2 co_vdd co_bl_n co_bit co_bit_n NoConn_PAD0x7 NoConn_PAD0x8 NoConn_PAD0x9 vss noco_bl noco_bl_n vss co_bl co_wl NoConn_PAD1x6 NoConn_PAD1x7 NoConn_PAD1x8 NoConn_PAD1x9 PadFrame_SP05
Xtestarray_noco vss noco_vdd noco_bl noco_bl_n noco_wl SP6TVar5TestArray_16X8
Xtestarray_co vss co_vdd co_bl co_bl_n co_bit co_bit_n co_wl SP6TVar5TestArray_16X8C
.ends SP6TVar5

.subckt DP8TVar5Cell wl1 wl2 bl1 bl1_n bl2 bl2_n vdd vss
Xpu1 vdd bit_n bit vdd sg13_lv_pmos l=1.3e-07 w=2e-07
Xpd1 bit bit_n vss vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpu2 vdd bit bit_n vdd sg13_lv_pmos l=1.3e-07 w=2e-07
Xpd2 bit_n bit vss vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg1 bit wl1 bl1 vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg1n bit_n wl1 bl1_n vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg2 bit wl2 bl2 vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg2n bit_n wl2 bl2_n vss sg13_lv_nmos l=1.3e-07 w=2e-07
.ends DP8TVar5Cell

.subckt DP8TVar5Array_2X1 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0]
Xinst0x0 wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] vdd vss DP8TVar5Cell
Xinst1x0 wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0] vdd vss DP8TVar5Cell
.ends DP8TVar5Array_2X1

.subckt DP8TVar5Array_2X2 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0] DP8TVar5Array_2X1
Xinst0x1 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TVar5Array_2X1
.ends DP8TVar5Array_2X2

.subckt DP8TVar5Array_4X2 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TVar5Array_2X2
Xinst1x0 vss vdd wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TVar5Array_2X2
.ends DP8TVar5Array_4X2

.subckt DP8TVar5Array_4X4 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TVar5Array_4X2
Xinst0x1 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar5Array_4X2
.ends DP8TVar5Array_4X4

.subckt DP8TVar5Array_8X4 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar5Array_4X4
Xinst1x0 vss vdd wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar5Array_4X4
.ends DP8TVar5Array_8X4

.subckt DP8TVar5Array_8X8 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar5Array_8X4
Xinst0x1 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar5Array_8X4
.ends DP8TVar5Array_8X8

.subckt DP8TVar5BulkConn vdd vss bl1 bl2 bl1_n bl2_n
.ends DP8TVar5BulkConn

.subckt DP8TVar5BulkConnRow_2 vss vdd bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1]
Xinst0 vdd vss bl1[0] bl2[0] bl1_n[0] bl2_n[0] DP8TVar5BulkConn
Xinst1 vdd vss bl1[1] bl2[1] bl1_n[1] bl2_n[1] DP8TVar5BulkConn
.ends DP8TVar5BulkConnRow_2

.subckt DP8TVar5BulkConnRow_4 vss vdd bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3]
Xinst0 vss vdd bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TVar5BulkConnRow_2
Xinst1 vss vdd bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar5BulkConnRow_2
.ends DP8TVar5BulkConnRow_4

.subckt DP8TVar5BulkConnRow_8 vss vdd bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0 vss vdd bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar5BulkConnRow_4
Xinst1 vss vdd bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar5BulkConnRow_4
.ends DP8TVar5BulkConnRow_8

.subckt DP8TVar5Array_16X8BC vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] wl1[8] wl2[8] wl1[9] wl2[9] wl1[10] wl2[10] wl1[11] wl2[11] wl1[12] wl2[12] wl1[13] wl2[13] wl1[14] wl2[14] wl1[15] wl2[15] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar5Array_8X8
Xinst1x0 vss vdd wl1[8] wl2[8] wl1[9] wl2[9] wl1[10] wl2[10] wl1[11] wl2[11] wl1[12] wl2[12] wl1[13] wl2[13] wl1[14] wl2[14] wl1[15] wl2[15] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar5Array_8X8
Xbottombcrow vss vdd bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar5BulkConnRow_8
Xtopbcrow vss vdd bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar5BulkConnRow_8
.ends DP8TVar5Array_16X8BC

.subckt DP8TVar5TestArray_16X8 vss vdd wl1 wl2 bl1 bl1_n bl2 bl2_n
Xarray vss vdd zero zero zero zero zero zero zero zero zero zero zero zero zero zero zero zero wl1 wl2 zero zero zero zero zero zero zero zero zero zero zero zero zero zero bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1 bl1_n bl2 bl2_n bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar5Array_16X8BC
Xzero vdd vss zero zero_x1
.ends DP8TVar5TestArray_16X8

.subckt DP8TVar5Array_4X8 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar5Array_4X4
Xinst0x1 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar5Array_4X4
.ends DP8TVar5Array_4X8

.subckt DP8TVar5Array_2X4 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TVar5Array_2X2
Xinst0x1 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar5Array_2X2
.ends DP8TVar5Array_2X4

.subckt DP8TVar5Array_2X8 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar5Array_2X4
Xinst0x1 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar5Array_2X4
.ends DP8TVar5Array_2X8

.subckt DP8TVar5Array_1X2 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1]
Xinst0x0 wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] vdd vss DP8TVar5Cell
Xinst0x1 wl1[0] wl2[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] vdd vss DP8TVar5Cell
.ends DP8TVar5Array_1X2

.subckt DP8TVar5Array_1X4 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3]
Xinst0x0 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TVar5Array_1X2
Xinst0x1 vss vdd wl1[0] wl2[0] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar5Array_1X2
.ends DP8TVar5Array_1X4

.subckt DP8TVar5Array_1X8 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar5Array_1X4
Xinst0x1 vss vdd wl1[0] wl2[0] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar5Array_1X4
.ends DP8TVar5Array_1X8

.subckt DP8TVar5Array_7X8 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar5Array_4X8
Xinst1x0 vss vdd wl1[4] wl2[4] wl1[5] wl2[5] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar5Array_2X8
Xinst2x0 vss vdd wl1[6] wl2[6] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar5Array_1X8
.ends DP8TVar5Array_7X8

.subckt DP8TVar5CellShWL1 wl1 wl2 bl1 bl1_n bl2 bl2_n vdd vss
Xpu1 vdd bit_n bit vdd sg13_lv_pmos l=1.3e-07 w=2e-07
Xpd1 bit bit_n vss vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpu2 vdd bit bit_n vdd sg13_lv_pmos l=1.3e-07 w=2e-07
Xpd2 bit_n bit vss vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg1 bit wl1 bl1 vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg1n bit_n wl1 bl1_n vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg2 bit wl1 bl2 vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg2n bit_n wl1 bl2_n vss sg13_lv_nmos l=1.3e-07 w=2e-07
.ends DP8TVar5CellShWL1

.subckt DP8TVar5ArrayShWL1_1X2 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1]
Xinst0x0 wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] vdd vss DP8TVar5CellShWL1
Xinst0x1 wl1[0] wl2[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] vdd vss DP8TVar5CellShWL1
.ends DP8TVar5ArrayShWL1_1X2

.subckt DP8TVar5ArrayShWL1_1X4 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3]
Xinst0x0 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TVar5ArrayShWL1_1X2
Xinst0x1 vss vdd wl1[0] wl2[0] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar5ArrayShWL1_1X2
.ends DP8TVar5ArrayShWL1_1X4

.subckt DP8TVar5ArrayShWL1_1X8 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar5ArrayShWL1_1X4
Xinst0x1 vss vdd wl1[0] wl2[0] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar5ArrayShWL1_1X4
.ends DP8TVar5ArrayShWL1_1X8

.subckt DP8TVar5CellConnectOut wl1 wl2 bl1 bl1_n bl2 bl2_n vdd vss bit bit_n
Xpu1 vdd bit_n bit vdd sg13_lv_pmos l=1.3e-07 w=2e-07
Xpd1 bit bit_n vss vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpu2 vdd bit bit_n vdd sg13_lv_pmos l=1.3e-07 w=2e-07
Xpd2 bit_n bit vss vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg1 bit wl1 bl1 vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg1n bit_n wl1 bl1_n vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg2 bit wl2 bl2 vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg2n bit_n wl2 bl2_n vss sg13_lv_nmos l=1.3e-07 w=2e-07
.ends DP8TVar5CellConnectOut

.subckt DP8TVar5CellShWL2 wl1 wl2 bl1 bl1_n bl2 bl2_n vdd vss
Xpu1 vdd bit_n bit vdd sg13_lv_pmos l=1.3e-07 w=2e-07
Xpd1 bit bit_n vss vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpu2 vdd bit bit_n vdd sg13_lv_pmos l=1.3e-07 w=2e-07
Xpd2 bit_n bit vss vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg1 bit wl2 bl1 vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg1n bit_n wl2 bl1_n vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg2 bit wl2 bl2 vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg2n bit_n wl2 bl2_n vss sg13_lv_nmos l=1.3e-07 w=2e-07
.ends DP8TVar5CellShWL2

.subckt DP8TVar5ArrayShWL2_1X2 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1]
Xinst0x0 wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] vdd vss DP8TVar5CellShWL2
Xinst0x1 wl1[0] wl2[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] vdd vss DP8TVar5CellShWL2
.ends DP8TVar5ArrayShWL2_1X2

.subckt DP8TVar5ArrayShWL2_1X4 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3]
Xinst0x0 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TVar5ArrayShWL2_1X2
Xinst0x1 vss vdd wl1[0] wl2[0] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar5ArrayShWL2_1X2
.ends DP8TVar5ArrayShWL2_1X4

.subckt DP8TVar5ArrayShWL2_1X8 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar5ArrayShWL2_1X4
Xinst0x1 vss vdd wl1[0] wl2[0] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar5ArrayShWL2_1X4
.ends DP8TVar5ArrayShWL2_1X8

.subckt DP8TVar5Array_6X8 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar5Array_4X8
Xinst1x0 vss vdd wl1[4] wl2[4] wl1[5] wl2[5] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar5Array_2X8
.ends DP8TVar5Array_6X8

.subckt DP8TVar5TestArray_16X8C vss vdd wl1 wl2 bl1 bl1_n bl2 bl2_n bit bit_n
Xbcconn_bot vss vdd bcconn_bot_bl1[0] bcconn_bot_bl1_n[0] bcconn_bot_bl2[0] bcconn_bot_bl2_n[0] bcconn_bot_bl1[1] bcconn_bot_bl1_n[1] bcconn_bot_bl2[1] bcconn_bot_bl2_n[1] bcconn_bot_bl1[2] bcconn_bot_bl1_n[2] bcconn_bot_bl2[2] bcconn_bot_bl2_n[2] bcconn_bot_bl1[3] bcconn_bot_bl1_n[3] bcconn_bot_bl2[3] bcconn_bot_bl2_n[3] bl1 bl1_n bl2 bl2_n bcconn_bot_bl1[5] bcconn_bot_bl1_n[5] bcconn_bot_bl2[5] bcconn_bot_bl2_n[5] bcconn_bot_bl1[6] bcconn_bot_bl1_n[6] bcconn_bot_bl2[6] bcconn_bot_bl2_n[6] bcconn_bot_bl1[7] bcconn_bot_bl1_n[7] bcconn_bot_bl2[7] bcconn_bot_bl2_n[7] DP8TVar5BulkConnRow_8
Xbcconn_top vss vdd bcconn_top_bl1[0] bcconn_top_bl1_n[0] bcconn_top_bl2[0] bcconn_top_bl2_n[0] bcconn_top_bl1[1] bcconn_top_bl1_n[1] bcconn_top_bl2[1] bcconn_top_bl2_n[1] bcconn_top_bl1[2] bcconn_top_bl1_n[2] bcconn_top_bl2[2] bcconn_top_bl2_n[2] bcconn_top_bl1[3] bcconn_top_bl1_n[3] bcconn_top_bl2[3] bcconn_top_bl2_n[3] bl1 bl1_n bl2 bl2_n bcconn_top_bl1[5] bcconn_top_bl1_n[5] bcconn_top_bl2[5] bcconn_top_bl2_n[5] bcconn_top_bl1[6] bcconn_top_bl1_n[6] bcconn_top_bl2[6] bcconn_top_bl2_n[6] bcconn_top_bl1[7] bcconn_top_bl1_n[7] bcconn_top_bl2[7] bcconn_top_bl2_n[7] DP8TVar5BulkConnRow_8
Xarray_bot vss vdd zero zero zero zero zero zero zero zero zero zero zero zero zero zero array_bot_bl1[0] array_bot_bl1_n[0] array_bot_bl2[0] array_bot_bl2_n[0] array_bot_bl1[1] array_bot_bl1_n[1] array_bot_bl2[1] array_bot_bl2_n[1] array_bot_bl1[2] array_bot_bl1_n[2] array_bot_bl2[2] array_bot_bl2_n[2] array_bot_bl1[3] array_bot_bl1_n[3] array_bot_bl2[3] array_bot_bl2_n[3] bl1 bl1_n bl2 bl2_n array_bot_bl1[5] array_bot_bl1_n[5] array_bot_bl2[5] array_bot_bl2_n[5] array_bot_bl1[6] array_bot_bl1_n[6] array_bot_bl2[6] array_bot_bl2_n[6] array_bot_bl1[7] array_bot_bl1_n[7] array_bot_bl2[7] array_bot_bl2_n[7] DP8TVar5Array_7X8
Xshwl1_row vss vdd zero bit shwl1_row_bl1[0] shwl1_row_bl1_n[0] shwl1_row_bl2[0] shwl1_row_bl2_n[0] shwl1_row_bl1[1] shwl1_row_bl1_n[1] shwl1_row_bl2[1] shwl1_row_bl2_n[1] shwl1_row_bl1[2] shwl1_row_bl1_n[2] shwl1_row_bl2[2] shwl1_row_bl2_n[2] shwl1_row_bl1[3] shwl1_row_bl1_n[3] shwl1_row_bl2[3] shwl1_row_bl2_n[3] bl1 bl1_n bl2 bl2_n shwl1_row_bl1[5] shwl1_row_bl1_n[5] shwl1_row_bl2[5] shwl1_row_bl2_n[5] shwl1_row_bl1[6] shwl1_row_bl1_n[6] shwl1_row_bl2[6] shwl1_row_bl2_n[6] shwl1_row_bl1[7] shwl1_row_bl1_n[7] shwl1_row_bl2[7] shwl1_row_bl2_n[7] DP8TVar5ArrayShWL1_1X8
Xcell_cols_left vss vdd wl1 wl2 cell_cols_left_bl1[0] cell_cols_left_bl1_n[0] cell_cols_left_bl2[0] cell_cols_left_bl2_n[0] cell_cols_left_bl1[1] cell_cols_left_bl1_n[1] cell_cols_left_bl2[1] cell_cols_left_bl2_n[1] cell_cols_left_bl1[2] cell_cols_left_bl1_n[2] cell_cols_left_bl2[2] cell_cols_left_bl2_n[2] cell_cols_left_bl1[3] cell_cols_left_bl1_n[3] cell_cols_left_bl2[3] cell_cols_left_bl2_n[3] DP8TVar5Array_1X4
Xconncell wl1 wl2 bl1 bl1_n bl2 bl2_n vdd vss bit bit_n DP8TVar5CellConnectOut
Xfillcell wl1 wl2 fillcell_bl1 fillcell_bl1_n fillcell_bl2 fillcell_bl2_n vdd vss DP8TVar5Cell
Xcell_cols_right vss vdd wl1 wl2 cell_cols_right_bl1[0] cell_cols_right_bl1_n[0] cell_cols_right_bl2[0] cell_cols_right_bl2_n[0] cell_cols_right_bl1[1] cell_cols_right_bl1_n[1] cell_cols_right_bl2[1] cell_cols_right_bl2_n[1] DP8TVar5Array_1X2
Xshwl2_row vss vdd bit_n zero shwl2_row_bl1[0] shwl2_row_bl1_n[0] shwl2_row_bl2[0] shwl2_row_bl2_n[0] shwl2_row_bl1[1] shwl2_row_bl1_n[1] shwl2_row_bl2[1] shwl2_row_bl2_n[1] shwl2_row_bl1[2] shwl2_row_bl1_n[2] shwl2_row_bl2[2] shwl2_row_bl2_n[2] shwl2_row_bl1[3] shwl2_row_bl1_n[3] shwl2_row_bl2[3] shwl2_row_bl2_n[3] bl1 bl1_n bl2 bl2_n shwl2_row_bl1[5] shwl2_row_bl1_n[5] shwl2_row_bl2[5] shwl2_row_bl2_n[5] shwl2_row_bl1[6] shwl2_row_bl1_n[6] shwl2_row_bl2[6] shwl2_row_bl2_n[6] shwl2_row_bl1[7] shwl2_row_bl1_n[7] shwl2_row_bl2[7] shwl2_row_bl2_n[7] DP8TVar5ArrayShWL2_1X8
Xarray_top vss vdd zero zero zero zero zero zero zero zero zero zero zero zero array_top_bl1[0] array_top_bl1_n[0] array_top_bl2[0] array_top_bl2_n[0] array_top_bl1[1] array_top_bl1_n[1] array_top_bl2[1] array_top_bl2_n[1] array_top_bl1[2] array_top_bl1_n[2] array_top_bl2[2] array_top_bl2_n[2] array_top_bl1[3] array_top_bl1_n[3] array_top_bl2[3] array_top_bl2_n[3] bl1 bl1_n bl2 bl2_n array_top_bl1[5] array_top_bl1_n[5] array_top_bl2[5] array_top_bl2_n[5] array_top_bl1[6] array_top_bl1_n[6] array_top_bl2[6] array_top_bl2_n[6] array_top_bl1[7] array_top_bl1_n[7] array_top_bl2[7] array_top_bl2_n[7] DP8TVar5Array_6X8
Xzero vdd vss zero zero_x1
.ends DP8TVar5TestArray_16X8C

.subckt PadFrame_DP05 PAD0x0 PAD0x1 PAD0x2 PAD0x3 PAD0x4 PAD0x5 PAD0x6 PAD0x7 PAD0x8 PAD0x9 PAD1x0 PAD1x1 PAD1x2 PAD1x3 PAD1x4 PAD1x5 PAD1x6 PAD1x7 PAD1x8 PAD1x9
XPAD0x0 PAD0x0 BondPad
XPAD0x1 PAD0x1 BondPad
XPAD0x2 PAD0x2 BondPad
XPAD0x3 PAD0x3 BondPad
XPAD0x4 PAD0x4 BondPad
XPAD0x5 PAD0x5 BondPad
XPAD0x6 PAD0x6 BondPad
XPAD0x7 PAD0x7 BondPad
XPAD0x8 PAD0x8 BondPad
XPAD0x9 PAD0x9 BondPad
XPAD1x0 PAD1x0 BondPad
XPAD1x1 PAD1x1 BondPad
XPAD1x2 PAD1x2 BondPad
XPAD1x3 PAD1x3 BondPad
XPAD1x4 PAD1x4 BondPad
XPAD1x5 PAD1x5 BondPad
XPAD1x6 PAD1x6 BondPad
XPAD1x7 PAD1x7 BondPad
XPAD1x8 PAD1x8 BondPad
XPAD1x9 PAD1x9 BondPad
.ends PadFrame_DP05

.subckt DP8TVar5 vss noco_vdd noco_wl1 noco_wl2 noco_bl1 noco_bl1_n noco_bl2 noco_bl2_n co_vdd co_bit co_bit_n co_wl1 co_wl2 co_bl1 co_bl1_n co_bl2_n co_bl2
Xframe noco_vdd noco_wl1 noco_wl2 noco_bl2 co_vdd co_bit co_bit_n co_wl1 co_wl2 NoConn_PAD0x9 vss noco_bl1 noco_bl1_n noco_bl2_n vss co_bl1 co_bl1_n co_bl2_n co_bl2 NoConn_PAD1x9 PadFrame_DP05
Xtestarray_noco vss noco_vdd noco_wl1 noco_wl2 noco_bl1 noco_bl1_n noco_bl2 noco_bl2_n DP8TVar5TestArray_16X8
Xtestarray_co vss co_vdd co_wl1 co_wl2 co_bl1 co_bl1_n co_bl2 co_bl2_n co_bit co_bit_n DP8TVar5TestArray_16X8C
.ends DP8TVar5

.subckt SP6TVar6Cell wl bl bl_n vdd vss
Xpu1 vdd bit_n bit vdd sg13_lv_pmos l=1.3e-07 w=1.5e-07
Xpd1 bit bit_n vss vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpu2 vdd bit bit_n vdd sg13_lv_pmos l=1.3e-07 w=1.5e-07
Xpd2 bit_n bit vss vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg1 bit wl bl vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg2 bit_n wl bl_n vss sg13_lv_nmos l=1.3e-07 w=2e-07
.ends SP6TVar6Cell

.subckt SP6TVar6Array_2X1 vss vdd wl[0] wl[1] bl[0] bl_n[0]
Xinst0x0 wl[0] bl[0] bl_n[0] vdd vss SP6TVar6Cell
Xinst1x0 wl[1] bl[0] bl_n[0] vdd vss SP6TVar6Cell
.ends SP6TVar6Array_2X1

.subckt SP6TVar6Array_2X2 vss vdd wl[0] wl[1] bl[0] bl_n[0] bl[1] bl_n[1]
Xinst0x0 vss vdd wl[0] wl[1] bl[0] bl_n[0] SP6TVar6Array_2X1
Xinst0x1 vss vdd wl[0] wl[1] bl[1] bl_n[1] SP6TVar6Array_2X1
.ends SP6TVar6Array_2X2

.subckt SP6TVar6Array_4X2 vss vdd wl[0] wl[1] wl[2] wl[3] bl[0] bl_n[0] bl[1] bl_n[1]
Xinst0x0 vss vdd wl[0] wl[1] bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar6Array_2X2
Xinst1x0 vss vdd wl[2] wl[3] bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar6Array_2X2
.ends SP6TVar6Array_4X2

.subckt SP6TVar6Array_4X4 vss vdd wl[0] wl[1] wl[2] wl[3] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar6Array_4X2
Xinst0x1 vss vdd wl[0] wl[1] wl[2] wl[3] bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar6Array_4X2
.ends SP6TVar6Array_4X4

.subckt SP6TVar6Array_8X4 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar6Array_4X4
Xinst1x0 vss vdd wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar6Array_4X4
.ends SP6TVar6Array_8X4

.subckt SP6TVar6Array_8X8 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar6Array_8X4
Xinst0x1 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7] SP6TVar6Array_8X4
.ends SP6TVar6Array_8X8

.subckt SP6TVar6BulkConn vdd vss bl bl_n
.ends SP6TVar6BulkConn

.subckt SP6TVar6BulkConnRow_2 vss vdd bl[0] bl_n[0] bl[1] bl_n[1]
Xinst0 vdd vss bl[0] bl_n[0] SP6TVar6BulkConn
Xinst1 vdd vss bl[1] bl_n[1] SP6TVar6BulkConn
.ends SP6TVar6BulkConnRow_2

.subckt SP6TVar6BulkConnRow_4 vss vdd bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3]
Xinst0 vss vdd bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar6BulkConnRow_2
Xinst1 vss vdd bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar6BulkConnRow_2
.ends SP6TVar6BulkConnRow_4

.subckt SP6TVar6BulkConnRow_8 vss vdd bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7]
Xinst0 vss vdd bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar6BulkConnRow_4
Xinst1 vss vdd bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7] SP6TVar6BulkConnRow_4
.ends SP6TVar6BulkConnRow_8

.subckt SP6TVar6Array_16X8BC vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7] SP6TVar6Array_8X8
Xinst1x0 vss vdd wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7] SP6TVar6Array_8X8
Xbottombcrow vss vdd bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7] SP6TVar6BulkConnRow_8
Xtopbcrow vss vdd bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7] SP6TVar6BulkConnRow_8
.ends SP6TVar6Array_16X8BC

.subckt SP6TVar6TestArray_16X8 vss vdd bl bl_n wl
Xarray vss vdd zero zero zero zero zero zero zero zero wl zero zero zero zero zero zero zero bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl bl_n bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7] SP6TVar6Array_16X8BC
Xzero vdd vss zero zero_x1
.ends SP6TVar6TestArray_16X8

.subckt SP6TVar6Array_4X1 vss vdd wl[0] wl[1] wl[2] wl[3] bl[0] bl_n[0]
Xinst0x0 vss vdd wl[0] wl[1] bl[0] bl_n[0] SP6TVar6Array_2X1
Xinst1x0 vss vdd wl[2] wl[3] bl[0] bl_n[0] SP6TVar6Array_2X1
.ends SP6TVar6Array_4X1

.subckt SP6TVar6Array_8X1 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] bl[0] bl_n[0] SP6TVar6Array_4X1
Xinst1x0 vss vdd wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] SP6TVar6Array_4X1
.ends SP6TVar6Array_8X1

.subckt SP6TVar6Array_16X1BC vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] bl[0] bl_n[0]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] SP6TVar6Array_8X1
Xinst1x0 vss vdd wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] bl[0] bl_n[0] SP6TVar6Array_8X1
Xbottombcrow vdd vss bl[0] bl_n[0] SP6TVar6BulkConn
Xtopbcrow vdd vss bl[0] bl_n[0] SP6TVar6BulkConn
.ends SP6TVar6Array_16X1BC

.subckt SP6TVar6Array_8X2 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar6Array_4X2
Xinst1x0 vss vdd wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar6Array_4X2
.ends SP6TVar6Array_8X2

.subckt SP6TVar6Array_16X2BC vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] bl[0] bl_n[0] bl[1] bl_n[1]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar6Array_8X2
Xinst1x0 vss vdd wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar6Array_8X2
Xbottombcrow vss vdd bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar6BulkConnRow_2
Xtopbcrow vss vdd bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar6BulkConnRow_2
.ends SP6TVar6Array_16X2BC

.subckt SP6TVar6Array_16X4BC vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar6Array_8X4
Xinst1x0 vss vdd wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar6Array_8X4
Xbottombcrow vss vdd bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar6BulkConnRow_4
Xtopbcrow vss vdd bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar6BulkConnRow_4
.ends SP6TVar6Array_16X4BC

.subckt SP6TVar6Array_6X1 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] bl[0] bl_n[0]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] bl[0] bl_n[0] SP6TVar6Array_4X1
Xinst1x0 vss vdd wl[4] wl[5] bl[0] bl_n[0] SP6TVar6Array_2X1
.ends SP6TVar6Array_6X1

.subckt SP6TVar6CellConnectOut wl bl bl_n vdd vss bit bit_n
Xpu1 vdd bit_n bit vdd sg13_lv_pmos l=1.3e-07 w=1.5e-07
Xpd1 bit bit_n vss vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpu2 vdd bit bit_n vdd sg13_lv_pmos l=1.3e-07 w=1.5e-07
Xpd2 bit_n bit vss vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg1 bit wl bl vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg2 bit_n wl bl_n vss sg13_lv_nmos l=1.3e-07 w=2e-07
.ends SP6TVar6CellConnectOut

.subckt SP6TVar6TestArray_16X8C vss vdd bl bl_n bit bit_n wl
Xarray_0 vss vdd zero zero zero zero zero zero zero zero wl zero zero zero zero zero zero zero array_0_bl[0] array_0_bl_n[0] SP6TVar6Array_16X1BC
Xarray_1 vss vdd zero zero zero zero zero zero zero zero wl zero zero zero zero zero zero zero array_1_bl[0] array_1_bl_n[0] array_1_bl[1] array_1_bl_n[1] SP6TVar6Array_16X2BC
Xarray_2 vss vdd zero zero zero zero zero zero zero zero wl zero zero zero zero zero zero zero array_2_bl[0] array_2_bl_n[0] array_2_bl[1] array_2_bl_n[1] array_2_bl[2] array_2_bl_n[2] array_2_bl[3] array_2_bl_n[3] SP6TVar6Array_16X4BC
Xcolbc_0 vdd vss bl bl_n SP6TVar6BulkConn
Xcolbc_1 vdd vss bl bl_n SP6TVar6BulkConn
Xcolarray_0 vss vdd zero zero zero zero zero zero zero zero bl bl_n SP6TVar6Array_8X1
Xcolarray_1 vss vdd zero zero zero zero zero zero bl bl_n SP6TVar6Array_6X1
Xbc_noconn zero bl bl_n vdd vss SP6TVar6Cell
Xbc_conn wl bl bl_n vdd vss bit bit_n SP6TVar6CellConnectOut
Xzero vdd vss zero zero_x1
.ends SP6TVar6TestArray_16X8C

.subckt PadFrame_SP06 PAD0x0 PAD0x1 PAD0x2 PAD0x3 PAD0x4 PAD0x5 PAD0x6 PAD0x7 PAD0x8 PAD0x9 PAD1x0 PAD1x1 PAD1x2 PAD1x3 PAD1x4 PAD1x5 PAD1x6 PAD1x7 PAD1x8 PAD1x9
XPAD0x0 PAD0x0 BondPad
XPAD0x1 PAD0x1 BondPad
XPAD0x2 PAD0x2 BondPad
XPAD0x3 PAD0x3 BondPad
XPAD0x4 PAD0x4 BondPad
XPAD0x5 PAD0x5 BondPad
XPAD0x6 PAD0x6 BondPad
XPAD0x7 PAD0x7 BondPad
XPAD0x8 PAD0x8 BondPad
XPAD0x9 PAD0x9 BondPad
XPAD1x0 PAD1x0 BondPad
XPAD1x1 PAD1x1 BondPad
XPAD1x2 PAD1x2 BondPad
XPAD1x3 PAD1x3 BondPad
XPAD1x4 PAD1x4 BondPad
XPAD1x5 PAD1x5 BondPad
XPAD1x6 PAD1x6 BondPad
XPAD1x7 PAD1x7 BondPad
XPAD1x8 PAD1x8 BondPad
XPAD1x9 PAD1x9 BondPad
.ends PadFrame_SP06

.subckt SP6TVar6 vss noco_vdd noco_wl noco_bl noco_bl_n co_vdd co_bl co_bl_n co_bit co_bit_n co_wl
Xframe noco_vdd noco_wl NoConn_PAD0x2 co_vdd co_bl_n co_bit co_bit_n NoConn_PAD0x7 NoConn_PAD0x8 NoConn_PAD0x9 vss noco_bl noco_bl_n vss co_bl co_wl NoConn_PAD1x6 NoConn_PAD1x7 NoConn_PAD1x8 NoConn_PAD1x9 PadFrame_SP06
Xtestarray_noco vss noco_vdd noco_bl noco_bl_n noco_wl SP6TVar6TestArray_16X8
Xtestarray_co vss co_vdd co_bl co_bl_n co_bit co_bit_n co_wl SP6TVar6TestArray_16X8C
.ends SP6TVar6

.subckt DP8TVar6Cell wl1 wl2 bl1 bl1_n bl2 bl2_n vdd vss
Xpu1 vdd bit_n bit vdd sg13_lv_pmos l=1.3e-07 w=1.5e-07
Xpd1 bit bit_n vss vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpu2 vdd bit bit_n vdd sg13_lv_pmos l=1.3e-07 w=1.5e-07
Xpd2 bit_n bit vss vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg1 bit wl1 bl1 vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg1n bit_n wl1 bl1_n vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg2 bit wl2 bl2 vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg2n bit_n wl2 bl2_n vss sg13_lv_nmos l=1.3e-07 w=2e-07
.ends DP8TVar6Cell

.subckt DP8TVar6Array_2X1 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0]
Xinst0x0 wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] vdd vss DP8TVar6Cell
Xinst1x0 wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0] vdd vss DP8TVar6Cell
.ends DP8TVar6Array_2X1

.subckt DP8TVar6Array_2X2 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0] DP8TVar6Array_2X1
Xinst0x1 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TVar6Array_2X1
.ends DP8TVar6Array_2X2

.subckt DP8TVar6Array_4X2 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TVar6Array_2X2
Xinst1x0 vss vdd wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TVar6Array_2X2
.ends DP8TVar6Array_4X2

.subckt DP8TVar6Array_4X4 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TVar6Array_4X2
Xinst0x1 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar6Array_4X2
.ends DP8TVar6Array_4X4

.subckt DP8TVar6Array_8X4 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar6Array_4X4
Xinst1x0 vss vdd wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar6Array_4X4
.ends DP8TVar6Array_8X4

.subckt DP8TVar6Array_8X8 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar6Array_8X4
Xinst0x1 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar6Array_8X4
.ends DP8TVar6Array_8X8

.subckt DP8TVar6BulkConn vdd vss bl1 bl2 bl1_n bl2_n
.ends DP8TVar6BulkConn

.subckt DP8TVar6BulkConnRow_2 vss vdd bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1]
Xinst0 vdd vss bl1[0] bl2[0] bl1_n[0] bl2_n[0] DP8TVar6BulkConn
Xinst1 vdd vss bl1[1] bl2[1] bl1_n[1] bl2_n[1] DP8TVar6BulkConn
.ends DP8TVar6BulkConnRow_2

.subckt DP8TVar6BulkConnRow_4 vss vdd bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3]
Xinst0 vss vdd bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TVar6BulkConnRow_2
Xinst1 vss vdd bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar6BulkConnRow_2
.ends DP8TVar6BulkConnRow_4

.subckt DP8TVar6BulkConnRow_8 vss vdd bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0 vss vdd bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar6BulkConnRow_4
Xinst1 vss vdd bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar6BulkConnRow_4
.ends DP8TVar6BulkConnRow_8

.subckt DP8TVar6Array_16X8BC vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] wl1[8] wl2[8] wl1[9] wl2[9] wl1[10] wl2[10] wl1[11] wl2[11] wl1[12] wl2[12] wl1[13] wl2[13] wl1[14] wl2[14] wl1[15] wl2[15] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar6Array_8X8
Xinst1x0 vss vdd wl1[8] wl2[8] wl1[9] wl2[9] wl1[10] wl2[10] wl1[11] wl2[11] wl1[12] wl2[12] wl1[13] wl2[13] wl1[14] wl2[14] wl1[15] wl2[15] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar6Array_8X8
Xbottombcrow vss vdd bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar6BulkConnRow_8
Xtopbcrow vss vdd bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar6BulkConnRow_8
.ends DP8TVar6Array_16X8BC

.subckt DP8TVar6TestArray_16X8 vss vdd wl1 wl2 bl1 bl1_n bl2 bl2_n
Xarray vss vdd zero zero zero zero zero zero zero zero zero zero zero zero zero zero zero zero wl1 wl2 zero zero zero zero zero zero zero zero zero zero zero zero zero zero bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1 bl1_n bl2 bl2_n bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar6Array_16X8BC
Xzero vdd vss zero zero_x1
.ends DP8TVar6TestArray_16X8

.subckt DP8TVar6Array_4X8 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar6Array_4X4
Xinst0x1 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar6Array_4X4
.ends DP8TVar6Array_4X8

.subckt DP8TVar6Array_2X4 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TVar6Array_2X2
Xinst0x1 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar6Array_2X2
.ends DP8TVar6Array_2X4

.subckt DP8TVar6Array_2X8 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar6Array_2X4
Xinst0x1 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar6Array_2X4
.ends DP8TVar6Array_2X8

.subckt DP8TVar6Array_1X2 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1]
Xinst0x0 wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] vdd vss DP8TVar6Cell
Xinst0x1 wl1[0] wl2[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] vdd vss DP8TVar6Cell
.ends DP8TVar6Array_1X2

.subckt DP8TVar6Array_1X4 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3]
Xinst0x0 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TVar6Array_1X2
Xinst0x1 vss vdd wl1[0] wl2[0] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar6Array_1X2
.ends DP8TVar6Array_1X4

.subckt DP8TVar6Array_1X8 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar6Array_1X4
Xinst0x1 vss vdd wl1[0] wl2[0] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar6Array_1X4
.ends DP8TVar6Array_1X8

.subckt DP8TVar6Array_7X8 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar6Array_4X8
Xinst1x0 vss vdd wl1[4] wl2[4] wl1[5] wl2[5] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar6Array_2X8
Xinst2x0 vss vdd wl1[6] wl2[6] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar6Array_1X8
.ends DP8TVar6Array_7X8

.subckt DP8TVar6CellShWL1 wl1 wl2 bl1 bl1_n bl2 bl2_n vdd vss
Xpu1 vdd bit_n bit vdd sg13_lv_pmos l=1.3e-07 w=1.5e-07
Xpd1 bit bit_n vss vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpu2 vdd bit bit_n vdd sg13_lv_pmos l=1.3e-07 w=1.5e-07
Xpd2 bit_n bit vss vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg1 bit wl1 bl1 vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg1n bit_n wl1 bl1_n vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg2 bit wl1 bl2 vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg2n bit_n wl1 bl2_n vss sg13_lv_nmos l=1.3e-07 w=2e-07
.ends DP8TVar6CellShWL1

.subckt DP8TVar6ArrayShWL1_1X2 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1]
Xinst0x0 wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] vdd vss DP8TVar6CellShWL1
Xinst0x1 wl1[0] wl2[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] vdd vss DP8TVar6CellShWL1
.ends DP8TVar6ArrayShWL1_1X2

.subckt DP8TVar6ArrayShWL1_1X4 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3]
Xinst0x0 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TVar6ArrayShWL1_1X2
Xinst0x1 vss vdd wl1[0] wl2[0] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar6ArrayShWL1_1X2
.ends DP8TVar6ArrayShWL1_1X4

.subckt DP8TVar6ArrayShWL1_1X8 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar6ArrayShWL1_1X4
Xinst0x1 vss vdd wl1[0] wl2[0] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar6ArrayShWL1_1X4
.ends DP8TVar6ArrayShWL1_1X8

.subckt DP8TVar6CellConnectOut wl1 wl2 bl1 bl1_n bl2 bl2_n vdd vss bit bit_n
Xpu1 vdd bit_n bit vdd sg13_lv_pmos l=1.3e-07 w=1.5e-07
Xpd1 bit bit_n vss vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpu2 vdd bit bit_n vdd sg13_lv_pmos l=1.3e-07 w=1.5e-07
Xpd2 bit_n bit vss vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg1 bit wl1 bl1 vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg1n bit_n wl1 bl1_n vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg2 bit wl2 bl2 vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg2n bit_n wl2 bl2_n vss sg13_lv_nmos l=1.3e-07 w=2e-07
.ends DP8TVar6CellConnectOut

.subckt DP8TVar6CellShWL2 wl1 wl2 bl1 bl1_n bl2 bl2_n vdd vss
Xpu1 vdd bit_n bit vdd sg13_lv_pmos l=1.3e-07 w=1.5e-07
Xpd1 bit bit_n vss vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpu2 vdd bit bit_n vdd sg13_lv_pmos l=1.3e-07 w=1.5e-07
Xpd2 bit_n bit vss vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg1 bit wl2 bl1 vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg1n bit_n wl2 bl1_n vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg2 bit wl2 bl2 vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg2n bit_n wl2 bl2_n vss sg13_lv_nmos l=1.3e-07 w=2e-07
.ends DP8TVar6CellShWL2

.subckt DP8TVar6ArrayShWL2_1X2 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1]
Xinst0x0 wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] vdd vss DP8TVar6CellShWL2
Xinst0x1 wl1[0] wl2[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] vdd vss DP8TVar6CellShWL2
.ends DP8TVar6ArrayShWL2_1X2

.subckt DP8TVar6ArrayShWL2_1X4 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3]
Xinst0x0 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TVar6ArrayShWL2_1X2
Xinst0x1 vss vdd wl1[0] wl2[0] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar6ArrayShWL2_1X2
.ends DP8TVar6ArrayShWL2_1X4

.subckt DP8TVar6ArrayShWL2_1X8 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar6ArrayShWL2_1X4
Xinst0x1 vss vdd wl1[0] wl2[0] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar6ArrayShWL2_1X4
.ends DP8TVar6ArrayShWL2_1X8

.subckt DP8TVar6Array_6X8 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar6Array_4X8
Xinst1x0 vss vdd wl1[4] wl2[4] wl1[5] wl2[5] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar6Array_2X8
.ends DP8TVar6Array_6X8

.subckt DP8TVar6TestArray_16X8C vss vdd wl1 wl2 bl1 bl1_n bl2 bl2_n bit bit_n
Xbcconn_bot vss vdd bcconn_bot_bl1[0] bcconn_bot_bl1_n[0] bcconn_bot_bl2[0] bcconn_bot_bl2_n[0] bcconn_bot_bl1[1] bcconn_bot_bl1_n[1] bcconn_bot_bl2[1] bcconn_bot_bl2_n[1] bcconn_bot_bl1[2] bcconn_bot_bl1_n[2] bcconn_bot_bl2[2] bcconn_bot_bl2_n[2] bcconn_bot_bl1[3] bcconn_bot_bl1_n[3] bcconn_bot_bl2[3] bcconn_bot_bl2_n[3] bl1 bl1_n bl2 bl2_n bcconn_bot_bl1[5] bcconn_bot_bl1_n[5] bcconn_bot_bl2[5] bcconn_bot_bl2_n[5] bcconn_bot_bl1[6] bcconn_bot_bl1_n[6] bcconn_bot_bl2[6] bcconn_bot_bl2_n[6] bcconn_bot_bl1[7] bcconn_bot_bl1_n[7] bcconn_bot_bl2[7] bcconn_bot_bl2_n[7] DP8TVar6BulkConnRow_8
Xbcconn_top vss vdd bcconn_top_bl1[0] bcconn_top_bl1_n[0] bcconn_top_bl2[0] bcconn_top_bl2_n[0] bcconn_top_bl1[1] bcconn_top_bl1_n[1] bcconn_top_bl2[1] bcconn_top_bl2_n[1] bcconn_top_bl1[2] bcconn_top_bl1_n[2] bcconn_top_bl2[2] bcconn_top_bl2_n[2] bcconn_top_bl1[3] bcconn_top_bl1_n[3] bcconn_top_bl2[3] bcconn_top_bl2_n[3] bl1 bl1_n bl2 bl2_n bcconn_top_bl1[5] bcconn_top_bl1_n[5] bcconn_top_bl2[5] bcconn_top_bl2_n[5] bcconn_top_bl1[6] bcconn_top_bl1_n[6] bcconn_top_bl2[6] bcconn_top_bl2_n[6] bcconn_top_bl1[7] bcconn_top_bl1_n[7] bcconn_top_bl2[7] bcconn_top_bl2_n[7] DP8TVar6BulkConnRow_8
Xarray_bot vss vdd zero zero zero zero zero zero zero zero zero zero zero zero zero zero array_bot_bl1[0] array_bot_bl1_n[0] array_bot_bl2[0] array_bot_bl2_n[0] array_bot_bl1[1] array_bot_bl1_n[1] array_bot_bl2[1] array_bot_bl2_n[1] array_bot_bl1[2] array_bot_bl1_n[2] array_bot_bl2[2] array_bot_bl2_n[2] array_bot_bl1[3] array_bot_bl1_n[3] array_bot_bl2[3] array_bot_bl2_n[3] bl1 bl1_n bl2 bl2_n array_bot_bl1[5] array_bot_bl1_n[5] array_bot_bl2[5] array_bot_bl2_n[5] array_bot_bl1[6] array_bot_bl1_n[6] array_bot_bl2[6] array_bot_bl2_n[6] array_bot_bl1[7] array_bot_bl1_n[7] array_bot_bl2[7] array_bot_bl2_n[7] DP8TVar6Array_7X8
Xshwl1_row vss vdd zero bit shwl1_row_bl1[0] shwl1_row_bl1_n[0] shwl1_row_bl2[0] shwl1_row_bl2_n[0] shwl1_row_bl1[1] shwl1_row_bl1_n[1] shwl1_row_bl2[1] shwl1_row_bl2_n[1] shwl1_row_bl1[2] shwl1_row_bl1_n[2] shwl1_row_bl2[2] shwl1_row_bl2_n[2] shwl1_row_bl1[3] shwl1_row_bl1_n[3] shwl1_row_bl2[3] shwl1_row_bl2_n[3] bl1 bl1_n bl2 bl2_n shwl1_row_bl1[5] shwl1_row_bl1_n[5] shwl1_row_bl2[5] shwl1_row_bl2_n[5] shwl1_row_bl1[6] shwl1_row_bl1_n[6] shwl1_row_bl2[6] shwl1_row_bl2_n[6] shwl1_row_bl1[7] shwl1_row_bl1_n[7] shwl1_row_bl2[7] shwl1_row_bl2_n[7] DP8TVar6ArrayShWL1_1X8
Xcell_cols_left vss vdd wl1 wl2 cell_cols_left_bl1[0] cell_cols_left_bl1_n[0] cell_cols_left_bl2[0] cell_cols_left_bl2_n[0] cell_cols_left_bl1[1] cell_cols_left_bl1_n[1] cell_cols_left_bl2[1] cell_cols_left_bl2_n[1] cell_cols_left_bl1[2] cell_cols_left_bl1_n[2] cell_cols_left_bl2[2] cell_cols_left_bl2_n[2] cell_cols_left_bl1[3] cell_cols_left_bl1_n[3] cell_cols_left_bl2[3] cell_cols_left_bl2_n[3] DP8TVar6Array_1X4
Xconncell wl1 wl2 bl1 bl1_n bl2 bl2_n vdd vss bit bit_n DP8TVar6CellConnectOut
Xfillcell wl1 wl2 fillcell_bl1 fillcell_bl1_n fillcell_bl2 fillcell_bl2_n vdd vss DP8TVar6Cell
Xcell_cols_right vss vdd wl1 wl2 cell_cols_right_bl1[0] cell_cols_right_bl1_n[0] cell_cols_right_bl2[0] cell_cols_right_bl2_n[0] cell_cols_right_bl1[1] cell_cols_right_bl1_n[1] cell_cols_right_bl2[1] cell_cols_right_bl2_n[1] DP8TVar6Array_1X2
Xshwl2_row vss vdd bit_n zero shwl2_row_bl1[0] shwl2_row_bl1_n[0] shwl2_row_bl2[0] shwl2_row_bl2_n[0] shwl2_row_bl1[1] shwl2_row_bl1_n[1] shwl2_row_bl2[1] shwl2_row_bl2_n[1] shwl2_row_bl1[2] shwl2_row_bl1_n[2] shwl2_row_bl2[2] shwl2_row_bl2_n[2] shwl2_row_bl1[3] shwl2_row_bl1_n[3] shwl2_row_bl2[3] shwl2_row_bl2_n[3] bl1 bl1_n bl2 bl2_n shwl2_row_bl1[5] shwl2_row_bl1_n[5] shwl2_row_bl2[5] shwl2_row_bl2_n[5] shwl2_row_bl1[6] shwl2_row_bl1_n[6] shwl2_row_bl2[6] shwl2_row_bl2_n[6] shwl2_row_bl1[7] shwl2_row_bl1_n[7] shwl2_row_bl2[7] shwl2_row_bl2_n[7] DP8TVar6ArrayShWL2_1X8
Xarray_top vss vdd zero zero zero zero zero zero zero zero zero zero zero zero array_top_bl1[0] array_top_bl1_n[0] array_top_bl2[0] array_top_bl2_n[0] array_top_bl1[1] array_top_bl1_n[1] array_top_bl2[1] array_top_bl2_n[1] array_top_bl1[2] array_top_bl1_n[2] array_top_bl2[2] array_top_bl2_n[2] array_top_bl1[3] array_top_bl1_n[3] array_top_bl2[3] array_top_bl2_n[3] bl1 bl1_n bl2 bl2_n array_top_bl1[5] array_top_bl1_n[5] array_top_bl2[5] array_top_bl2_n[5] array_top_bl1[6] array_top_bl1_n[6] array_top_bl2[6] array_top_bl2_n[6] array_top_bl1[7] array_top_bl1_n[7] array_top_bl2[7] array_top_bl2_n[7] DP8TVar6Array_6X8
Xzero vdd vss zero zero_x1
.ends DP8TVar6TestArray_16X8C

.subckt PadFrame_DP06 PAD0x0 PAD0x1 PAD0x2 PAD0x3 PAD0x4 PAD0x5 PAD0x6 PAD0x7 PAD0x8 PAD0x9 PAD1x0 PAD1x1 PAD1x2 PAD1x3 PAD1x4 PAD1x5 PAD1x6 PAD1x7 PAD1x8 PAD1x9
XPAD0x0 PAD0x0 BondPad
XPAD0x1 PAD0x1 BondPad
XPAD0x2 PAD0x2 BondPad
XPAD0x3 PAD0x3 BondPad
XPAD0x4 PAD0x4 BondPad
XPAD0x5 PAD0x5 BondPad
XPAD0x6 PAD0x6 BondPad
XPAD0x7 PAD0x7 BondPad
XPAD0x8 PAD0x8 BondPad
XPAD0x9 PAD0x9 BondPad
XPAD1x0 PAD1x0 BondPad
XPAD1x1 PAD1x1 BondPad
XPAD1x2 PAD1x2 BondPad
XPAD1x3 PAD1x3 BondPad
XPAD1x4 PAD1x4 BondPad
XPAD1x5 PAD1x5 BondPad
XPAD1x6 PAD1x6 BondPad
XPAD1x7 PAD1x7 BondPad
XPAD1x8 PAD1x8 BondPad
XPAD1x9 PAD1x9 BondPad
.ends PadFrame_DP06

.subckt DP8TVar6 vss noco_vdd noco_wl1 noco_wl2 noco_bl1 noco_bl1_n noco_bl2 noco_bl2_n co_vdd co_bit co_bit_n co_wl1 co_wl2 co_bl1 co_bl1_n co_bl2_n co_bl2
Xframe noco_vdd noco_wl1 noco_wl2 noco_bl2 co_vdd co_bit co_bit_n co_wl1 co_wl2 NoConn_PAD0x9 vss noco_bl1 noco_bl1_n noco_bl2_n vss co_bl1 co_bl1_n co_bl2_n co_bl2 NoConn_PAD1x9 PadFrame_DP06
Xtestarray_noco vss noco_vdd noco_wl1 noco_wl2 noco_bl1 noco_bl1_n noco_bl2 noco_bl2_n DP8TVar6TestArray_16X8
Xtestarray_co vss co_vdd co_wl1 co_wl2 co_bl1 co_bl1_n co_bl2 co_bl2_n co_bit co_bit_n DP8TVar6TestArray_16X8C
.ends DP8TVar6

.subckt PadFrame_SP22 PAD0x0 PAD0x1 PAD0x2 PAD0x3 PAD0x4 PAD0x5 PAD0x6 PAD0x7 PAD0x8 PAD0x9 PAD1x0 PAD1x1 PAD1x2 PAD1x3 PAD1x4 PAD1x5 PAD1x6 PAD1x7 PAD1x8 PAD1x9
XPAD0x0 PAD0x0 BondPad
XPAD0x1 PAD0x1 BondPad
XPAD0x2 PAD0x2 BondPad
XPAD0x3 PAD0x3 BondPad
XPAD0x4 PAD0x4 BondPad
XPAD0x5 PAD0x5 BondPad
XPAD0x6 PAD0x6 BondPad
XPAD0x7 PAD0x7 BondPad
XPAD0x8 PAD0x8 BondPad
XPAD0x9 PAD0x9 BondPad
XPAD1x0 PAD1x0 BondPad
XPAD1x1 PAD1x1 BondPad
XPAD1x2 PAD1x2 BondPad
XPAD1x3 PAD1x3 BondPad
XPAD1x4 PAD1x4 BondPad
XPAD1x5 PAD1x5 BondPad
XPAD1x6 PAD1x6 BondPad
XPAD1x7 PAD1x7 BondPad
XPAD1x8 PAD1x8 BondPad
XPAD1x9 PAD1x9 BondPad
.ends PadFrame_SP22

.subckt SP6TVar22Cell wl bl bl_n vdd vss
Xpu1 vdd bit_n bit vdd sg13_lv_pmos l=1.3e-07 w=3e-07
Xpd1 bit bit_n vss vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpu2 vdd bit bit_n vdd sg13_lv_pmos l=1.3e-07 w=3e-07
Xpd2 bit_n bit vss vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg1 bit wl bl vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg2 bit_n wl bl_n vss sg13_lv_nmos l=1.3e-07 w=3e-07
.ends SP6TVar22Cell

.subckt SP6TVar22Array_2X1 vss vdd wl[0] wl[1] bl[0] bl_n[0]
Xinst0x0 wl[0] bl[0] bl_n[0] vdd vss SP6TVar22Cell
Xinst1x0 wl[1] bl[0] bl_n[0] vdd vss SP6TVar22Cell
.ends SP6TVar22Array_2X1

.subckt SP6TVar22Array_2X2 vss vdd wl[0] wl[1] bl[0] bl_n[0] bl[1] bl_n[1]
Xinst0x0 vss vdd wl[0] wl[1] bl[0] bl_n[0] SP6TVar22Array_2X1
Xinst0x1 vss vdd wl[0] wl[1] bl[1] bl_n[1] SP6TVar22Array_2X1
.ends SP6TVar22Array_2X2

.subckt SP6TVar22Array_4X2 vss vdd wl[0] wl[1] wl[2] wl[3] bl[0] bl_n[0] bl[1] bl_n[1]
Xinst0x0 vss vdd wl[0] wl[1] bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar22Array_2X2
Xinst1x0 vss vdd wl[2] wl[3] bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar22Array_2X2
.ends SP6TVar22Array_4X2

.subckt SP6TVar22Array_4X4 vss vdd wl[0] wl[1] wl[2] wl[3] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar22Array_4X2
Xinst0x1 vss vdd wl[0] wl[1] wl[2] wl[3] bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar22Array_4X2
.ends SP6TVar22Array_4X4

.subckt SP6TVar22Array_8X4 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar22Array_4X4
Xinst1x0 vss vdd wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar22Array_4X4
.ends SP6TVar22Array_8X4

.subckt SP6TVar22Array_8X8 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar22Array_8X4
Xinst0x1 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7] SP6TVar22Array_8X4
.ends SP6TVar22Array_8X8

.subckt SP6TVar22Array_8X16 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7] bl[8] bl_n[8] bl[9] bl_n[9] bl[10] bl_n[10] bl[11] bl_n[11] bl[12] bl_n[12] bl[13] bl_n[13] bl[14] bl_n[14] bl[15] bl_n[15]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7] SP6TVar22Array_8X8
Xinst0x1 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[8] bl_n[8] bl[9] bl_n[9] bl[10] bl_n[10] bl[11] bl_n[11] bl[12] bl_n[12] bl[13] bl_n[13] bl[14] bl_n[14] bl[15] bl_n[15] SP6TVar22Array_8X8
.ends SP6TVar22Array_8X16

.subckt SP6TVar22TestArray_8X16 vss vdd bl bl_n wl
Xarray vss vdd zero zero zero zero wl zero zero zero bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7] bl bl_n bl[9] bl_n[9] bl[10] bl_n[10] bl[11] bl_n[11] bl[12] bl_n[12] bl[13] bl_n[13] bl[14] bl_n[14] bl[15] bl_n[15] SP6TVar22Array_8X16
Xzero vdd vss zero zero_x1
.ends SP6TVar22TestArray_8X16

.subckt SP6TVar22Array_4X1 vss vdd wl[0] wl[1] wl[2] wl[3] bl[0] bl_n[0]
Xinst0x0 vss vdd wl[0] wl[1] bl[0] bl_n[0] SP6TVar22Array_2X1
Xinst1x0 vss vdd wl[2] wl[3] bl[0] bl_n[0] SP6TVar22Array_2X1
.ends SP6TVar22Array_4X1

.subckt SP6TVar22Array_8X1 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] bl[0] bl_n[0] SP6TVar22Array_4X1
Xinst1x0 vss vdd wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] SP6TVar22Array_4X1
.ends SP6TVar22Array_8X1

.subckt SP6TVar22Array_8X2 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar22Array_4X2
Xinst1x0 vss vdd wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar22Array_4X2
.ends SP6TVar22Array_8X2

.subckt SP6TVar22CellConnectOut wl bl bl_n vdd vss bit bit_n
Xpu1 vdd bit_n bit vdd sg13_lv_pmos l=1.3e-07 w=3e-07
Xpd1 bit bit_n vss vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpu2 vdd bit bit_n vdd sg13_lv_pmos l=1.3e-07 w=3e-07
Xpd2 bit_n bit vss vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg1 bit wl bl vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg2 bit_n wl bl_n vss sg13_lv_nmos l=1.3e-07 w=3e-07
.ends SP6TVar22CellConnectOut

.subckt SP6TVar22TestArray_8X16C vss vdd bl bl_n bit bit_n wl
Xarray_0 vss vdd zero zero zero zero wl zero zero zero array_0_bl[0] array_0_bl_n[0] SP6TVar22Array_8X1
Xarray_1 vss vdd zero zero zero zero wl zero zero zero array_1_bl[0] array_1_bl_n[0] array_1_bl[1] array_1_bl_n[1] SP6TVar22Array_8X2
Xarray_2 vss vdd zero zero zero zero wl zero zero zero array_2_bl[0] array_2_bl_n[0] array_2_bl[1] array_2_bl_n[1] array_2_bl[2] array_2_bl_n[2] array_2_bl[3] array_2_bl_n[3] SP6TVar22Array_8X4
Xarray_3 vss vdd zero zero zero zero wl zero zero zero array_3_bl[0] array_3_bl_n[0] array_3_bl[1] array_3_bl_n[1] array_3_bl[2] array_3_bl_n[2] array_3_bl[3] array_3_bl_n[3] array_3_bl[4] array_3_bl_n[4] array_3_bl[5] array_3_bl_n[5] array_3_bl[6] array_3_bl_n[6] array_3_bl[7] array_3_bl_n[7] SP6TVar22Array_8X8
Xcolarray_0 vss vdd zero zero zero zero bl bl_n SP6TVar22Array_4X1
Xcolarray_1 vss vdd zero zero bl bl_n SP6TVar22Array_2X1
Xbc_noconn zero bl bl_n vdd vss SP6TVar22Cell
Xbc_conn wl bl bl_n vdd vss bit bit_n SP6TVar22CellConnectOut
Xzero vdd vss zero zero_x1
.ends SP6TVar22TestArray_8X16C

.subckt SP6TVar22 vss noco_vdd noco_wl noco_bl noco_bl_n co_vdd co_bl co_bl_n co_bit co_bit_n co_wl
Xframe noco_vdd noco_wl NoConn_PAD0x2 co_vdd co_bl_n co_bit co_bit_n NoConn_PAD0x7 NoConn_PAD0x8 NoConn_PAD0x9 vss noco_bl noco_bl_n vss co_bl co_wl NoConn_PAD1x6 NoConn_PAD1x7 NoConn_PAD1x8 NoConn_PAD1x9 PadFrame_SP22
Xtestarray_noco vss noco_vdd noco_bl noco_bl_n noco_wl SP6TVar22TestArray_8X16
Xtestarray_co vss co_vdd co_bl co_bl_n co_bit co_bit_n co_wl SP6TVar22TestArray_8X16C
.ends SP6TVar22

.subckt PadFrame_SP07 PAD0x0 PAD0x1 PAD0x2 PAD0x3 PAD0x4 PAD0x5 PAD0x6 PAD0x7 PAD0x8 PAD0x9 PAD1x0 PAD1x1 PAD1x2 PAD1x3 PAD1x4 PAD1x5 PAD1x6 PAD1x7 PAD1x8 PAD1x9
XPAD0x0 PAD0x0 BondPad
XPAD0x1 PAD0x1 BondPad
XPAD0x2 PAD0x2 BondPad
XPAD0x3 PAD0x3 BondPad
XPAD0x4 PAD0x4 BondPad
XPAD0x5 PAD0x5 BondPad
XPAD0x6 PAD0x6 BondPad
XPAD0x7 PAD0x7 BondPad
XPAD0x8 PAD0x8 BondPad
XPAD0x9 PAD0x9 BondPad
XPAD1x0 PAD1x0 BondPad
XPAD1x1 PAD1x1 BondPad
XPAD1x2 PAD1x2 BondPad
XPAD1x3 PAD1x3 BondPad
XPAD1x4 PAD1x4 BondPad
XPAD1x5 PAD1x5 BondPad
XPAD1x6 PAD1x6 BondPad
XPAD1x7 PAD1x7 BondPad
XPAD1x8 PAD1x8 BondPad
XPAD1x9 PAD1x9 BondPad
.ends PadFrame_SP07

.subckt SP6TVar7Cell wl bl bl_n vdd vss
Xpu1 vdd bit_n bit vdd sg13_lv_pmos l=1.3e-07 w=3e-07
Xpd1 bit bit_n vss vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpu2 vdd bit bit_n vdd sg13_lv_pmos l=1.3e-07 w=3e-07
Xpd2 bit_n bit vss vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg1 bit wl bl vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg2 bit_n wl bl_n vss sg13_lv_nmos l=1.3e-07 w=3e-07
.ends SP6TVar7Cell

.subckt SP6TVar7Array_2X1 vss vdd wl[0] wl[1] bl[0] bl_n[0]
Xinst0x0 wl[0] bl[0] bl_n[0] vdd vss SP6TVar7Cell
Xinst1x0 wl[1] bl[0] bl_n[0] vdd vss SP6TVar7Cell
.ends SP6TVar7Array_2X1

.subckt SP6TVar7Array_2X2 vss vdd wl[0] wl[1] bl[0] bl_n[0] bl[1] bl_n[1]
Xinst0x0 vss vdd wl[0] wl[1] bl[0] bl_n[0] SP6TVar7Array_2X1
Xinst0x1 vss vdd wl[0] wl[1] bl[1] bl_n[1] SP6TVar7Array_2X1
.ends SP6TVar7Array_2X2

.subckt SP6TVar7Array_4X2 vss vdd wl[0] wl[1] wl[2] wl[3] bl[0] bl_n[0] bl[1] bl_n[1]
Xinst0x0 vss vdd wl[0] wl[1] bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar7Array_2X2
Xinst1x0 vss vdd wl[2] wl[3] bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar7Array_2X2
.ends SP6TVar7Array_4X2

.subckt SP6TVar7Array_4X4 vss vdd wl[0] wl[1] wl[2] wl[3] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar7Array_4X2
Xinst0x1 vss vdd wl[0] wl[1] wl[2] wl[3] bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar7Array_4X2
.ends SP6TVar7Array_4X4

.subckt SP6TVar7Array_8X4 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar7Array_4X4
Xinst1x0 vss vdd wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar7Array_4X4
.ends SP6TVar7Array_8X4

.subckt SP6TVar7Array_8X8 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar7Array_8X4
Xinst0x1 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7] SP6TVar7Array_8X4
.ends SP6TVar7Array_8X8

.subckt SP6TVar7BulkConn vdd vss bl bl_n
.ends SP6TVar7BulkConn

.subckt SP6TVar7BulkConnRow_2 vss vdd bl[0] bl_n[0] bl[1] bl_n[1]
Xinst0 vdd vss bl[0] bl_n[0] SP6TVar7BulkConn
Xinst1 vdd vss bl[1] bl_n[1] SP6TVar7BulkConn
.ends SP6TVar7BulkConnRow_2

.subckt SP6TVar7BulkConnRow_4 vss vdd bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3]
Xinst0 vss vdd bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar7BulkConnRow_2
Xinst1 vss vdd bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar7BulkConnRow_2
.ends SP6TVar7BulkConnRow_4

.subckt SP6TVar7BulkConnRow_8 vss vdd bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7]
Xinst0 vss vdd bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar7BulkConnRow_4
Xinst1 vss vdd bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7] SP6TVar7BulkConnRow_4
.ends SP6TVar7BulkConnRow_8

.subckt SP6TVar7Array_16X8BC vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7] SP6TVar7Array_8X8
Xinst1x0 vss vdd wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7] SP6TVar7Array_8X8
Xbottombcrow vss vdd bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7] SP6TVar7BulkConnRow_8
Xtopbcrow vss vdd bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7] SP6TVar7BulkConnRow_8
.ends SP6TVar7Array_16X8BC

.subckt SP6TVar7TestArray_16X8 vss vdd bl bl_n wl
Xarray vss vdd zero zero zero zero zero zero zero zero wl zero zero zero zero zero zero zero bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl bl_n bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7] SP6TVar7Array_16X8BC
Xzero vdd vss zero zero_x1
.ends SP6TVar7TestArray_16X8

.subckt SP6TVar7Array_4X1 vss vdd wl[0] wl[1] wl[2] wl[3] bl[0] bl_n[0]
Xinst0x0 vss vdd wl[0] wl[1] bl[0] bl_n[0] SP6TVar7Array_2X1
Xinst1x0 vss vdd wl[2] wl[3] bl[0] bl_n[0] SP6TVar7Array_2X1
.ends SP6TVar7Array_4X1

.subckt SP6TVar7Array_8X1 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] bl[0] bl_n[0] SP6TVar7Array_4X1
Xinst1x0 vss vdd wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] SP6TVar7Array_4X1
.ends SP6TVar7Array_8X1

.subckt SP6TVar7Array_16X1BC vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] bl[0] bl_n[0]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] SP6TVar7Array_8X1
Xinst1x0 vss vdd wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] bl[0] bl_n[0] SP6TVar7Array_8X1
Xbottombcrow vdd vss bl[0] bl_n[0] SP6TVar7BulkConn
Xtopbcrow vdd vss bl[0] bl_n[0] SP6TVar7BulkConn
.ends SP6TVar7Array_16X1BC

.subckt SP6TVar7Array_8X2 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar7Array_4X2
Xinst1x0 vss vdd wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar7Array_4X2
.ends SP6TVar7Array_8X2

.subckt SP6TVar7Array_16X2BC vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] bl[0] bl_n[0] bl[1] bl_n[1]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar7Array_8X2
Xinst1x0 vss vdd wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar7Array_8X2
Xbottombcrow vss vdd bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar7BulkConnRow_2
Xtopbcrow vss vdd bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar7BulkConnRow_2
.ends SP6TVar7Array_16X2BC

.subckt SP6TVar7Array_16X4BC vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar7Array_8X4
Xinst1x0 vss vdd wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar7Array_8X4
Xbottombcrow vss vdd bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar7BulkConnRow_4
Xtopbcrow vss vdd bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar7BulkConnRow_4
.ends SP6TVar7Array_16X4BC

.subckt SP6TVar7Array_6X1 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] bl[0] bl_n[0]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] bl[0] bl_n[0] SP6TVar7Array_4X1
Xinst1x0 vss vdd wl[4] wl[5] bl[0] bl_n[0] SP6TVar7Array_2X1
.ends SP6TVar7Array_6X1

.subckt SP6TVar7CellConnectOut wl bl bl_n vdd vss bit bit_n
Xpu1 vdd bit_n bit vdd sg13_lv_pmos l=1.3e-07 w=3e-07
Xpd1 bit bit_n vss vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpu2 vdd bit bit_n vdd sg13_lv_pmos l=1.3e-07 w=3e-07
Xpd2 bit_n bit vss vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg1 bit wl bl vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg2 bit_n wl bl_n vss sg13_lv_nmos l=1.3e-07 w=3e-07
.ends SP6TVar7CellConnectOut

.subckt SP6TVar7TestArray_16X8C vss vdd bl bl_n bit bit_n wl
Xarray_0 vss vdd zero zero zero zero zero zero zero zero wl zero zero zero zero zero zero zero array_0_bl[0] array_0_bl_n[0] SP6TVar7Array_16X1BC
Xarray_1 vss vdd zero zero zero zero zero zero zero zero wl zero zero zero zero zero zero zero array_1_bl[0] array_1_bl_n[0] array_1_bl[1] array_1_bl_n[1] SP6TVar7Array_16X2BC
Xarray_2 vss vdd zero zero zero zero zero zero zero zero wl zero zero zero zero zero zero zero array_2_bl[0] array_2_bl_n[0] array_2_bl[1] array_2_bl_n[1] array_2_bl[2] array_2_bl_n[2] array_2_bl[3] array_2_bl_n[3] SP6TVar7Array_16X4BC
Xcolbc_0 vdd vss bl bl_n SP6TVar7BulkConn
Xcolbc_1 vdd vss bl bl_n SP6TVar7BulkConn
Xcolarray_0 vss vdd zero zero zero zero zero zero zero zero bl bl_n SP6TVar7Array_8X1
Xcolarray_1 vss vdd zero zero zero zero zero zero bl bl_n SP6TVar7Array_6X1
Xbc_noconn zero bl bl_n vdd vss SP6TVar7Cell
Xbc_conn wl bl bl_n vdd vss bit bit_n SP6TVar7CellConnectOut
Xzero vdd vss zero zero_x1
.ends SP6TVar7TestArray_16X8C

.subckt SP6TVar7 vss noco_vdd noco_wl noco_bl noco_bl_n co_vdd co_bl co_bl_n co_bit co_bit_n co_wl
Xframe noco_vdd noco_wl NoConn_PAD0x2 co_vdd co_bl_n co_bit co_bit_n NoConn_PAD0x7 NoConn_PAD0x8 NoConn_PAD0x9 vss noco_bl noco_bl_n vss co_bl co_wl NoConn_PAD1x6 NoConn_PAD1x7 NoConn_PAD1x8 NoConn_PAD1x9 PadFrame_SP07
Xtestarray_noco vss noco_vdd noco_bl noco_bl_n noco_wl SP6TVar7TestArray_16X8
Xtestarray_co vss co_vdd co_bl co_bl_n co_bit co_bit_n co_wl SP6TVar7TestArray_16X8C
.ends SP6TVar7

.subckt PadFrame_SP08 PAD0x0 PAD0x1 PAD0x2 PAD0x3 PAD0x4 PAD0x5 PAD0x6 PAD0x7 PAD0x8 PAD0x9 PAD1x0 PAD1x1 PAD1x2 PAD1x3 PAD1x4 PAD1x5 PAD1x6 PAD1x7 PAD1x8 PAD1x9
XPAD0x0 PAD0x0 BondPad
XPAD0x1 PAD0x1 BondPad
XPAD0x2 PAD0x2 BondPad
XPAD0x3 PAD0x3 BondPad
XPAD0x4 PAD0x4 BondPad
XPAD0x5 PAD0x5 BondPad
XPAD0x6 PAD0x6 BondPad
XPAD0x7 PAD0x7 BondPad
XPAD0x8 PAD0x8 BondPad
XPAD0x9 PAD0x9 BondPad
XPAD1x0 PAD1x0 BondPad
XPAD1x1 PAD1x1 BondPad
XPAD1x2 PAD1x2 BondPad
XPAD1x3 PAD1x3 BondPad
XPAD1x4 PAD1x4 BondPad
XPAD1x5 PAD1x5 BondPad
XPAD1x6 PAD1x6 BondPad
XPAD1x7 PAD1x7 BondPad
XPAD1x8 PAD1x8 BondPad
XPAD1x9 PAD1x9 BondPad
.ends PadFrame_SP08

.subckt SP6TVar8Cell wl bl bl_n vdd vss
Xpu1 vdd bit_n bit vdd sg13_lv_pmos l=1.3e-07 w=2e-07
Xpd1 bit bit_n vss vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpu2 vdd bit bit_n vdd sg13_lv_pmos l=1.3e-07 w=2e-07
Xpd2 bit_n bit vss vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg1 bit wl bl vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg2 bit_n wl bl_n vss sg13_lv_nmos l=1.3e-07 w=3e-07
.ends SP6TVar8Cell

.subckt SP6TVar8Array_2X1 vss vdd wl[0] wl[1] bl[0] bl_n[0]
Xinst0x0 wl[0] bl[0] bl_n[0] vdd vss SP6TVar8Cell
Xinst1x0 wl[1] bl[0] bl_n[0] vdd vss SP6TVar8Cell
.ends SP6TVar8Array_2X1

.subckt SP6TVar8Array_2X2 vss vdd wl[0] wl[1] bl[0] bl_n[0] bl[1] bl_n[1]
Xinst0x0 vss vdd wl[0] wl[1] bl[0] bl_n[0] SP6TVar8Array_2X1
Xinst0x1 vss vdd wl[0] wl[1] bl[1] bl_n[1] SP6TVar8Array_2X1
.ends SP6TVar8Array_2X2

.subckt SP6TVar8Array_4X2 vss vdd wl[0] wl[1] wl[2] wl[3] bl[0] bl_n[0] bl[1] bl_n[1]
Xinst0x0 vss vdd wl[0] wl[1] bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar8Array_2X2
Xinst1x0 vss vdd wl[2] wl[3] bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar8Array_2X2
.ends SP6TVar8Array_4X2

.subckt SP6TVar8Array_4X4 vss vdd wl[0] wl[1] wl[2] wl[3] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar8Array_4X2
Xinst0x1 vss vdd wl[0] wl[1] wl[2] wl[3] bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar8Array_4X2
.ends SP6TVar8Array_4X4

.subckt SP6TVar8Array_8X4 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar8Array_4X4
Xinst1x0 vss vdd wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar8Array_4X4
.ends SP6TVar8Array_8X4

.subckt SP6TVar8Array_8X8 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar8Array_8X4
Xinst0x1 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7] SP6TVar8Array_8X4
.ends SP6TVar8Array_8X8

.subckt SP6TVar8BulkConn vdd vss bl bl_n
.ends SP6TVar8BulkConn

.subckt SP6TVar8BulkConnRow_2 vss vdd bl[0] bl_n[0] bl[1] bl_n[1]
Xinst0 vdd vss bl[0] bl_n[0] SP6TVar8BulkConn
Xinst1 vdd vss bl[1] bl_n[1] SP6TVar8BulkConn
.ends SP6TVar8BulkConnRow_2

.subckt SP6TVar8BulkConnRow_4 vss vdd bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3]
Xinst0 vss vdd bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar8BulkConnRow_2
Xinst1 vss vdd bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar8BulkConnRow_2
.ends SP6TVar8BulkConnRow_4

.subckt SP6TVar8BulkConnRow_8 vss vdd bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7]
Xinst0 vss vdd bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar8BulkConnRow_4
Xinst1 vss vdd bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7] SP6TVar8BulkConnRow_4
.ends SP6TVar8BulkConnRow_8

.subckt SP6TVar8Array_16X8BC vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7] SP6TVar8Array_8X8
Xinst1x0 vss vdd wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7] SP6TVar8Array_8X8
Xbottombcrow vss vdd bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7] SP6TVar8BulkConnRow_8
Xtopbcrow vss vdd bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7] SP6TVar8BulkConnRow_8
.ends SP6TVar8Array_16X8BC

.subckt SP6TVar8TestArray_16X8 vss vdd bl bl_n wl
Xarray vss vdd zero zero zero zero zero zero zero zero wl zero zero zero zero zero zero zero bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl bl_n bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7] SP6TVar8Array_16X8BC
Xzero vdd vss zero zero_x1
.ends SP6TVar8TestArray_16X8

.subckt SP6TVar8Array_4X1 vss vdd wl[0] wl[1] wl[2] wl[3] bl[0] bl_n[0]
Xinst0x0 vss vdd wl[0] wl[1] bl[0] bl_n[0] SP6TVar8Array_2X1
Xinst1x0 vss vdd wl[2] wl[3] bl[0] bl_n[0] SP6TVar8Array_2X1
.ends SP6TVar8Array_4X1

.subckt SP6TVar8Array_8X1 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] bl[0] bl_n[0] SP6TVar8Array_4X1
Xinst1x0 vss vdd wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] SP6TVar8Array_4X1
.ends SP6TVar8Array_8X1

.subckt SP6TVar8Array_16X1BC vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] bl[0] bl_n[0]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] SP6TVar8Array_8X1
Xinst1x0 vss vdd wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] bl[0] bl_n[0] SP6TVar8Array_8X1
Xbottombcrow vdd vss bl[0] bl_n[0] SP6TVar8BulkConn
Xtopbcrow vdd vss bl[0] bl_n[0] SP6TVar8BulkConn
.ends SP6TVar8Array_16X1BC

.subckt SP6TVar8Array_8X2 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar8Array_4X2
Xinst1x0 vss vdd wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar8Array_4X2
.ends SP6TVar8Array_8X2

.subckt SP6TVar8Array_16X2BC vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] bl[0] bl_n[0] bl[1] bl_n[1]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar8Array_8X2
Xinst1x0 vss vdd wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar8Array_8X2
Xbottombcrow vss vdd bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar8BulkConnRow_2
Xtopbcrow vss vdd bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar8BulkConnRow_2
.ends SP6TVar8Array_16X2BC

.subckt SP6TVar8Array_16X4BC vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar8Array_8X4
Xinst1x0 vss vdd wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar8Array_8X4
Xbottombcrow vss vdd bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar8BulkConnRow_4
Xtopbcrow vss vdd bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar8BulkConnRow_4
.ends SP6TVar8Array_16X4BC

.subckt SP6TVar8Array_6X1 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] bl[0] bl_n[0]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] bl[0] bl_n[0] SP6TVar8Array_4X1
Xinst1x0 vss vdd wl[4] wl[5] bl[0] bl_n[0] SP6TVar8Array_2X1
.ends SP6TVar8Array_6X1

.subckt SP6TVar8CellConnectOut wl bl bl_n vdd vss bit bit_n
Xpu1 vdd bit_n bit vdd sg13_lv_pmos l=1.3e-07 w=2e-07
Xpd1 bit bit_n vss vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpu2 vdd bit bit_n vdd sg13_lv_pmos l=1.3e-07 w=2e-07
Xpd2 bit_n bit vss vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg1 bit wl bl vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg2 bit_n wl bl_n vss sg13_lv_nmos l=1.3e-07 w=3e-07
.ends SP6TVar8CellConnectOut

.subckt SP6TVar8TestArray_16X8C vss vdd bl bl_n bit bit_n wl
Xarray_0 vss vdd zero zero zero zero zero zero zero zero wl zero zero zero zero zero zero zero array_0_bl[0] array_0_bl_n[0] SP6TVar8Array_16X1BC
Xarray_1 vss vdd zero zero zero zero zero zero zero zero wl zero zero zero zero zero zero zero array_1_bl[0] array_1_bl_n[0] array_1_bl[1] array_1_bl_n[1] SP6TVar8Array_16X2BC
Xarray_2 vss vdd zero zero zero zero zero zero zero zero wl zero zero zero zero zero zero zero array_2_bl[0] array_2_bl_n[0] array_2_bl[1] array_2_bl_n[1] array_2_bl[2] array_2_bl_n[2] array_2_bl[3] array_2_bl_n[3] SP6TVar8Array_16X4BC
Xcolbc_0 vdd vss bl bl_n SP6TVar8BulkConn
Xcolbc_1 vdd vss bl bl_n SP6TVar8BulkConn
Xcolarray_0 vss vdd zero zero zero zero zero zero zero zero bl bl_n SP6TVar8Array_8X1
Xcolarray_1 vss vdd zero zero zero zero zero zero bl bl_n SP6TVar8Array_6X1
Xbc_noconn zero bl bl_n vdd vss SP6TVar8Cell
Xbc_conn wl bl bl_n vdd vss bit bit_n SP6TVar8CellConnectOut
Xzero vdd vss zero zero_x1
.ends SP6TVar8TestArray_16X8C

.subckt SP6TVar8 vss noco_vdd noco_wl noco_bl noco_bl_n co_vdd co_bl co_bl_n co_bit co_bit_n co_wl
Xframe noco_vdd noco_wl NoConn_PAD0x2 co_vdd co_bl_n co_bit co_bit_n NoConn_PAD0x7 NoConn_PAD0x8 NoConn_PAD0x9 vss noco_bl noco_bl_n vss co_bl co_wl NoConn_PAD1x6 NoConn_PAD1x7 NoConn_PAD1x8 NoConn_PAD1x9 PadFrame_SP08
Xtestarray_noco vss noco_vdd noco_bl noco_bl_n noco_wl SP6TVar8TestArray_16X8
Xtestarray_co vss co_vdd co_bl co_bl_n co_bit co_bit_n co_wl SP6TVar8TestArray_16X8C
.ends SP6TVar8

.subckt PadFrame_SP09 PAD0x0 PAD0x1 PAD0x2 PAD0x3 PAD0x4 PAD0x5 PAD0x6 PAD0x7 PAD0x8 PAD0x9 PAD1x0 PAD1x1 PAD1x2 PAD1x3 PAD1x4 PAD1x5 PAD1x6 PAD1x7 PAD1x8 PAD1x9
XPAD0x0 PAD0x0 BondPad
XPAD0x1 PAD0x1 BondPad
XPAD0x2 PAD0x2 BondPad
XPAD0x3 PAD0x3 BondPad
XPAD0x4 PAD0x4 BondPad
XPAD0x5 PAD0x5 BondPad
XPAD0x6 PAD0x6 BondPad
XPAD0x7 PAD0x7 BondPad
XPAD0x8 PAD0x8 BondPad
XPAD0x9 PAD0x9 BondPad
XPAD1x0 PAD1x0 BondPad
XPAD1x1 PAD1x1 BondPad
XPAD1x2 PAD1x2 BondPad
XPAD1x3 PAD1x3 BondPad
XPAD1x4 PAD1x4 BondPad
XPAD1x5 PAD1x5 BondPad
XPAD1x6 PAD1x6 BondPad
XPAD1x7 PAD1x7 BondPad
XPAD1x8 PAD1x8 BondPad
XPAD1x9 PAD1x9 BondPad
.ends PadFrame_SP09

.subckt SP6TVar9Cell wl bl bl_n vdd vss
Xpu1 vdd bit_n bit vdd sg13_lv_pmos l=1.3e-07 w=1.5e-07
Xpd1 bit bit_n vss vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpu2 vdd bit bit_n vdd sg13_lv_pmos l=1.3e-07 w=1.5e-07
Xpd2 bit_n bit vss vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg1 bit wl bl vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg2 bit_n wl bl_n vss sg13_lv_nmos l=1.3e-07 w=3e-07
.ends SP6TVar9Cell

.subckt SP6TVar9Array_2X1 vss vdd wl[0] wl[1] bl[0] bl_n[0]
Xinst0x0 wl[0] bl[0] bl_n[0] vdd vss SP6TVar9Cell
Xinst1x0 wl[1] bl[0] bl_n[0] vdd vss SP6TVar9Cell
.ends SP6TVar9Array_2X1

.subckt SP6TVar9Array_2X2 vss vdd wl[0] wl[1] bl[0] bl_n[0] bl[1] bl_n[1]
Xinst0x0 vss vdd wl[0] wl[1] bl[0] bl_n[0] SP6TVar9Array_2X1
Xinst0x1 vss vdd wl[0] wl[1] bl[1] bl_n[1] SP6TVar9Array_2X1
.ends SP6TVar9Array_2X2

.subckt SP6TVar9Array_4X2 vss vdd wl[0] wl[1] wl[2] wl[3] bl[0] bl_n[0] bl[1] bl_n[1]
Xinst0x0 vss vdd wl[0] wl[1] bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar9Array_2X2
Xinst1x0 vss vdd wl[2] wl[3] bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar9Array_2X2
.ends SP6TVar9Array_4X2

.subckt SP6TVar9Array_4X4 vss vdd wl[0] wl[1] wl[2] wl[3] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar9Array_4X2
Xinst0x1 vss vdd wl[0] wl[1] wl[2] wl[3] bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar9Array_4X2
.ends SP6TVar9Array_4X4

.subckt SP6TVar9Array_8X4 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar9Array_4X4
Xinst1x0 vss vdd wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar9Array_4X4
.ends SP6TVar9Array_8X4

.subckt SP6TVar9Array_8X8 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar9Array_8X4
Xinst0x1 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7] SP6TVar9Array_8X4
.ends SP6TVar9Array_8X8

.subckt SP6TVar9BulkConn vdd vss bl bl_n
.ends SP6TVar9BulkConn

.subckt SP6TVar9BulkConnRow_2 vss vdd bl[0] bl_n[0] bl[1] bl_n[1]
Xinst0 vdd vss bl[0] bl_n[0] SP6TVar9BulkConn
Xinst1 vdd vss bl[1] bl_n[1] SP6TVar9BulkConn
.ends SP6TVar9BulkConnRow_2

.subckt SP6TVar9BulkConnRow_4 vss vdd bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3]
Xinst0 vss vdd bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar9BulkConnRow_2
Xinst1 vss vdd bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar9BulkConnRow_2
.ends SP6TVar9BulkConnRow_4

.subckt SP6TVar9BulkConnRow_8 vss vdd bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7]
Xinst0 vss vdd bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar9BulkConnRow_4
Xinst1 vss vdd bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7] SP6TVar9BulkConnRow_4
.ends SP6TVar9BulkConnRow_8

.subckt SP6TVar9Array_16X8BC vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7] SP6TVar9Array_8X8
Xinst1x0 vss vdd wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7] SP6TVar9Array_8X8
Xbottombcrow vss vdd bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7] SP6TVar9BulkConnRow_8
Xtopbcrow vss vdd bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7] SP6TVar9BulkConnRow_8
.ends SP6TVar9Array_16X8BC

.subckt SP6TVar9TestArray_16X8 vss vdd bl bl_n wl
Xarray vss vdd zero zero zero zero zero zero zero zero wl zero zero zero zero zero zero zero bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl bl_n bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7] SP6TVar9Array_16X8BC
Xzero vdd vss zero zero_x1
.ends SP6TVar9TestArray_16X8

.subckt SP6TVar9Array_4X1 vss vdd wl[0] wl[1] wl[2] wl[3] bl[0] bl_n[0]
Xinst0x0 vss vdd wl[0] wl[1] bl[0] bl_n[0] SP6TVar9Array_2X1
Xinst1x0 vss vdd wl[2] wl[3] bl[0] bl_n[0] SP6TVar9Array_2X1
.ends SP6TVar9Array_4X1

.subckt SP6TVar9Array_8X1 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] bl[0] bl_n[0] SP6TVar9Array_4X1
Xinst1x0 vss vdd wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] SP6TVar9Array_4X1
.ends SP6TVar9Array_8X1

.subckt SP6TVar9Array_16X1BC vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] bl[0] bl_n[0]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] SP6TVar9Array_8X1
Xinst1x0 vss vdd wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] bl[0] bl_n[0] SP6TVar9Array_8X1
Xbottombcrow vdd vss bl[0] bl_n[0] SP6TVar9BulkConn
Xtopbcrow vdd vss bl[0] bl_n[0] SP6TVar9BulkConn
.ends SP6TVar9Array_16X1BC

.subckt SP6TVar9Array_8X2 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar9Array_4X2
Xinst1x0 vss vdd wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar9Array_4X2
.ends SP6TVar9Array_8X2

.subckt SP6TVar9Array_16X2BC vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] bl[0] bl_n[0] bl[1] bl_n[1]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar9Array_8X2
Xinst1x0 vss vdd wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar9Array_8X2
Xbottombcrow vss vdd bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar9BulkConnRow_2
Xtopbcrow vss vdd bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar9BulkConnRow_2
.ends SP6TVar9Array_16X2BC

.subckt SP6TVar9Array_16X4BC vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar9Array_8X4
Xinst1x0 vss vdd wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar9Array_8X4
Xbottombcrow vss vdd bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar9BulkConnRow_4
Xtopbcrow vss vdd bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar9BulkConnRow_4
.ends SP6TVar9Array_16X4BC

.subckt SP6TVar9Array_6X1 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] bl[0] bl_n[0]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] bl[0] bl_n[0] SP6TVar9Array_4X1
Xinst1x0 vss vdd wl[4] wl[5] bl[0] bl_n[0] SP6TVar9Array_2X1
.ends SP6TVar9Array_6X1

.subckt SP6TVar9CellConnectOut wl bl bl_n vdd vss bit bit_n
Xpu1 vdd bit_n bit vdd sg13_lv_pmos l=1.3e-07 w=1.5e-07
Xpd1 bit bit_n vss vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpu2 vdd bit bit_n vdd sg13_lv_pmos l=1.3e-07 w=1.5e-07
Xpd2 bit_n bit vss vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg1 bit wl bl vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg2 bit_n wl bl_n vss sg13_lv_nmos l=1.3e-07 w=3e-07
.ends SP6TVar9CellConnectOut

.subckt SP6TVar9TestArray_16X8C vss vdd bl bl_n bit bit_n wl
Xarray_0 vss vdd zero zero zero zero zero zero zero zero wl zero zero zero zero zero zero zero array_0_bl[0] array_0_bl_n[0] SP6TVar9Array_16X1BC
Xarray_1 vss vdd zero zero zero zero zero zero zero zero wl zero zero zero zero zero zero zero array_1_bl[0] array_1_bl_n[0] array_1_bl[1] array_1_bl_n[1] SP6TVar9Array_16X2BC
Xarray_2 vss vdd zero zero zero zero zero zero zero zero wl zero zero zero zero zero zero zero array_2_bl[0] array_2_bl_n[0] array_2_bl[1] array_2_bl_n[1] array_2_bl[2] array_2_bl_n[2] array_2_bl[3] array_2_bl_n[3] SP6TVar9Array_16X4BC
Xcolbc_0 vdd vss bl bl_n SP6TVar9BulkConn
Xcolbc_1 vdd vss bl bl_n SP6TVar9BulkConn
Xcolarray_0 vss vdd zero zero zero zero zero zero zero zero bl bl_n SP6TVar9Array_8X1
Xcolarray_1 vss vdd zero zero zero zero zero zero bl bl_n SP6TVar9Array_6X1
Xbc_noconn zero bl bl_n vdd vss SP6TVar9Cell
Xbc_conn wl bl bl_n vdd vss bit bit_n SP6TVar9CellConnectOut
Xzero vdd vss zero zero_x1
.ends SP6TVar9TestArray_16X8C

.subckt SP6TVar9 vss noco_vdd noco_wl noco_bl noco_bl_n co_vdd co_bl co_bl_n co_bit co_bit_n co_wl
Xframe noco_vdd noco_wl NoConn_PAD0x2 co_vdd co_bl_n co_bit co_bit_n NoConn_PAD0x7 NoConn_PAD0x8 NoConn_PAD0x9 vss noco_bl noco_bl_n vss co_bl co_wl NoConn_PAD1x6 NoConn_PAD1x7 NoConn_PAD1x8 NoConn_PAD1x9 PadFrame_SP09
Xtestarray_noco vss noco_vdd noco_bl noco_bl_n noco_wl SP6TVar9TestArray_16X8
Xtestarray_co vss co_vdd co_bl co_bl_n co_bit co_bit_n co_wl SP6TVar9TestArray_16X8C
.ends SP6TVar9

.subckt PadFrame_SP10 PAD0x0 PAD0x1 PAD0x2 PAD0x3 PAD0x4 PAD0x5 PAD0x6 PAD0x7 PAD0x8 PAD0x9 PAD1x0 PAD1x1 PAD1x2 PAD1x3 PAD1x4 PAD1x5 PAD1x6 PAD1x7 PAD1x8 PAD1x9
XPAD0x0 PAD0x0 BondPad
XPAD0x1 PAD0x1 BondPad
XPAD0x2 PAD0x2 BondPad
XPAD0x3 PAD0x3 BondPad
XPAD0x4 PAD0x4 BondPad
XPAD0x5 PAD0x5 BondPad
XPAD0x6 PAD0x6 BondPad
XPAD0x7 PAD0x7 BondPad
XPAD0x8 PAD0x8 BondPad
XPAD0x9 PAD0x9 BondPad
XPAD1x0 PAD1x0 BondPad
XPAD1x1 PAD1x1 BondPad
XPAD1x2 PAD1x2 BondPad
XPAD1x3 PAD1x3 BondPad
XPAD1x4 PAD1x4 BondPad
XPAD1x5 PAD1x5 BondPad
XPAD1x6 PAD1x6 BondPad
XPAD1x7 PAD1x7 BondPad
XPAD1x8 PAD1x8 BondPad
XPAD1x9 PAD1x9 BondPad
.ends PadFrame_SP10

.subckt SP6TVar10Cell wl bl bl_n vdd vss
Xpu1 vdd bit_n bit vdd sg13_lv_pmos l=1.3e-07 w=2e-07
Xpd1 bit bit_n vss vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpu2 vdd bit bit_n vdd sg13_lv_pmos l=1.3e-07 w=2e-07
Xpd2 bit_n bit vss vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg1 bit wl bl vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg2 bit_n wl bl_n vss sg13_lv_nmos l=1.3e-07 w=2e-07
.ends SP6TVar10Cell

.subckt SP6TVar10Array_2X1 vss vdd wl[0] wl[1] bl[0] bl_n[0]
Xinst0x0 wl[0] bl[0] bl_n[0] vdd vss SP6TVar10Cell
Xinst1x0 wl[1] bl[0] bl_n[0] vdd vss SP6TVar10Cell
.ends SP6TVar10Array_2X1

.subckt SP6TVar10Array_2X2 vss vdd wl[0] wl[1] bl[0] bl_n[0] bl[1] bl_n[1]
Xinst0x0 vss vdd wl[0] wl[1] bl[0] bl_n[0] SP6TVar10Array_2X1
Xinst0x1 vss vdd wl[0] wl[1] bl[1] bl_n[1] SP6TVar10Array_2X1
.ends SP6TVar10Array_2X2

.subckt SP6TVar10Array_4X2 vss vdd wl[0] wl[1] wl[2] wl[3] bl[0] bl_n[0] bl[1] bl_n[1]
Xinst0x0 vss vdd wl[0] wl[1] bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar10Array_2X2
Xinst1x0 vss vdd wl[2] wl[3] bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar10Array_2X2
.ends SP6TVar10Array_4X2

.subckt SP6TVar10Array_4X4 vss vdd wl[0] wl[1] wl[2] wl[3] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar10Array_4X2
Xinst0x1 vss vdd wl[0] wl[1] wl[2] wl[3] bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar10Array_4X2
.ends SP6TVar10Array_4X4

.subckt SP6TVar10Array_8X4 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar10Array_4X4
Xinst1x0 vss vdd wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar10Array_4X4
.ends SP6TVar10Array_8X4

.subckt SP6TVar10Array_8X8 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar10Array_8X4
Xinst0x1 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7] SP6TVar10Array_8X4
.ends SP6TVar10Array_8X8

.subckt SP6TVar10BulkConn vdd vss bl bl_n
.ends SP6TVar10BulkConn

.subckt SP6TVar10BulkConnRow_2 vss vdd bl[0] bl_n[0] bl[1] bl_n[1]
Xinst0 vdd vss bl[0] bl_n[0] SP6TVar10BulkConn
Xinst1 vdd vss bl[1] bl_n[1] SP6TVar10BulkConn
.ends SP6TVar10BulkConnRow_2

.subckt SP6TVar10BulkConnRow_4 vss vdd bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3]
Xinst0 vss vdd bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar10BulkConnRow_2
Xinst1 vss vdd bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar10BulkConnRow_2
.ends SP6TVar10BulkConnRow_4

.subckt SP6TVar10BulkConnRow_8 vss vdd bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7]
Xinst0 vss vdd bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar10BulkConnRow_4
Xinst1 vss vdd bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7] SP6TVar10BulkConnRow_4
.ends SP6TVar10BulkConnRow_8

.subckt SP6TVar10Array_16X8BC vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7] SP6TVar10Array_8X8
Xinst1x0 vss vdd wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7] SP6TVar10Array_8X8
Xbottombcrow vss vdd bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7] SP6TVar10BulkConnRow_8
Xtopbcrow vss vdd bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7] SP6TVar10BulkConnRow_8
.ends SP6TVar10Array_16X8BC

.subckt SP6TVar10TestArray_16X8 vss vdd bl bl_n wl
Xarray vss vdd zero zero zero zero zero zero zero zero wl zero zero zero zero zero zero zero bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl bl_n bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7] SP6TVar10Array_16X8BC
Xzero vdd vss zero zero_x1
.ends SP6TVar10TestArray_16X8

.subckt SP6TVar10Array_4X1 vss vdd wl[0] wl[1] wl[2] wl[3] bl[0] bl_n[0]
Xinst0x0 vss vdd wl[0] wl[1] bl[0] bl_n[0] SP6TVar10Array_2X1
Xinst1x0 vss vdd wl[2] wl[3] bl[0] bl_n[0] SP6TVar10Array_2X1
.ends SP6TVar10Array_4X1

.subckt SP6TVar10Array_8X1 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] bl[0] bl_n[0] SP6TVar10Array_4X1
Xinst1x0 vss vdd wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] SP6TVar10Array_4X1
.ends SP6TVar10Array_8X1

.subckt SP6TVar10Array_16X1BC vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] bl[0] bl_n[0]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] SP6TVar10Array_8X1
Xinst1x0 vss vdd wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] bl[0] bl_n[0] SP6TVar10Array_8X1
Xbottombcrow vdd vss bl[0] bl_n[0] SP6TVar10BulkConn
Xtopbcrow vdd vss bl[0] bl_n[0] SP6TVar10BulkConn
.ends SP6TVar10Array_16X1BC

.subckt SP6TVar10Array_8X2 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar10Array_4X2
Xinst1x0 vss vdd wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar10Array_4X2
.ends SP6TVar10Array_8X2

.subckt SP6TVar10Array_16X2BC vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] bl[0] bl_n[0] bl[1] bl_n[1]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar10Array_8X2
Xinst1x0 vss vdd wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar10Array_8X2
Xbottombcrow vss vdd bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar10BulkConnRow_2
Xtopbcrow vss vdd bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar10BulkConnRow_2
.ends SP6TVar10Array_16X2BC

.subckt SP6TVar10Array_16X4BC vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar10Array_8X4
Xinst1x0 vss vdd wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar10Array_8X4
Xbottombcrow vss vdd bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar10BulkConnRow_4
Xtopbcrow vss vdd bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar10BulkConnRow_4
.ends SP6TVar10Array_16X4BC

.subckt SP6TVar10Array_6X1 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] bl[0] bl_n[0]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] bl[0] bl_n[0] SP6TVar10Array_4X1
Xinst1x0 vss vdd wl[4] wl[5] bl[0] bl_n[0] SP6TVar10Array_2X1
.ends SP6TVar10Array_6X1

.subckt SP6TVar10CellConnectOut wl bl bl_n vdd vss bit bit_n
Xpu1 vdd bit_n bit vdd sg13_lv_pmos l=1.3e-07 w=2e-07
Xpd1 bit bit_n vss vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpu2 vdd bit bit_n vdd sg13_lv_pmos l=1.3e-07 w=2e-07
Xpd2 bit_n bit vss vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg1 bit wl bl vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg2 bit_n wl bl_n vss sg13_lv_nmos l=1.3e-07 w=2e-07
.ends SP6TVar10CellConnectOut

.subckt SP6TVar10TestArray_16X8C vss vdd bl bl_n bit bit_n wl
Xarray_0 vss vdd zero zero zero zero zero zero zero zero wl zero zero zero zero zero zero zero array_0_bl[0] array_0_bl_n[0] SP6TVar10Array_16X1BC
Xarray_1 vss vdd zero zero zero zero zero zero zero zero wl zero zero zero zero zero zero zero array_1_bl[0] array_1_bl_n[0] array_1_bl[1] array_1_bl_n[1] SP6TVar10Array_16X2BC
Xarray_2 vss vdd zero zero zero zero zero zero zero zero wl zero zero zero zero zero zero zero array_2_bl[0] array_2_bl_n[0] array_2_bl[1] array_2_bl_n[1] array_2_bl[2] array_2_bl_n[2] array_2_bl[3] array_2_bl_n[3] SP6TVar10Array_16X4BC
Xcolbc_0 vdd vss bl bl_n SP6TVar10BulkConn
Xcolbc_1 vdd vss bl bl_n SP6TVar10BulkConn
Xcolarray_0 vss vdd zero zero zero zero zero zero zero zero bl bl_n SP6TVar10Array_8X1
Xcolarray_1 vss vdd zero zero zero zero zero zero bl bl_n SP6TVar10Array_6X1
Xbc_noconn zero bl bl_n vdd vss SP6TVar10Cell
Xbc_conn wl bl bl_n vdd vss bit bit_n SP6TVar10CellConnectOut
Xzero vdd vss zero zero_x1
.ends SP6TVar10TestArray_16X8C

.subckt SP6TVar10 vss noco_vdd noco_wl noco_bl noco_bl_n co_vdd co_bl co_bl_n co_bit co_bit_n co_wl
Xframe noco_vdd noco_wl NoConn_PAD0x2 co_vdd co_bl_n co_bit co_bit_n NoConn_PAD0x7 NoConn_PAD0x8 NoConn_PAD0x9 vss noco_bl noco_bl_n vss co_bl co_wl NoConn_PAD1x6 NoConn_PAD1x7 NoConn_PAD1x8 NoConn_PAD1x9 PadFrame_SP10
Xtestarray_noco vss noco_vdd noco_bl noco_bl_n noco_wl SP6TVar10TestArray_16X8
Xtestarray_co vss co_vdd co_bl co_bl_n co_bit co_bit_n co_wl SP6TVar10TestArray_16X8C
.ends SP6TVar10

.subckt PadFrame_SP11 PAD0x0 PAD0x1 PAD0x2 PAD0x3 PAD0x4 PAD0x5 PAD0x6 PAD0x7 PAD0x8 PAD0x9 PAD1x0 PAD1x1 PAD1x2 PAD1x3 PAD1x4 PAD1x5 PAD1x6 PAD1x7 PAD1x8 PAD1x9
XPAD0x0 PAD0x0 BondPad
XPAD0x1 PAD0x1 BondPad
XPAD0x2 PAD0x2 BondPad
XPAD0x3 PAD0x3 BondPad
XPAD0x4 PAD0x4 BondPad
XPAD0x5 PAD0x5 BondPad
XPAD0x6 PAD0x6 BondPad
XPAD0x7 PAD0x7 BondPad
XPAD0x8 PAD0x8 BondPad
XPAD0x9 PAD0x9 BondPad
XPAD1x0 PAD1x0 BondPad
XPAD1x1 PAD1x1 BondPad
XPAD1x2 PAD1x2 BondPad
XPAD1x3 PAD1x3 BondPad
XPAD1x4 PAD1x4 BondPad
XPAD1x5 PAD1x5 BondPad
XPAD1x6 PAD1x6 BondPad
XPAD1x7 PAD1x7 BondPad
XPAD1x8 PAD1x8 BondPad
XPAD1x9 PAD1x9 BondPad
.ends PadFrame_SP11

.subckt SP6TVar11Cell wl bl bl_n vdd vss
Xpu1 vdd bit_n bit vdd sg13_lv_pmos l=1.3e-07 w=1.5e-07
Xpd1 bit bit_n vss vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpu2 vdd bit bit_n vdd sg13_lv_pmos l=1.3e-07 w=1.5e-07
Xpd2 bit_n bit vss vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg1 bit wl bl vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg2 bit_n wl bl_n vss sg13_lv_nmos l=1.3e-07 w=2e-07
.ends SP6TVar11Cell

.subckt SP6TVar11Array_2X1 vss vdd wl[0] wl[1] bl[0] bl_n[0]
Xinst0x0 wl[0] bl[0] bl_n[0] vdd vss SP6TVar11Cell
Xinst1x0 wl[1] bl[0] bl_n[0] vdd vss SP6TVar11Cell
.ends SP6TVar11Array_2X1

.subckt SP6TVar11Array_2X2 vss vdd wl[0] wl[1] bl[0] bl_n[0] bl[1] bl_n[1]
Xinst0x0 vss vdd wl[0] wl[1] bl[0] bl_n[0] SP6TVar11Array_2X1
Xinst0x1 vss vdd wl[0] wl[1] bl[1] bl_n[1] SP6TVar11Array_2X1
.ends SP6TVar11Array_2X2

.subckt SP6TVar11Array_4X2 vss vdd wl[0] wl[1] wl[2] wl[3] bl[0] bl_n[0] bl[1] bl_n[1]
Xinst0x0 vss vdd wl[0] wl[1] bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar11Array_2X2
Xinst1x0 vss vdd wl[2] wl[3] bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar11Array_2X2
.ends SP6TVar11Array_4X2

.subckt SP6TVar11Array_4X4 vss vdd wl[0] wl[1] wl[2] wl[3] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar11Array_4X2
Xinst0x1 vss vdd wl[0] wl[1] wl[2] wl[3] bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar11Array_4X2
.ends SP6TVar11Array_4X4

.subckt SP6TVar11Array_8X4 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar11Array_4X4
Xinst1x0 vss vdd wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar11Array_4X4
.ends SP6TVar11Array_8X4

.subckt SP6TVar11Array_8X8 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar11Array_8X4
Xinst0x1 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7] SP6TVar11Array_8X4
.ends SP6TVar11Array_8X8

.subckt SP6TVar11BulkConn vdd vss bl bl_n
.ends SP6TVar11BulkConn

.subckt SP6TVar11BulkConnRow_2 vss vdd bl[0] bl_n[0] bl[1] bl_n[1]
Xinst0 vdd vss bl[0] bl_n[0] SP6TVar11BulkConn
Xinst1 vdd vss bl[1] bl_n[1] SP6TVar11BulkConn
.ends SP6TVar11BulkConnRow_2

.subckt SP6TVar11BulkConnRow_4 vss vdd bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3]
Xinst0 vss vdd bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar11BulkConnRow_2
Xinst1 vss vdd bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar11BulkConnRow_2
.ends SP6TVar11BulkConnRow_4

.subckt SP6TVar11BulkConnRow_8 vss vdd bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7]
Xinst0 vss vdd bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar11BulkConnRow_4
Xinst1 vss vdd bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7] SP6TVar11BulkConnRow_4
.ends SP6TVar11BulkConnRow_8

.subckt SP6TVar11Array_16X8BC vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7] SP6TVar11Array_8X8
Xinst1x0 vss vdd wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7] SP6TVar11Array_8X8
Xbottombcrow vss vdd bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7] SP6TVar11BulkConnRow_8
Xtopbcrow vss vdd bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7] SP6TVar11BulkConnRow_8
.ends SP6TVar11Array_16X8BC

.subckt SP6TVar11TestArray_16X8 vss vdd bl bl_n wl
Xarray vss vdd zero zero zero zero zero zero zero zero wl zero zero zero zero zero zero zero bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl bl_n bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7] SP6TVar11Array_16X8BC
Xzero vdd vss zero zero_x1
.ends SP6TVar11TestArray_16X8

.subckt SP6TVar11Array_4X1 vss vdd wl[0] wl[1] wl[2] wl[3] bl[0] bl_n[0]
Xinst0x0 vss vdd wl[0] wl[1] bl[0] bl_n[0] SP6TVar11Array_2X1
Xinst1x0 vss vdd wl[2] wl[3] bl[0] bl_n[0] SP6TVar11Array_2X1
.ends SP6TVar11Array_4X1

.subckt SP6TVar11Array_8X1 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] bl[0] bl_n[0] SP6TVar11Array_4X1
Xinst1x0 vss vdd wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] SP6TVar11Array_4X1
.ends SP6TVar11Array_8X1

.subckt SP6TVar11Array_16X1BC vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] bl[0] bl_n[0]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] SP6TVar11Array_8X1
Xinst1x0 vss vdd wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] bl[0] bl_n[0] SP6TVar11Array_8X1
Xbottombcrow vdd vss bl[0] bl_n[0] SP6TVar11BulkConn
Xtopbcrow vdd vss bl[0] bl_n[0] SP6TVar11BulkConn
.ends SP6TVar11Array_16X1BC

.subckt SP6TVar11Array_8X2 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar11Array_4X2
Xinst1x0 vss vdd wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar11Array_4X2
.ends SP6TVar11Array_8X2

.subckt SP6TVar11Array_16X2BC vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] bl[0] bl_n[0] bl[1] bl_n[1]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar11Array_8X2
Xinst1x0 vss vdd wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar11Array_8X2
Xbottombcrow vss vdd bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar11BulkConnRow_2
Xtopbcrow vss vdd bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar11BulkConnRow_2
.ends SP6TVar11Array_16X2BC

.subckt SP6TVar11Array_16X4BC vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar11Array_8X4
Xinst1x0 vss vdd wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar11Array_8X4
Xbottombcrow vss vdd bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar11BulkConnRow_4
Xtopbcrow vss vdd bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar11BulkConnRow_4
.ends SP6TVar11Array_16X4BC

.subckt SP6TVar11Array_6X1 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] bl[0] bl_n[0]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] bl[0] bl_n[0] SP6TVar11Array_4X1
Xinst1x0 vss vdd wl[4] wl[5] bl[0] bl_n[0] SP6TVar11Array_2X1
.ends SP6TVar11Array_6X1

.subckt SP6TVar11CellConnectOut wl bl bl_n vdd vss bit bit_n
Xpu1 vdd bit_n bit vdd sg13_lv_pmos l=1.3e-07 w=1.5e-07
Xpd1 bit bit_n vss vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpu2 vdd bit bit_n vdd sg13_lv_pmos l=1.3e-07 w=1.5e-07
Xpd2 bit_n bit vss vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg1 bit wl bl vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg2 bit_n wl bl_n vss sg13_lv_nmos l=1.3e-07 w=2e-07
.ends SP6TVar11CellConnectOut

.subckt SP6TVar11TestArray_16X8C vss vdd bl bl_n bit bit_n wl
Xarray_0 vss vdd zero zero zero zero zero zero zero zero wl zero zero zero zero zero zero zero array_0_bl[0] array_0_bl_n[0] SP6TVar11Array_16X1BC
Xarray_1 vss vdd zero zero zero zero zero zero zero zero wl zero zero zero zero zero zero zero array_1_bl[0] array_1_bl_n[0] array_1_bl[1] array_1_bl_n[1] SP6TVar11Array_16X2BC
Xarray_2 vss vdd zero zero zero zero zero zero zero zero wl zero zero zero zero zero zero zero array_2_bl[0] array_2_bl_n[0] array_2_bl[1] array_2_bl_n[1] array_2_bl[2] array_2_bl_n[2] array_2_bl[3] array_2_bl_n[3] SP6TVar11Array_16X4BC
Xcolbc_0 vdd vss bl bl_n SP6TVar11BulkConn
Xcolbc_1 vdd vss bl bl_n SP6TVar11BulkConn
Xcolarray_0 vss vdd zero zero zero zero zero zero zero zero bl bl_n SP6TVar11Array_8X1
Xcolarray_1 vss vdd zero zero zero zero zero zero bl bl_n SP6TVar11Array_6X1
Xbc_noconn zero bl bl_n vdd vss SP6TVar11Cell
Xbc_conn wl bl bl_n vdd vss bit bit_n SP6TVar11CellConnectOut
Xzero vdd vss zero zero_x1
.ends SP6TVar11TestArray_16X8C

.subckt SP6TVar11 vss noco_vdd noco_wl noco_bl noco_bl_n co_vdd co_bl co_bl_n co_bit co_bit_n co_wl
Xframe noco_vdd noco_wl NoConn_PAD0x2 co_vdd co_bl_n co_bit co_bit_n NoConn_PAD0x7 NoConn_PAD0x8 NoConn_PAD0x9 vss noco_bl noco_bl_n vss co_bl co_wl NoConn_PAD1x6 NoConn_PAD1x7 NoConn_PAD1x8 NoConn_PAD1x9 PadFrame_SP11
Xtestarray_noco vss noco_vdd noco_bl noco_bl_n noco_wl SP6TVar11TestArray_16X8
Xtestarray_co vss co_vdd co_bl co_bl_n co_bit co_bit_n co_wl SP6TVar11TestArray_16X8C
.ends SP6TVar11

.subckt PadFrame_SP12 PAD0x0 PAD0x1 PAD0x2 PAD0x3 PAD0x4 PAD0x5 PAD0x6 PAD0x7 PAD0x8 PAD0x9 PAD1x0 PAD1x1 PAD1x2 PAD1x3 PAD1x4 PAD1x5 PAD1x6 PAD1x7 PAD1x8 PAD1x9
XPAD0x0 PAD0x0 BondPad
XPAD0x1 PAD0x1 BondPad
XPAD0x2 PAD0x2 BondPad
XPAD0x3 PAD0x3 BondPad
XPAD0x4 PAD0x4 BondPad
XPAD0x5 PAD0x5 BondPad
XPAD0x6 PAD0x6 BondPad
XPAD0x7 PAD0x7 BondPad
XPAD0x8 PAD0x8 BondPad
XPAD0x9 PAD0x9 BondPad
XPAD1x0 PAD1x0 BondPad
XPAD1x1 PAD1x1 BondPad
XPAD1x2 PAD1x2 BondPad
XPAD1x3 PAD1x3 BondPad
XPAD1x4 PAD1x4 BondPad
XPAD1x5 PAD1x5 BondPad
XPAD1x6 PAD1x6 BondPad
XPAD1x7 PAD1x7 BondPad
XPAD1x8 PAD1x8 BondPad
XPAD1x9 PAD1x9 BondPad
.ends PadFrame_SP12

.subckt SP6TVar12Cell wl bl bl_n vdd vss
Xpu1 vdd bit_n bit vdd sg13_lv_pmos l=1.3e-07 w=2e-07
Xpd1 bit bit_n vss vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpu2 vdd bit bit_n vdd sg13_lv_pmos l=1.3e-07 w=2e-07
Xpd2 bit_n bit vss vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg1 bit wl bl vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg2 bit_n wl bl_n vss sg13_lv_nmos l=1.3e-07 w=2e-07
.ends SP6TVar12Cell

.subckt SP6TVar12Array_2X1 vss vdd wl[0] wl[1] bl[0] bl_n[0]
Xinst0x0 wl[0] bl[0] bl_n[0] vdd vss SP6TVar12Cell
Xinst1x0 wl[1] bl[0] bl_n[0] vdd vss SP6TVar12Cell
.ends SP6TVar12Array_2X1

.subckt SP6TVar12Array_2X2 vss vdd wl[0] wl[1] bl[0] bl_n[0] bl[1] bl_n[1]
Xinst0x0 vss vdd wl[0] wl[1] bl[0] bl_n[0] SP6TVar12Array_2X1
Xinst0x1 vss vdd wl[0] wl[1] bl[1] bl_n[1] SP6TVar12Array_2X1
.ends SP6TVar12Array_2X2

.subckt SP6TVar12Array_4X2 vss vdd wl[0] wl[1] wl[2] wl[3] bl[0] bl_n[0] bl[1] bl_n[1]
Xinst0x0 vss vdd wl[0] wl[1] bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar12Array_2X2
Xinst1x0 vss vdd wl[2] wl[3] bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar12Array_2X2
.ends SP6TVar12Array_4X2

.subckt SP6TVar12Array_4X4 vss vdd wl[0] wl[1] wl[2] wl[3] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar12Array_4X2
Xinst0x1 vss vdd wl[0] wl[1] wl[2] wl[3] bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar12Array_4X2
.ends SP6TVar12Array_4X4

.subckt SP6TVar12Array_8X4 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar12Array_4X4
Xinst1x0 vss vdd wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar12Array_4X4
.ends SP6TVar12Array_8X4

.subckt SP6TVar12Array_8X8 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar12Array_8X4
Xinst0x1 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7] SP6TVar12Array_8X4
.ends SP6TVar12Array_8X8

.subckt SP6TVar12BulkConn vdd vss bl bl_n
.ends SP6TVar12BulkConn

.subckt SP6TVar12BulkConnRow_2 vss vdd bl[0] bl_n[0] bl[1] bl_n[1]
Xinst0 vdd vss bl[0] bl_n[0] SP6TVar12BulkConn
Xinst1 vdd vss bl[1] bl_n[1] SP6TVar12BulkConn
.ends SP6TVar12BulkConnRow_2

.subckt SP6TVar12BulkConnRow_4 vss vdd bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3]
Xinst0 vss vdd bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar12BulkConnRow_2
Xinst1 vss vdd bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar12BulkConnRow_2
.ends SP6TVar12BulkConnRow_4

.subckt SP6TVar12BulkConnRow_8 vss vdd bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7]
Xinst0 vss vdd bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar12BulkConnRow_4
Xinst1 vss vdd bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7] SP6TVar12BulkConnRow_4
.ends SP6TVar12BulkConnRow_8

.subckt SP6TVar12Array_16X8BC vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7] SP6TVar12Array_8X8
Xinst1x0 vss vdd wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7] SP6TVar12Array_8X8
Xbottombcrow vss vdd bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7] SP6TVar12BulkConnRow_8
Xtopbcrow vss vdd bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7] SP6TVar12BulkConnRow_8
.ends SP6TVar12Array_16X8BC

.subckt SP6TVar12TestArray_16X8 vss vdd bl bl_n wl
Xarray vss vdd zero zero zero zero zero zero zero zero wl zero zero zero zero zero zero zero bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl bl_n bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7] SP6TVar12Array_16X8BC
Xzero vdd vss zero zero_x1
.ends SP6TVar12TestArray_16X8

.subckt SP6TVar12Array_4X1 vss vdd wl[0] wl[1] wl[2] wl[3] bl[0] bl_n[0]
Xinst0x0 vss vdd wl[0] wl[1] bl[0] bl_n[0] SP6TVar12Array_2X1
Xinst1x0 vss vdd wl[2] wl[3] bl[0] bl_n[0] SP6TVar12Array_2X1
.ends SP6TVar12Array_4X1

.subckt SP6TVar12Array_8X1 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] bl[0] bl_n[0] SP6TVar12Array_4X1
Xinst1x0 vss vdd wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] SP6TVar12Array_4X1
.ends SP6TVar12Array_8X1

.subckt SP6TVar12Array_16X1BC vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] bl[0] bl_n[0]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] SP6TVar12Array_8X1
Xinst1x0 vss vdd wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] bl[0] bl_n[0] SP6TVar12Array_8X1
Xbottombcrow vdd vss bl[0] bl_n[0] SP6TVar12BulkConn
Xtopbcrow vdd vss bl[0] bl_n[0] SP6TVar12BulkConn
.ends SP6TVar12Array_16X1BC

.subckt SP6TVar12Array_8X2 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar12Array_4X2
Xinst1x0 vss vdd wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar12Array_4X2
.ends SP6TVar12Array_8X2

.subckt SP6TVar12Array_16X2BC vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] bl[0] bl_n[0] bl[1] bl_n[1]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar12Array_8X2
Xinst1x0 vss vdd wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar12Array_8X2
Xbottombcrow vss vdd bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar12BulkConnRow_2
Xtopbcrow vss vdd bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar12BulkConnRow_2
.ends SP6TVar12Array_16X2BC

.subckt SP6TVar12Array_16X4BC vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar12Array_8X4
Xinst1x0 vss vdd wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar12Array_8X4
Xbottombcrow vss vdd bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar12BulkConnRow_4
Xtopbcrow vss vdd bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar12BulkConnRow_4
.ends SP6TVar12Array_16X4BC

.subckt SP6TVar12Array_6X1 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] bl[0] bl_n[0]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] bl[0] bl_n[0] SP6TVar12Array_4X1
Xinst1x0 vss vdd wl[4] wl[5] bl[0] bl_n[0] SP6TVar12Array_2X1
.ends SP6TVar12Array_6X1

.subckt SP6TVar12CellConnectOut wl bl bl_n vdd vss bit bit_n
Xpu1 vdd bit_n bit vdd sg13_lv_pmos l=1.3e-07 w=2e-07
Xpd1 bit bit_n vss vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpu2 vdd bit bit_n vdd sg13_lv_pmos l=1.3e-07 w=2e-07
Xpd2 bit_n bit vss vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg1 bit wl bl vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg2 bit_n wl bl_n vss sg13_lv_nmos l=1.3e-07 w=2e-07
.ends SP6TVar12CellConnectOut

.subckt SP6TVar12TestArray_16X8C vss vdd bl bl_n bit bit_n wl
Xarray_0 vss vdd zero zero zero zero zero zero zero zero wl zero zero zero zero zero zero zero array_0_bl[0] array_0_bl_n[0] SP6TVar12Array_16X1BC
Xarray_1 vss vdd zero zero zero zero zero zero zero zero wl zero zero zero zero zero zero zero array_1_bl[0] array_1_bl_n[0] array_1_bl[1] array_1_bl_n[1] SP6TVar12Array_16X2BC
Xarray_2 vss vdd zero zero zero zero zero zero zero zero wl zero zero zero zero zero zero zero array_2_bl[0] array_2_bl_n[0] array_2_bl[1] array_2_bl_n[1] array_2_bl[2] array_2_bl_n[2] array_2_bl[3] array_2_bl_n[3] SP6TVar12Array_16X4BC
Xcolbc_0 vdd vss bl bl_n SP6TVar12BulkConn
Xcolbc_1 vdd vss bl bl_n SP6TVar12BulkConn
Xcolarray_0 vss vdd zero zero zero zero zero zero zero zero bl bl_n SP6TVar12Array_8X1
Xcolarray_1 vss vdd zero zero zero zero zero zero bl bl_n SP6TVar12Array_6X1
Xbc_noconn zero bl bl_n vdd vss SP6TVar12Cell
Xbc_conn wl bl bl_n vdd vss bit bit_n SP6TVar12CellConnectOut
Xzero vdd vss zero zero_x1
.ends SP6TVar12TestArray_16X8C

.subckt SP6TVar12 vss noco_vdd noco_wl noco_bl noco_bl_n co_vdd co_bl co_bl_n co_bit co_bit_n co_wl
Xframe noco_vdd noco_wl NoConn_PAD0x2 co_vdd co_bl_n co_bit co_bit_n NoConn_PAD0x7 NoConn_PAD0x8 NoConn_PAD0x9 vss noco_bl noco_bl_n vss co_bl co_wl NoConn_PAD1x6 NoConn_PAD1x7 NoConn_PAD1x8 NoConn_PAD1x9 PadFrame_SP12
Xtestarray_noco vss noco_vdd noco_bl noco_bl_n noco_wl SP6TVar12TestArray_16X8
Xtestarray_co vss co_vdd co_bl co_bl_n co_bit co_bit_n co_wl SP6TVar12TestArray_16X8C
.ends SP6TVar12

.subckt PadFrame_SP13 PAD0x0 PAD0x1 PAD0x2 PAD0x3 PAD0x4 PAD0x5 PAD0x6 PAD0x7 PAD0x8 PAD0x9 PAD1x0 PAD1x1 PAD1x2 PAD1x3 PAD1x4 PAD1x5 PAD1x6 PAD1x7 PAD1x8 PAD1x9
XPAD0x0 PAD0x0 BondPad
XPAD0x1 PAD0x1 BondPad
XPAD0x2 PAD0x2 BondPad
XPAD0x3 PAD0x3 BondPad
XPAD0x4 PAD0x4 BondPad
XPAD0x5 PAD0x5 BondPad
XPAD0x6 PAD0x6 BondPad
XPAD0x7 PAD0x7 BondPad
XPAD0x8 PAD0x8 BondPad
XPAD0x9 PAD0x9 BondPad
XPAD1x0 PAD1x0 BondPad
XPAD1x1 PAD1x1 BondPad
XPAD1x2 PAD1x2 BondPad
XPAD1x3 PAD1x3 BondPad
XPAD1x4 PAD1x4 BondPad
XPAD1x5 PAD1x5 BondPad
XPAD1x6 PAD1x6 BondPad
XPAD1x7 PAD1x7 BondPad
XPAD1x8 PAD1x8 BondPad
XPAD1x9 PAD1x9 BondPad
.ends PadFrame_SP13

.subckt SP6TVar13Cell wl bl bl_n vdd vss
Xpu1 vdd bit_n bit vdd sg13_lv_pmos l=1.3e-07 w=1.5e-07
Xpd1 bit bit_n vss vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpu2 vdd bit bit_n vdd sg13_lv_pmos l=1.3e-07 w=1.5e-07
Xpd2 bit_n bit vss vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg1 bit wl bl vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg2 bit_n wl bl_n vss sg13_lv_nmos l=1.3e-07 w=2e-07
.ends SP6TVar13Cell

.subckt SP6TVar13Array_2X1 vss vdd wl[0] wl[1] bl[0] bl_n[0]
Xinst0x0 wl[0] bl[0] bl_n[0] vdd vss SP6TVar13Cell
Xinst1x0 wl[1] bl[0] bl_n[0] vdd vss SP6TVar13Cell
.ends SP6TVar13Array_2X1

.subckt SP6TVar13Array_2X2 vss vdd wl[0] wl[1] bl[0] bl_n[0] bl[1] bl_n[1]
Xinst0x0 vss vdd wl[0] wl[1] bl[0] bl_n[0] SP6TVar13Array_2X1
Xinst0x1 vss vdd wl[0] wl[1] bl[1] bl_n[1] SP6TVar13Array_2X1
.ends SP6TVar13Array_2X2

.subckt SP6TVar13Array_4X2 vss vdd wl[0] wl[1] wl[2] wl[3] bl[0] bl_n[0] bl[1] bl_n[1]
Xinst0x0 vss vdd wl[0] wl[1] bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar13Array_2X2
Xinst1x0 vss vdd wl[2] wl[3] bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar13Array_2X2
.ends SP6TVar13Array_4X2

.subckt SP6TVar13Array_4X4 vss vdd wl[0] wl[1] wl[2] wl[3] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar13Array_4X2
Xinst0x1 vss vdd wl[0] wl[1] wl[2] wl[3] bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar13Array_4X2
.ends SP6TVar13Array_4X4

.subckt SP6TVar13Array_8X4 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar13Array_4X4
Xinst1x0 vss vdd wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar13Array_4X4
.ends SP6TVar13Array_8X4

.subckt SP6TVar13Array_8X8 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar13Array_8X4
Xinst0x1 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7] SP6TVar13Array_8X4
.ends SP6TVar13Array_8X8

.subckt SP6TVar13BulkConn vdd vss bl bl_n
.ends SP6TVar13BulkConn

.subckt SP6TVar13BulkConnRow_2 vss vdd bl[0] bl_n[0] bl[1] bl_n[1]
Xinst0 vdd vss bl[0] bl_n[0] SP6TVar13BulkConn
Xinst1 vdd vss bl[1] bl_n[1] SP6TVar13BulkConn
.ends SP6TVar13BulkConnRow_2

.subckt SP6TVar13BulkConnRow_4 vss vdd bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3]
Xinst0 vss vdd bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar13BulkConnRow_2
Xinst1 vss vdd bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar13BulkConnRow_2
.ends SP6TVar13BulkConnRow_4

.subckt SP6TVar13BulkConnRow_8 vss vdd bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7]
Xinst0 vss vdd bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar13BulkConnRow_4
Xinst1 vss vdd bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7] SP6TVar13BulkConnRow_4
.ends SP6TVar13BulkConnRow_8

.subckt SP6TVar13Array_16X8BC vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7] SP6TVar13Array_8X8
Xinst1x0 vss vdd wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7] SP6TVar13Array_8X8
Xbottombcrow vss vdd bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7] SP6TVar13BulkConnRow_8
Xtopbcrow vss vdd bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7] SP6TVar13BulkConnRow_8
.ends SP6TVar13Array_16X8BC

.subckt SP6TVar13TestArray_16X8 vss vdd bl bl_n wl
Xarray vss vdd zero zero zero zero zero zero zero zero wl zero zero zero zero zero zero zero bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl bl_n bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7] SP6TVar13Array_16X8BC
Xzero vdd vss zero zero_x1
.ends SP6TVar13TestArray_16X8

.subckt SP6TVar13Array_4X1 vss vdd wl[0] wl[1] wl[2] wl[3] bl[0] bl_n[0]
Xinst0x0 vss vdd wl[0] wl[1] bl[0] bl_n[0] SP6TVar13Array_2X1
Xinst1x0 vss vdd wl[2] wl[3] bl[0] bl_n[0] SP6TVar13Array_2X1
.ends SP6TVar13Array_4X1

.subckt SP6TVar13Array_8X1 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] bl[0] bl_n[0] SP6TVar13Array_4X1
Xinst1x0 vss vdd wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] SP6TVar13Array_4X1
.ends SP6TVar13Array_8X1

.subckt SP6TVar13Array_16X1BC vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] bl[0] bl_n[0]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] SP6TVar13Array_8X1
Xinst1x0 vss vdd wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] bl[0] bl_n[0] SP6TVar13Array_8X1
Xbottombcrow vdd vss bl[0] bl_n[0] SP6TVar13BulkConn
Xtopbcrow vdd vss bl[0] bl_n[0] SP6TVar13BulkConn
.ends SP6TVar13Array_16X1BC

.subckt SP6TVar13Array_8X2 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar13Array_4X2
Xinst1x0 vss vdd wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar13Array_4X2
.ends SP6TVar13Array_8X2

.subckt SP6TVar13Array_16X2BC vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] bl[0] bl_n[0] bl[1] bl_n[1]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar13Array_8X2
Xinst1x0 vss vdd wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar13Array_8X2
Xbottombcrow vss vdd bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar13BulkConnRow_2
Xtopbcrow vss vdd bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar13BulkConnRow_2
.ends SP6TVar13Array_16X2BC

.subckt SP6TVar13Array_16X4BC vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar13Array_8X4
Xinst1x0 vss vdd wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar13Array_8X4
Xbottombcrow vss vdd bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar13BulkConnRow_4
Xtopbcrow vss vdd bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar13BulkConnRow_4
.ends SP6TVar13Array_16X4BC

.subckt SP6TVar13Array_6X1 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] bl[0] bl_n[0]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] bl[0] bl_n[0] SP6TVar13Array_4X1
Xinst1x0 vss vdd wl[4] wl[5] bl[0] bl_n[0] SP6TVar13Array_2X1
.ends SP6TVar13Array_6X1

.subckt SP6TVar13CellConnectOut wl bl bl_n vdd vss bit bit_n
Xpu1 vdd bit_n bit vdd sg13_lv_pmos l=1.3e-07 w=1.5e-07
Xpd1 bit bit_n vss vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpu2 vdd bit bit_n vdd sg13_lv_pmos l=1.3e-07 w=1.5e-07
Xpd2 bit_n bit vss vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg1 bit wl bl vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg2 bit_n wl bl_n vss sg13_lv_nmos l=1.3e-07 w=2e-07
.ends SP6TVar13CellConnectOut

.subckt SP6TVar13TestArray_16X8C vss vdd bl bl_n bit bit_n wl
Xarray_0 vss vdd zero zero zero zero zero zero zero zero wl zero zero zero zero zero zero zero array_0_bl[0] array_0_bl_n[0] SP6TVar13Array_16X1BC
Xarray_1 vss vdd zero zero zero zero zero zero zero zero wl zero zero zero zero zero zero zero array_1_bl[0] array_1_bl_n[0] array_1_bl[1] array_1_bl_n[1] SP6TVar13Array_16X2BC
Xarray_2 vss vdd zero zero zero zero zero zero zero zero wl zero zero zero zero zero zero zero array_2_bl[0] array_2_bl_n[0] array_2_bl[1] array_2_bl_n[1] array_2_bl[2] array_2_bl_n[2] array_2_bl[3] array_2_bl_n[3] SP6TVar13Array_16X4BC
Xcolbc_0 vdd vss bl bl_n SP6TVar13BulkConn
Xcolbc_1 vdd vss bl bl_n SP6TVar13BulkConn
Xcolarray_0 vss vdd zero zero zero zero zero zero zero zero bl bl_n SP6TVar13Array_8X1
Xcolarray_1 vss vdd zero zero zero zero zero zero bl bl_n SP6TVar13Array_6X1
Xbc_noconn zero bl bl_n vdd vss SP6TVar13Cell
Xbc_conn wl bl bl_n vdd vss bit bit_n SP6TVar13CellConnectOut
Xzero vdd vss zero zero_x1
.ends SP6TVar13TestArray_16X8C

.subckt SP6TVar13 vss noco_vdd noco_wl noco_bl noco_bl_n co_vdd co_bl co_bl_n co_bit co_bit_n co_wl
Xframe noco_vdd noco_wl NoConn_PAD0x2 co_vdd co_bl_n co_bit co_bit_n NoConn_PAD0x7 NoConn_PAD0x8 NoConn_PAD0x9 vss noco_bl noco_bl_n vss co_bl co_wl NoConn_PAD1x6 NoConn_PAD1x7 NoConn_PAD1x8 NoConn_PAD1x9 PadFrame_SP13
Xtestarray_noco vss noco_vdd noco_bl noco_bl_n noco_wl SP6TVar13TestArray_16X8
Xtestarray_co vss co_vdd co_bl co_bl_n co_bit co_bit_n co_wl SP6TVar13TestArray_16X8C
.ends SP6TVar13

.subckt PadFrame_SP14 PAD0x0 PAD0x1 PAD0x2 PAD0x3 PAD0x4 PAD0x5 PAD0x6 PAD0x7 PAD0x8 PAD0x9 PAD1x0 PAD1x1 PAD1x2 PAD1x3 PAD1x4 PAD1x5 PAD1x6 PAD1x7 PAD1x8 PAD1x9
XPAD0x0 PAD0x0 BondPad
XPAD0x1 PAD0x1 BondPad
XPAD0x2 PAD0x2 BondPad
XPAD0x3 PAD0x3 BondPad
XPAD0x4 PAD0x4 BondPad
XPAD0x5 PAD0x5 BondPad
XPAD0x6 PAD0x6 BondPad
XPAD0x7 PAD0x7 BondPad
XPAD0x8 PAD0x8 BondPad
XPAD0x9 PAD0x9 BondPad
XPAD1x0 PAD1x0 BondPad
XPAD1x1 PAD1x1 BondPad
XPAD1x2 PAD1x2 BondPad
XPAD1x3 PAD1x3 BondPad
XPAD1x4 PAD1x4 BondPad
XPAD1x5 PAD1x5 BondPad
XPAD1x6 PAD1x6 BondPad
XPAD1x7 PAD1x7 BondPad
XPAD1x8 PAD1x8 BondPad
XPAD1x9 PAD1x9 BondPad
.ends PadFrame_SP14

.subckt SP6TVar14Cell wl bl bl_n vdd vss
Xpu1 vdd bit_n bit vdd sg13_lv_pmos l=1.3e-07 w=3e-07
Xpd1 bit bit_n vss vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpu2 vdd bit bit_n vdd sg13_lv_pmos l=1.3e-07 w=3e-07
Xpd2 bit_n bit vss vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg1 bit wl bl vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg2 bit_n wl bl_n vss sg13_lv_nmos l=1.3e-07 w=3e-07
.ends SP6TVar14Cell

.subckt SP6TVar14Array_2X1 vss vdd wl[0] wl[1] bl[0] bl_n[0]
Xinst0x0 wl[0] bl[0] bl_n[0] vdd vss SP6TVar14Cell
Xinst1x0 wl[1] bl[0] bl_n[0] vdd vss SP6TVar14Cell
.ends SP6TVar14Array_2X1

.subckt SP6TVar14Array_2X2 vss vdd wl[0] wl[1] bl[0] bl_n[0] bl[1] bl_n[1]
Xinst0x0 vss vdd wl[0] wl[1] bl[0] bl_n[0] SP6TVar14Array_2X1
Xinst0x1 vss vdd wl[0] wl[1] bl[1] bl_n[1] SP6TVar14Array_2X1
.ends SP6TVar14Array_2X2

.subckt SP6TVar14Array_4X2 vss vdd wl[0] wl[1] wl[2] wl[3] bl[0] bl_n[0] bl[1] bl_n[1]
Xinst0x0 vss vdd wl[0] wl[1] bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar14Array_2X2
Xinst1x0 vss vdd wl[2] wl[3] bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar14Array_2X2
.ends SP6TVar14Array_4X2

.subckt SP6TVar14Array_4X4 vss vdd wl[0] wl[1] wl[2] wl[3] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar14Array_4X2
Xinst0x1 vss vdd wl[0] wl[1] wl[2] wl[3] bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar14Array_4X2
.ends SP6TVar14Array_4X4

.subckt SP6TVar14Array_8X4 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar14Array_4X4
Xinst1x0 vss vdd wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar14Array_4X4
.ends SP6TVar14Array_8X4

.subckt SP6TVar14Array_8X8 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar14Array_8X4
Xinst0x1 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7] SP6TVar14Array_8X4
.ends SP6TVar14Array_8X8

.subckt SP6TVar14BulkConn vdd vss bl bl_n
.ends SP6TVar14BulkConn

.subckt SP6TVar14BulkConnRow_2 vss vdd bl[0] bl_n[0] bl[1] bl_n[1]
Xinst0 vdd vss bl[0] bl_n[0] SP6TVar14BulkConn
Xinst1 vdd vss bl[1] bl_n[1] SP6TVar14BulkConn
.ends SP6TVar14BulkConnRow_2

.subckt SP6TVar14BulkConnRow_4 vss vdd bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3]
Xinst0 vss vdd bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar14BulkConnRow_2
Xinst1 vss vdd bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar14BulkConnRow_2
.ends SP6TVar14BulkConnRow_4

.subckt SP6TVar14BulkConnRow_8 vss vdd bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7]
Xinst0 vss vdd bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar14BulkConnRow_4
Xinst1 vss vdd bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7] SP6TVar14BulkConnRow_4
.ends SP6TVar14BulkConnRow_8

.subckt SP6TVar14Array_16X8BC vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7] SP6TVar14Array_8X8
Xinst1x0 vss vdd wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7] SP6TVar14Array_8X8
Xbottombcrow vss vdd bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7] SP6TVar14BulkConnRow_8
Xtopbcrow vss vdd bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7] SP6TVar14BulkConnRow_8
.ends SP6TVar14Array_16X8BC

.subckt SP6TVar14TestArray_16X8 vss vdd bl bl_n wl
Xarray vss vdd zero zero zero zero zero zero zero zero wl zero zero zero zero zero zero zero bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl bl_n bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7] SP6TVar14Array_16X8BC
Xzero vdd vss zero zero_x1
.ends SP6TVar14TestArray_16X8

.subckt SP6TVar14Array_4X1 vss vdd wl[0] wl[1] wl[2] wl[3] bl[0] bl_n[0]
Xinst0x0 vss vdd wl[0] wl[1] bl[0] bl_n[0] SP6TVar14Array_2X1
Xinst1x0 vss vdd wl[2] wl[3] bl[0] bl_n[0] SP6TVar14Array_2X1
.ends SP6TVar14Array_4X1

.subckt SP6TVar14Array_8X1 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] bl[0] bl_n[0] SP6TVar14Array_4X1
Xinst1x0 vss vdd wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] SP6TVar14Array_4X1
.ends SP6TVar14Array_8X1

.subckt SP6TVar14Array_16X1BC vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] bl[0] bl_n[0]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] SP6TVar14Array_8X1
Xinst1x0 vss vdd wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] bl[0] bl_n[0] SP6TVar14Array_8X1
Xbottombcrow vdd vss bl[0] bl_n[0] SP6TVar14BulkConn
Xtopbcrow vdd vss bl[0] bl_n[0] SP6TVar14BulkConn
.ends SP6TVar14Array_16X1BC

.subckt SP6TVar14Array_8X2 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar14Array_4X2
Xinst1x0 vss vdd wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar14Array_4X2
.ends SP6TVar14Array_8X2

.subckt SP6TVar14Array_16X2BC vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] bl[0] bl_n[0] bl[1] bl_n[1]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar14Array_8X2
Xinst1x0 vss vdd wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar14Array_8X2
Xbottombcrow vss vdd bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar14BulkConnRow_2
Xtopbcrow vss vdd bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar14BulkConnRow_2
.ends SP6TVar14Array_16X2BC

.subckt SP6TVar14Array_16X4BC vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar14Array_8X4
Xinst1x0 vss vdd wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar14Array_8X4
Xbottombcrow vss vdd bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar14BulkConnRow_4
Xtopbcrow vss vdd bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar14BulkConnRow_4
.ends SP6TVar14Array_16X4BC

.subckt SP6TVar14Array_6X1 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] bl[0] bl_n[0]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] bl[0] bl_n[0] SP6TVar14Array_4X1
Xinst1x0 vss vdd wl[4] wl[5] bl[0] bl_n[0] SP6TVar14Array_2X1
.ends SP6TVar14Array_6X1

.subckt SP6TVar14CellConnectOut wl bl bl_n vdd vss bit bit_n
Xpu1 vdd bit_n bit vdd sg13_lv_pmos l=1.3e-07 w=3e-07
Xpd1 bit bit_n vss vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpu2 vdd bit bit_n vdd sg13_lv_pmos l=1.3e-07 w=3e-07
Xpd2 bit_n bit vss vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg1 bit wl bl vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg2 bit_n wl bl_n vss sg13_lv_nmos l=1.3e-07 w=3e-07
.ends SP6TVar14CellConnectOut

.subckt SP6TVar14TestArray_16X8C vss vdd bl bl_n bit bit_n wl
Xarray_0 vss vdd zero zero zero zero zero zero zero zero wl zero zero zero zero zero zero zero array_0_bl[0] array_0_bl_n[0] SP6TVar14Array_16X1BC
Xarray_1 vss vdd zero zero zero zero zero zero zero zero wl zero zero zero zero zero zero zero array_1_bl[0] array_1_bl_n[0] array_1_bl[1] array_1_bl_n[1] SP6TVar14Array_16X2BC
Xarray_2 vss vdd zero zero zero zero zero zero zero zero wl zero zero zero zero zero zero zero array_2_bl[0] array_2_bl_n[0] array_2_bl[1] array_2_bl_n[1] array_2_bl[2] array_2_bl_n[2] array_2_bl[3] array_2_bl_n[3] SP6TVar14Array_16X4BC
Xcolbc_0 vdd vss bl bl_n SP6TVar14BulkConn
Xcolbc_1 vdd vss bl bl_n SP6TVar14BulkConn
Xcolarray_0 vss vdd zero zero zero zero zero zero zero zero bl bl_n SP6TVar14Array_8X1
Xcolarray_1 vss vdd zero zero zero zero zero zero bl bl_n SP6TVar14Array_6X1
Xbc_noconn zero bl bl_n vdd vss SP6TVar14Cell
Xbc_conn wl bl bl_n vdd vss bit bit_n SP6TVar14CellConnectOut
Xzero vdd vss zero zero_x1
.ends SP6TVar14TestArray_16X8C

.subckt SP6TVar14 vss noco_vdd noco_wl noco_bl noco_bl_n co_vdd co_bl co_bl_n co_bit co_bit_n co_wl
Xframe noco_vdd noco_wl NoConn_PAD0x2 co_vdd co_bl_n co_bit co_bit_n NoConn_PAD0x7 NoConn_PAD0x8 NoConn_PAD0x9 vss noco_bl noco_bl_n vss co_bl co_wl NoConn_PAD1x6 NoConn_PAD1x7 NoConn_PAD1x8 NoConn_PAD1x9 PadFrame_SP14
Xtestarray_noco vss noco_vdd noco_bl noco_bl_n noco_wl SP6TVar14TestArray_16X8
Xtestarray_co vss co_vdd co_bl co_bl_n co_bit co_bit_n co_wl SP6TVar14TestArray_16X8C
.ends SP6TVar14

.subckt PadFrame_SP15 PAD0x0 PAD0x1 PAD0x2 PAD0x3 PAD0x4 PAD0x5 PAD0x6 PAD0x7 PAD0x8 PAD0x9 PAD1x0 PAD1x1 PAD1x2 PAD1x3 PAD1x4 PAD1x5 PAD1x6 PAD1x7 PAD1x8 PAD1x9
XPAD0x0 PAD0x0 BondPad
XPAD0x1 PAD0x1 BondPad
XPAD0x2 PAD0x2 BondPad
XPAD0x3 PAD0x3 BondPad
XPAD0x4 PAD0x4 BondPad
XPAD0x5 PAD0x5 BondPad
XPAD0x6 PAD0x6 BondPad
XPAD0x7 PAD0x7 BondPad
XPAD0x8 PAD0x8 BondPad
XPAD0x9 PAD0x9 BondPad
XPAD1x0 PAD1x0 BondPad
XPAD1x1 PAD1x1 BondPad
XPAD1x2 PAD1x2 BondPad
XPAD1x3 PAD1x3 BondPad
XPAD1x4 PAD1x4 BondPad
XPAD1x5 PAD1x5 BondPad
XPAD1x6 PAD1x6 BondPad
XPAD1x7 PAD1x7 BondPad
XPAD1x8 PAD1x8 BondPad
XPAD1x9 PAD1x9 BondPad
.ends PadFrame_SP15

.subckt SP6TVar15Cell wl bl bl_n vdd vss
Xpu1 vdd bit_n bit vdd sg13_lv_pmos l=1.3e-07 w=2e-07
Xpd1 bit bit_n vss vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpu2 vdd bit bit_n vdd sg13_lv_pmos l=1.3e-07 w=2e-07
Xpd2 bit_n bit vss vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg1 bit wl bl vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg2 bit_n wl bl_n vss sg13_lv_nmos l=1.3e-07 w=3e-07
.ends SP6TVar15Cell

.subckt SP6TVar15Array_2X1 vss vdd wl[0] wl[1] bl[0] bl_n[0]
Xinst0x0 wl[0] bl[0] bl_n[0] vdd vss SP6TVar15Cell
Xinst1x0 wl[1] bl[0] bl_n[0] vdd vss SP6TVar15Cell
.ends SP6TVar15Array_2X1

.subckt SP6TVar15Array_2X2 vss vdd wl[0] wl[1] bl[0] bl_n[0] bl[1] bl_n[1]
Xinst0x0 vss vdd wl[0] wl[1] bl[0] bl_n[0] SP6TVar15Array_2X1
Xinst0x1 vss vdd wl[0] wl[1] bl[1] bl_n[1] SP6TVar15Array_2X1
.ends SP6TVar15Array_2X2

.subckt SP6TVar15Array_4X2 vss vdd wl[0] wl[1] wl[2] wl[3] bl[0] bl_n[0] bl[1] bl_n[1]
Xinst0x0 vss vdd wl[0] wl[1] bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar15Array_2X2
Xinst1x0 vss vdd wl[2] wl[3] bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar15Array_2X2
.ends SP6TVar15Array_4X2

.subckt SP6TVar15Array_4X4 vss vdd wl[0] wl[1] wl[2] wl[3] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar15Array_4X2
Xinst0x1 vss vdd wl[0] wl[1] wl[2] wl[3] bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar15Array_4X2
.ends SP6TVar15Array_4X4

.subckt SP6TVar15Array_8X4 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar15Array_4X4
Xinst1x0 vss vdd wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar15Array_4X4
.ends SP6TVar15Array_8X4

.subckt SP6TVar15Array_8X8 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar15Array_8X4
Xinst0x1 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7] SP6TVar15Array_8X4
.ends SP6TVar15Array_8X8

.subckt SP6TVar15BulkConn vdd vss bl bl_n
.ends SP6TVar15BulkConn

.subckt SP6TVar15BulkConnRow_2 vss vdd bl[0] bl_n[0] bl[1] bl_n[1]
Xinst0 vdd vss bl[0] bl_n[0] SP6TVar15BulkConn
Xinst1 vdd vss bl[1] bl_n[1] SP6TVar15BulkConn
.ends SP6TVar15BulkConnRow_2

.subckt SP6TVar15BulkConnRow_4 vss vdd bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3]
Xinst0 vss vdd bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar15BulkConnRow_2
Xinst1 vss vdd bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar15BulkConnRow_2
.ends SP6TVar15BulkConnRow_4

.subckt SP6TVar15BulkConnRow_8 vss vdd bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7]
Xinst0 vss vdd bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar15BulkConnRow_4
Xinst1 vss vdd bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7] SP6TVar15BulkConnRow_4
.ends SP6TVar15BulkConnRow_8

.subckt SP6TVar15Array_16X8BC vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7] SP6TVar15Array_8X8
Xinst1x0 vss vdd wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7] SP6TVar15Array_8X8
Xbottombcrow vss vdd bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7] SP6TVar15BulkConnRow_8
Xtopbcrow vss vdd bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7] SP6TVar15BulkConnRow_8
.ends SP6TVar15Array_16X8BC

.subckt SP6TVar15TestArray_16X8 vss vdd bl bl_n wl
Xarray vss vdd zero zero zero zero zero zero zero zero wl zero zero zero zero zero zero zero bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl bl_n bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7] SP6TVar15Array_16X8BC
Xzero vdd vss zero zero_x1
.ends SP6TVar15TestArray_16X8

.subckt SP6TVar15Array_4X1 vss vdd wl[0] wl[1] wl[2] wl[3] bl[0] bl_n[0]
Xinst0x0 vss vdd wl[0] wl[1] bl[0] bl_n[0] SP6TVar15Array_2X1
Xinst1x0 vss vdd wl[2] wl[3] bl[0] bl_n[0] SP6TVar15Array_2X1
.ends SP6TVar15Array_4X1

.subckt SP6TVar15Array_8X1 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] bl[0] bl_n[0] SP6TVar15Array_4X1
Xinst1x0 vss vdd wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] SP6TVar15Array_4X1
.ends SP6TVar15Array_8X1

.subckt SP6TVar15Array_16X1BC vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] bl[0] bl_n[0]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] SP6TVar15Array_8X1
Xinst1x0 vss vdd wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] bl[0] bl_n[0] SP6TVar15Array_8X1
Xbottombcrow vdd vss bl[0] bl_n[0] SP6TVar15BulkConn
Xtopbcrow vdd vss bl[0] bl_n[0] SP6TVar15BulkConn
.ends SP6TVar15Array_16X1BC

.subckt SP6TVar15Array_8X2 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar15Array_4X2
Xinst1x0 vss vdd wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar15Array_4X2
.ends SP6TVar15Array_8X2

.subckt SP6TVar15Array_16X2BC vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] bl[0] bl_n[0] bl[1] bl_n[1]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar15Array_8X2
Xinst1x0 vss vdd wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar15Array_8X2
Xbottombcrow vss vdd bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar15BulkConnRow_2
Xtopbcrow vss vdd bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar15BulkConnRow_2
.ends SP6TVar15Array_16X2BC

.subckt SP6TVar15Array_16X4BC vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar15Array_8X4
Xinst1x0 vss vdd wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar15Array_8X4
Xbottombcrow vss vdd bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar15BulkConnRow_4
Xtopbcrow vss vdd bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar15BulkConnRow_4
.ends SP6TVar15Array_16X4BC

.subckt SP6TVar15Array_6X1 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] bl[0] bl_n[0]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] bl[0] bl_n[0] SP6TVar15Array_4X1
Xinst1x0 vss vdd wl[4] wl[5] bl[0] bl_n[0] SP6TVar15Array_2X1
.ends SP6TVar15Array_6X1

.subckt SP6TVar15CellConnectOut wl bl bl_n vdd vss bit bit_n
Xpu1 vdd bit_n bit vdd sg13_lv_pmos l=1.3e-07 w=2e-07
Xpd1 bit bit_n vss vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpu2 vdd bit bit_n vdd sg13_lv_pmos l=1.3e-07 w=2e-07
Xpd2 bit_n bit vss vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg1 bit wl bl vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg2 bit_n wl bl_n vss sg13_lv_nmos l=1.3e-07 w=3e-07
.ends SP6TVar15CellConnectOut

.subckt SP6TVar15TestArray_16X8C vss vdd bl bl_n bit bit_n wl
Xarray_0 vss vdd zero zero zero zero zero zero zero zero wl zero zero zero zero zero zero zero array_0_bl[0] array_0_bl_n[0] SP6TVar15Array_16X1BC
Xarray_1 vss vdd zero zero zero zero zero zero zero zero wl zero zero zero zero zero zero zero array_1_bl[0] array_1_bl_n[0] array_1_bl[1] array_1_bl_n[1] SP6TVar15Array_16X2BC
Xarray_2 vss vdd zero zero zero zero zero zero zero zero wl zero zero zero zero zero zero zero array_2_bl[0] array_2_bl_n[0] array_2_bl[1] array_2_bl_n[1] array_2_bl[2] array_2_bl_n[2] array_2_bl[3] array_2_bl_n[3] SP6TVar15Array_16X4BC
Xcolbc_0 vdd vss bl bl_n SP6TVar15BulkConn
Xcolbc_1 vdd vss bl bl_n SP6TVar15BulkConn
Xcolarray_0 vss vdd zero zero zero zero zero zero zero zero bl bl_n SP6TVar15Array_8X1
Xcolarray_1 vss vdd zero zero zero zero zero zero bl bl_n SP6TVar15Array_6X1
Xbc_noconn zero bl bl_n vdd vss SP6TVar15Cell
Xbc_conn wl bl bl_n vdd vss bit bit_n SP6TVar15CellConnectOut
Xzero vdd vss zero zero_x1
.ends SP6TVar15TestArray_16X8C

.subckt SP6TVar15 vss noco_vdd noco_wl noco_bl noco_bl_n co_vdd co_bl co_bl_n co_bit co_bit_n co_wl
Xframe noco_vdd noco_wl NoConn_PAD0x2 co_vdd co_bl_n co_bit co_bit_n NoConn_PAD0x7 NoConn_PAD0x8 NoConn_PAD0x9 vss noco_bl noco_bl_n vss co_bl co_wl NoConn_PAD1x6 NoConn_PAD1x7 NoConn_PAD1x8 NoConn_PAD1x9 PadFrame_SP15
Xtestarray_noco vss noco_vdd noco_bl noco_bl_n noco_wl SP6TVar15TestArray_16X8
Xtestarray_co vss co_vdd co_bl co_bl_n co_bit co_bit_n co_wl SP6TVar15TestArray_16X8C
.ends SP6TVar15

.subckt PadFrame_SP16 PAD0x0 PAD0x1 PAD0x2 PAD0x3 PAD0x4 PAD0x5 PAD0x6 PAD0x7 PAD0x8 PAD0x9 PAD1x0 PAD1x1 PAD1x2 PAD1x3 PAD1x4 PAD1x5 PAD1x6 PAD1x7 PAD1x8 PAD1x9
XPAD0x0 PAD0x0 BondPad
XPAD0x1 PAD0x1 BondPad
XPAD0x2 PAD0x2 BondPad
XPAD0x3 PAD0x3 BondPad
XPAD0x4 PAD0x4 BondPad
XPAD0x5 PAD0x5 BondPad
XPAD0x6 PAD0x6 BondPad
XPAD0x7 PAD0x7 BondPad
XPAD0x8 PAD0x8 BondPad
XPAD0x9 PAD0x9 BondPad
XPAD1x0 PAD1x0 BondPad
XPAD1x1 PAD1x1 BondPad
XPAD1x2 PAD1x2 BondPad
XPAD1x3 PAD1x3 BondPad
XPAD1x4 PAD1x4 BondPad
XPAD1x5 PAD1x5 BondPad
XPAD1x6 PAD1x6 BondPad
XPAD1x7 PAD1x7 BondPad
XPAD1x8 PAD1x8 BondPad
XPAD1x9 PAD1x9 BondPad
.ends PadFrame_SP16

.subckt SP6TVar16Cell wl bl bl_n vdd vss
Xpu1 vdd bit_n bit vdd sg13_lv_pmos l=1.3e-07 w=1.5e-07
Xpd1 bit bit_n vss vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpu2 vdd bit bit_n vdd sg13_lv_pmos l=1.3e-07 w=1.5e-07
Xpd2 bit_n bit vss vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg1 bit wl bl vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg2 bit_n wl bl_n vss sg13_lv_nmos l=1.3e-07 w=3e-07
.ends SP6TVar16Cell

.subckt SP6TVar16Array_2X1 vss vdd wl[0] wl[1] bl[0] bl_n[0]
Xinst0x0 wl[0] bl[0] bl_n[0] vdd vss SP6TVar16Cell
Xinst1x0 wl[1] bl[0] bl_n[0] vdd vss SP6TVar16Cell
.ends SP6TVar16Array_2X1

.subckt SP6TVar16Array_2X2 vss vdd wl[0] wl[1] bl[0] bl_n[0] bl[1] bl_n[1]
Xinst0x0 vss vdd wl[0] wl[1] bl[0] bl_n[0] SP6TVar16Array_2X1
Xinst0x1 vss vdd wl[0] wl[1] bl[1] bl_n[1] SP6TVar16Array_2X1
.ends SP6TVar16Array_2X2

.subckt SP6TVar16Array_4X2 vss vdd wl[0] wl[1] wl[2] wl[3] bl[0] bl_n[0] bl[1] bl_n[1]
Xinst0x0 vss vdd wl[0] wl[1] bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar16Array_2X2
Xinst1x0 vss vdd wl[2] wl[3] bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar16Array_2X2
.ends SP6TVar16Array_4X2

.subckt SP6TVar16Array_4X4 vss vdd wl[0] wl[1] wl[2] wl[3] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar16Array_4X2
Xinst0x1 vss vdd wl[0] wl[1] wl[2] wl[3] bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar16Array_4X2
.ends SP6TVar16Array_4X4

.subckt SP6TVar16Array_8X4 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar16Array_4X4
Xinst1x0 vss vdd wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar16Array_4X4
.ends SP6TVar16Array_8X4

.subckt SP6TVar16Array_8X8 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar16Array_8X4
Xinst0x1 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7] SP6TVar16Array_8X4
.ends SP6TVar16Array_8X8

.subckt SP6TVar16BulkConn vdd vss bl bl_n
.ends SP6TVar16BulkConn

.subckt SP6TVar16BulkConnRow_2 vss vdd bl[0] bl_n[0] bl[1] bl_n[1]
Xinst0 vdd vss bl[0] bl_n[0] SP6TVar16BulkConn
Xinst1 vdd vss bl[1] bl_n[1] SP6TVar16BulkConn
.ends SP6TVar16BulkConnRow_2

.subckt SP6TVar16BulkConnRow_4 vss vdd bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3]
Xinst0 vss vdd bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar16BulkConnRow_2
Xinst1 vss vdd bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar16BulkConnRow_2
.ends SP6TVar16BulkConnRow_4

.subckt SP6TVar16BulkConnRow_8 vss vdd bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7]
Xinst0 vss vdd bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar16BulkConnRow_4
Xinst1 vss vdd bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7] SP6TVar16BulkConnRow_4
.ends SP6TVar16BulkConnRow_8

.subckt SP6TVar16Array_16X8BC vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7] SP6TVar16Array_8X8
Xinst1x0 vss vdd wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7] SP6TVar16Array_8X8
Xbottombcrow vss vdd bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7] SP6TVar16BulkConnRow_8
Xtopbcrow vss vdd bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7] SP6TVar16BulkConnRow_8
.ends SP6TVar16Array_16X8BC

.subckt SP6TVar16TestArray_16X8 vss vdd bl bl_n wl
Xarray vss vdd zero zero zero zero zero zero zero zero wl zero zero zero zero zero zero zero bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl bl_n bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7] SP6TVar16Array_16X8BC
Xzero vdd vss zero zero_x1
.ends SP6TVar16TestArray_16X8

.subckt SP6TVar16Array_4X1 vss vdd wl[0] wl[1] wl[2] wl[3] bl[0] bl_n[0]
Xinst0x0 vss vdd wl[0] wl[1] bl[0] bl_n[0] SP6TVar16Array_2X1
Xinst1x0 vss vdd wl[2] wl[3] bl[0] bl_n[0] SP6TVar16Array_2X1
.ends SP6TVar16Array_4X1

.subckt SP6TVar16Array_8X1 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] bl[0] bl_n[0] SP6TVar16Array_4X1
Xinst1x0 vss vdd wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] SP6TVar16Array_4X1
.ends SP6TVar16Array_8X1

.subckt SP6TVar16Array_16X1BC vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] bl[0] bl_n[0]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] SP6TVar16Array_8X1
Xinst1x0 vss vdd wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] bl[0] bl_n[0] SP6TVar16Array_8X1
Xbottombcrow vdd vss bl[0] bl_n[0] SP6TVar16BulkConn
Xtopbcrow vdd vss bl[0] bl_n[0] SP6TVar16BulkConn
.ends SP6TVar16Array_16X1BC

.subckt SP6TVar16Array_8X2 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar16Array_4X2
Xinst1x0 vss vdd wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar16Array_4X2
.ends SP6TVar16Array_8X2

.subckt SP6TVar16Array_16X2BC vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] bl[0] bl_n[0] bl[1] bl_n[1]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar16Array_8X2
Xinst1x0 vss vdd wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar16Array_8X2
Xbottombcrow vss vdd bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar16BulkConnRow_2
Xtopbcrow vss vdd bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar16BulkConnRow_2
.ends SP6TVar16Array_16X2BC

.subckt SP6TVar16Array_16X4BC vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar16Array_8X4
Xinst1x0 vss vdd wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar16Array_8X4
Xbottombcrow vss vdd bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar16BulkConnRow_4
Xtopbcrow vss vdd bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar16BulkConnRow_4
.ends SP6TVar16Array_16X4BC

.subckt SP6TVar16Array_6X1 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] bl[0] bl_n[0]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] bl[0] bl_n[0] SP6TVar16Array_4X1
Xinst1x0 vss vdd wl[4] wl[5] bl[0] bl_n[0] SP6TVar16Array_2X1
.ends SP6TVar16Array_6X1

.subckt SP6TVar16CellConnectOut wl bl bl_n vdd vss bit bit_n
Xpu1 vdd bit_n bit vdd sg13_lv_pmos l=1.3e-07 w=1.5e-07
Xpd1 bit bit_n vss vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpu2 vdd bit bit_n vdd sg13_lv_pmos l=1.3e-07 w=1.5e-07
Xpd2 bit_n bit vss vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg1 bit wl bl vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg2 bit_n wl bl_n vss sg13_lv_nmos l=1.3e-07 w=3e-07
.ends SP6TVar16CellConnectOut

.subckt SP6TVar16TestArray_16X8C vss vdd bl bl_n bit bit_n wl
Xarray_0 vss vdd zero zero zero zero zero zero zero zero wl zero zero zero zero zero zero zero array_0_bl[0] array_0_bl_n[0] SP6TVar16Array_16X1BC
Xarray_1 vss vdd zero zero zero zero zero zero zero zero wl zero zero zero zero zero zero zero array_1_bl[0] array_1_bl_n[0] array_1_bl[1] array_1_bl_n[1] SP6TVar16Array_16X2BC
Xarray_2 vss vdd zero zero zero zero zero zero zero zero wl zero zero zero zero zero zero zero array_2_bl[0] array_2_bl_n[0] array_2_bl[1] array_2_bl_n[1] array_2_bl[2] array_2_bl_n[2] array_2_bl[3] array_2_bl_n[3] SP6TVar16Array_16X4BC
Xcolbc_0 vdd vss bl bl_n SP6TVar16BulkConn
Xcolbc_1 vdd vss bl bl_n SP6TVar16BulkConn
Xcolarray_0 vss vdd zero zero zero zero zero zero zero zero bl bl_n SP6TVar16Array_8X1
Xcolarray_1 vss vdd zero zero zero zero zero zero bl bl_n SP6TVar16Array_6X1
Xbc_noconn zero bl bl_n vdd vss SP6TVar16Cell
Xbc_conn wl bl bl_n vdd vss bit bit_n SP6TVar16CellConnectOut
Xzero vdd vss zero zero_x1
.ends SP6TVar16TestArray_16X8C

.subckt SP6TVar16 vss noco_vdd noco_wl noco_bl noco_bl_n co_vdd co_bl co_bl_n co_bit co_bit_n co_wl
Xframe noco_vdd noco_wl NoConn_PAD0x2 co_vdd co_bl_n co_bit co_bit_n NoConn_PAD0x7 NoConn_PAD0x8 NoConn_PAD0x9 vss noco_bl noco_bl_n vss co_bl co_wl NoConn_PAD1x6 NoConn_PAD1x7 NoConn_PAD1x8 NoConn_PAD1x9 PadFrame_SP16
Xtestarray_noco vss noco_vdd noco_bl noco_bl_n noco_wl SP6TVar16TestArray_16X8
Xtestarray_co vss co_vdd co_bl co_bl_n co_bit co_bit_n co_wl SP6TVar16TestArray_16X8C
.ends SP6TVar16

.subckt PadFrame_SP17 PAD0x0 PAD0x1 PAD0x2 PAD0x3 PAD0x4 PAD0x5 PAD0x6 PAD0x7 PAD0x8 PAD0x9 PAD1x0 PAD1x1 PAD1x2 PAD1x3 PAD1x4 PAD1x5 PAD1x6 PAD1x7 PAD1x8 PAD1x9
XPAD0x0 PAD0x0 BondPad
XPAD0x1 PAD0x1 BondPad
XPAD0x2 PAD0x2 BondPad
XPAD0x3 PAD0x3 BondPad
XPAD0x4 PAD0x4 BondPad
XPAD0x5 PAD0x5 BondPad
XPAD0x6 PAD0x6 BondPad
XPAD0x7 PAD0x7 BondPad
XPAD0x8 PAD0x8 BondPad
XPAD0x9 PAD0x9 BondPad
XPAD1x0 PAD1x0 BondPad
XPAD1x1 PAD1x1 BondPad
XPAD1x2 PAD1x2 BondPad
XPAD1x3 PAD1x3 BondPad
XPAD1x4 PAD1x4 BondPad
XPAD1x5 PAD1x5 BondPad
XPAD1x6 PAD1x6 BondPad
XPAD1x7 PAD1x7 BondPad
XPAD1x8 PAD1x8 BondPad
XPAD1x9 PAD1x9 BondPad
.ends PadFrame_SP17

.subckt SP6TVar17Cell wl bl bl_n vdd vss
Xpu1 vdd bit_n bit vdd sg13_lv_pmos l=1.3e-07 w=2e-07
Xpd1 bit bit_n vss vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpu2 vdd bit bit_n vdd sg13_lv_pmos l=1.3e-07 w=2e-07
Xpd2 bit_n bit vss vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg1 bit wl bl vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg2 bit_n wl bl_n vss sg13_lv_nmos l=1.3e-07 w=2e-07
.ends SP6TVar17Cell

.subckt SP6TVar17Array_2X1 vss vdd wl[0] wl[1] bl[0] bl_n[0]
Xinst0x0 wl[0] bl[0] bl_n[0] vdd vss SP6TVar17Cell
Xinst1x0 wl[1] bl[0] bl_n[0] vdd vss SP6TVar17Cell
.ends SP6TVar17Array_2X1

.subckt SP6TVar17Array_2X2 vss vdd wl[0] wl[1] bl[0] bl_n[0] bl[1] bl_n[1]
Xinst0x0 vss vdd wl[0] wl[1] bl[0] bl_n[0] SP6TVar17Array_2X1
Xinst0x1 vss vdd wl[0] wl[1] bl[1] bl_n[1] SP6TVar17Array_2X1
.ends SP6TVar17Array_2X2

.subckt SP6TVar17Array_4X2 vss vdd wl[0] wl[1] wl[2] wl[3] bl[0] bl_n[0] bl[1] bl_n[1]
Xinst0x0 vss vdd wl[0] wl[1] bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar17Array_2X2
Xinst1x0 vss vdd wl[2] wl[3] bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar17Array_2X2
.ends SP6TVar17Array_4X2

.subckt SP6TVar17Array_4X4 vss vdd wl[0] wl[1] wl[2] wl[3] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar17Array_4X2
Xinst0x1 vss vdd wl[0] wl[1] wl[2] wl[3] bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar17Array_4X2
.ends SP6TVar17Array_4X4

.subckt SP6TVar17Array_8X4 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar17Array_4X4
Xinst1x0 vss vdd wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar17Array_4X4
.ends SP6TVar17Array_8X4

.subckt SP6TVar17Array_8X8 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar17Array_8X4
Xinst0x1 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7] SP6TVar17Array_8X4
.ends SP6TVar17Array_8X8

.subckt SP6TVar17BulkConn vdd vss bl bl_n
.ends SP6TVar17BulkConn

.subckt SP6TVar17BulkConnRow_2 vss vdd bl[0] bl_n[0] bl[1] bl_n[1]
Xinst0 vdd vss bl[0] bl_n[0] SP6TVar17BulkConn
Xinst1 vdd vss bl[1] bl_n[1] SP6TVar17BulkConn
.ends SP6TVar17BulkConnRow_2

.subckt SP6TVar17BulkConnRow_4 vss vdd bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3]
Xinst0 vss vdd bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar17BulkConnRow_2
Xinst1 vss vdd bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar17BulkConnRow_2
.ends SP6TVar17BulkConnRow_4

.subckt SP6TVar17BulkConnRow_8 vss vdd bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7]
Xinst0 vss vdd bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar17BulkConnRow_4
Xinst1 vss vdd bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7] SP6TVar17BulkConnRow_4
.ends SP6TVar17BulkConnRow_8

.subckt SP6TVar17Array_16X8BC vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7] SP6TVar17Array_8X8
Xinst1x0 vss vdd wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7] SP6TVar17Array_8X8
Xbottombcrow vss vdd bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7] SP6TVar17BulkConnRow_8
Xtopbcrow vss vdd bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7] SP6TVar17BulkConnRow_8
.ends SP6TVar17Array_16X8BC

.subckt SP6TVar17TestArray_16X8 vss vdd bl bl_n wl
Xarray vss vdd zero zero zero zero zero zero zero zero wl zero zero zero zero zero zero zero bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl bl_n bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7] SP6TVar17Array_16X8BC
Xzero vdd vss zero zero_x1
.ends SP6TVar17TestArray_16X8

.subckt SP6TVar17Array_4X1 vss vdd wl[0] wl[1] wl[2] wl[3] bl[0] bl_n[0]
Xinst0x0 vss vdd wl[0] wl[1] bl[0] bl_n[0] SP6TVar17Array_2X1
Xinst1x0 vss vdd wl[2] wl[3] bl[0] bl_n[0] SP6TVar17Array_2X1
.ends SP6TVar17Array_4X1

.subckt SP6TVar17Array_8X1 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] bl[0] bl_n[0] SP6TVar17Array_4X1
Xinst1x0 vss vdd wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] SP6TVar17Array_4X1
.ends SP6TVar17Array_8X1

.subckt SP6TVar17Array_16X1BC vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] bl[0] bl_n[0]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] SP6TVar17Array_8X1
Xinst1x0 vss vdd wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] bl[0] bl_n[0] SP6TVar17Array_8X1
Xbottombcrow vdd vss bl[0] bl_n[0] SP6TVar17BulkConn
Xtopbcrow vdd vss bl[0] bl_n[0] SP6TVar17BulkConn
.ends SP6TVar17Array_16X1BC

.subckt SP6TVar17Array_8X2 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar17Array_4X2
Xinst1x0 vss vdd wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar17Array_4X2
.ends SP6TVar17Array_8X2

.subckt SP6TVar17Array_16X2BC vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] bl[0] bl_n[0] bl[1] bl_n[1]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar17Array_8X2
Xinst1x0 vss vdd wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar17Array_8X2
Xbottombcrow vss vdd bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar17BulkConnRow_2
Xtopbcrow vss vdd bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar17BulkConnRow_2
.ends SP6TVar17Array_16X2BC

.subckt SP6TVar17Array_16X4BC vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar17Array_8X4
Xinst1x0 vss vdd wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar17Array_8X4
Xbottombcrow vss vdd bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar17BulkConnRow_4
Xtopbcrow vss vdd bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar17BulkConnRow_4
.ends SP6TVar17Array_16X4BC

.subckt SP6TVar17Array_6X1 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] bl[0] bl_n[0]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] bl[0] bl_n[0] SP6TVar17Array_4X1
Xinst1x0 vss vdd wl[4] wl[5] bl[0] bl_n[0] SP6TVar17Array_2X1
.ends SP6TVar17Array_6X1

.subckt SP6TVar17CellConnectOut wl bl bl_n vdd vss bit bit_n
Xpu1 vdd bit_n bit vdd sg13_lv_pmos l=1.3e-07 w=2e-07
Xpd1 bit bit_n vss vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpu2 vdd bit bit_n vdd sg13_lv_pmos l=1.3e-07 w=2e-07
Xpd2 bit_n bit vss vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg1 bit wl bl vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg2 bit_n wl bl_n vss sg13_lv_nmos l=1.3e-07 w=2e-07
.ends SP6TVar17CellConnectOut

.subckt SP6TVar17TestArray_16X8C vss vdd bl bl_n bit bit_n wl
Xarray_0 vss vdd zero zero zero zero zero zero zero zero wl zero zero zero zero zero zero zero array_0_bl[0] array_0_bl_n[0] SP6TVar17Array_16X1BC
Xarray_1 vss vdd zero zero zero zero zero zero zero zero wl zero zero zero zero zero zero zero array_1_bl[0] array_1_bl_n[0] array_1_bl[1] array_1_bl_n[1] SP6TVar17Array_16X2BC
Xarray_2 vss vdd zero zero zero zero zero zero zero zero wl zero zero zero zero zero zero zero array_2_bl[0] array_2_bl_n[0] array_2_bl[1] array_2_bl_n[1] array_2_bl[2] array_2_bl_n[2] array_2_bl[3] array_2_bl_n[3] SP6TVar17Array_16X4BC
Xcolbc_0 vdd vss bl bl_n SP6TVar17BulkConn
Xcolbc_1 vdd vss bl bl_n SP6TVar17BulkConn
Xcolarray_0 vss vdd zero zero zero zero zero zero zero zero bl bl_n SP6TVar17Array_8X1
Xcolarray_1 vss vdd zero zero zero zero zero zero bl bl_n SP6TVar17Array_6X1
Xbc_noconn zero bl bl_n vdd vss SP6TVar17Cell
Xbc_conn wl bl bl_n vdd vss bit bit_n SP6TVar17CellConnectOut
Xzero vdd vss zero zero_x1
.ends SP6TVar17TestArray_16X8C

.subckt SP6TVar17 vss noco_vdd noco_wl noco_bl noco_bl_n co_vdd co_bl co_bl_n co_bit co_bit_n co_wl
Xframe noco_vdd noco_wl NoConn_PAD0x2 co_vdd co_bl_n co_bit co_bit_n NoConn_PAD0x7 NoConn_PAD0x8 NoConn_PAD0x9 vss noco_bl noco_bl_n vss co_bl co_wl NoConn_PAD1x6 NoConn_PAD1x7 NoConn_PAD1x8 NoConn_PAD1x9 PadFrame_SP17
Xtestarray_noco vss noco_vdd noco_bl noco_bl_n noco_wl SP6TVar17TestArray_16X8
Xtestarray_co vss co_vdd co_bl co_bl_n co_bit co_bit_n co_wl SP6TVar17TestArray_16X8C
.ends SP6TVar17

.subckt PadFrame_SP18 PAD0x0 PAD0x1 PAD0x2 PAD0x3 PAD0x4 PAD0x5 PAD0x6 PAD0x7 PAD0x8 PAD0x9 PAD1x0 PAD1x1 PAD1x2 PAD1x3 PAD1x4 PAD1x5 PAD1x6 PAD1x7 PAD1x8 PAD1x9
XPAD0x0 PAD0x0 BondPad
XPAD0x1 PAD0x1 BondPad
XPAD0x2 PAD0x2 BondPad
XPAD0x3 PAD0x3 BondPad
XPAD0x4 PAD0x4 BondPad
XPAD0x5 PAD0x5 BondPad
XPAD0x6 PAD0x6 BondPad
XPAD0x7 PAD0x7 BondPad
XPAD0x8 PAD0x8 BondPad
XPAD0x9 PAD0x9 BondPad
XPAD1x0 PAD1x0 BondPad
XPAD1x1 PAD1x1 BondPad
XPAD1x2 PAD1x2 BondPad
XPAD1x3 PAD1x3 BondPad
XPAD1x4 PAD1x4 BondPad
XPAD1x5 PAD1x5 BondPad
XPAD1x6 PAD1x6 BondPad
XPAD1x7 PAD1x7 BondPad
XPAD1x8 PAD1x8 BondPad
XPAD1x9 PAD1x9 BondPad
.ends PadFrame_SP18

.subckt SP6TVar18Cell wl bl bl_n vdd vss
Xpu1 vdd bit_n bit vdd sg13_lv_pmos l=1.3e-07 w=1.5e-07
Xpd1 bit bit_n vss vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpu2 vdd bit bit_n vdd sg13_lv_pmos l=1.3e-07 w=1.5e-07
Xpd2 bit_n bit vss vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg1 bit wl bl vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg2 bit_n wl bl_n vss sg13_lv_nmos l=1.3e-07 w=2e-07
.ends SP6TVar18Cell

.subckt SP6TVar18Array_2X1 vss vdd wl[0] wl[1] bl[0] bl_n[0]
Xinst0x0 wl[0] bl[0] bl_n[0] vdd vss SP6TVar18Cell
Xinst1x0 wl[1] bl[0] bl_n[0] vdd vss SP6TVar18Cell
.ends SP6TVar18Array_2X1

.subckt SP6TVar18Array_2X2 vss vdd wl[0] wl[1] bl[0] bl_n[0] bl[1] bl_n[1]
Xinst0x0 vss vdd wl[0] wl[1] bl[0] bl_n[0] SP6TVar18Array_2X1
Xinst0x1 vss vdd wl[0] wl[1] bl[1] bl_n[1] SP6TVar18Array_2X1
.ends SP6TVar18Array_2X2

.subckt SP6TVar18Array_4X2 vss vdd wl[0] wl[1] wl[2] wl[3] bl[0] bl_n[0] bl[1] bl_n[1]
Xinst0x0 vss vdd wl[0] wl[1] bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar18Array_2X2
Xinst1x0 vss vdd wl[2] wl[3] bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar18Array_2X2
.ends SP6TVar18Array_4X2

.subckt SP6TVar18Array_4X4 vss vdd wl[0] wl[1] wl[2] wl[3] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar18Array_4X2
Xinst0x1 vss vdd wl[0] wl[1] wl[2] wl[3] bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar18Array_4X2
.ends SP6TVar18Array_4X4

.subckt SP6TVar18Array_8X4 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar18Array_4X4
Xinst1x0 vss vdd wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar18Array_4X4
.ends SP6TVar18Array_8X4

.subckt SP6TVar18Array_8X8 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar18Array_8X4
Xinst0x1 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7] SP6TVar18Array_8X4
.ends SP6TVar18Array_8X8

.subckt SP6TVar18BulkConn vdd vss bl bl_n
.ends SP6TVar18BulkConn

.subckt SP6TVar18BulkConnRow_2 vss vdd bl[0] bl_n[0] bl[1] bl_n[1]
Xinst0 vdd vss bl[0] bl_n[0] SP6TVar18BulkConn
Xinst1 vdd vss bl[1] bl_n[1] SP6TVar18BulkConn
.ends SP6TVar18BulkConnRow_2

.subckt SP6TVar18BulkConnRow_4 vss vdd bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3]
Xinst0 vss vdd bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar18BulkConnRow_2
Xinst1 vss vdd bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar18BulkConnRow_2
.ends SP6TVar18BulkConnRow_4

.subckt SP6TVar18BulkConnRow_8 vss vdd bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7]
Xinst0 vss vdd bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar18BulkConnRow_4
Xinst1 vss vdd bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7] SP6TVar18BulkConnRow_4
.ends SP6TVar18BulkConnRow_8

.subckt SP6TVar18Array_16X8BC vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7] SP6TVar18Array_8X8
Xinst1x0 vss vdd wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7] SP6TVar18Array_8X8
Xbottombcrow vss vdd bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7] SP6TVar18BulkConnRow_8
Xtopbcrow vss vdd bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7] SP6TVar18BulkConnRow_8
.ends SP6TVar18Array_16X8BC

.subckt SP6TVar18TestArray_16X8 vss vdd bl bl_n wl
Xarray vss vdd zero zero zero zero zero zero zero zero wl zero zero zero zero zero zero zero bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl bl_n bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7] SP6TVar18Array_16X8BC
Xzero vdd vss zero zero_x1
.ends SP6TVar18TestArray_16X8

.subckt SP6TVar18Array_4X1 vss vdd wl[0] wl[1] wl[2] wl[3] bl[0] bl_n[0]
Xinst0x0 vss vdd wl[0] wl[1] bl[0] bl_n[0] SP6TVar18Array_2X1
Xinst1x0 vss vdd wl[2] wl[3] bl[0] bl_n[0] SP6TVar18Array_2X1
.ends SP6TVar18Array_4X1

.subckt SP6TVar18Array_8X1 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] bl[0] bl_n[0] SP6TVar18Array_4X1
Xinst1x0 vss vdd wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] SP6TVar18Array_4X1
.ends SP6TVar18Array_8X1

.subckt SP6TVar18Array_16X1BC vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] bl[0] bl_n[0]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] SP6TVar18Array_8X1
Xinst1x0 vss vdd wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] bl[0] bl_n[0] SP6TVar18Array_8X1
Xbottombcrow vdd vss bl[0] bl_n[0] SP6TVar18BulkConn
Xtopbcrow vdd vss bl[0] bl_n[0] SP6TVar18BulkConn
.ends SP6TVar18Array_16X1BC

.subckt SP6TVar18Array_8X2 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar18Array_4X2
Xinst1x0 vss vdd wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar18Array_4X2
.ends SP6TVar18Array_8X2

.subckt SP6TVar18Array_16X2BC vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] bl[0] bl_n[0] bl[1] bl_n[1]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar18Array_8X2
Xinst1x0 vss vdd wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar18Array_8X2
Xbottombcrow vss vdd bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar18BulkConnRow_2
Xtopbcrow vss vdd bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar18BulkConnRow_2
.ends SP6TVar18Array_16X2BC

.subckt SP6TVar18Array_16X4BC vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar18Array_8X4
Xinst1x0 vss vdd wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar18Array_8X4
Xbottombcrow vss vdd bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar18BulkConnRow_4
Xtopbcrow vss vdd bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar18BulkConnRow_4
.ends SP6TVar18Array_16X4BC

.subckt SP6TVar18Array_6X1 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] bl[0] bl_n[0]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] bl[0] bl_n[0] SP6TVar18Array_4X1
Xinst1x0 vss vdd wl[4] wl[5] bl[0] bl_n[0] SP6TVar18Array_2X1
.ends SP6TVar18Array_6X1

.subckt SP6TVar18CellConnectOut wl bl bl_n vdd vss bit bit_n
Xpu1 vdd bit_n bit vdd sg13_lv_pmos l=1.3e-07 w=1.5e-07
Xpd1 bit bit_n vss vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpu2 vdd bit bit_n vdd sg13_lv_pmos l=1.3e-07 w=1.5e-07
Xpd2 bit_n bit vss vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg1 bit wl bl vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg2 bit_n wl bl_n vss sg13_lv_nmos l=1.3e-07 w=2e-07
.ends SP6TVar18CellConnectOut

.subckt SP6TVar18TestArray_16X8C vss vdd bl bl_n bit bit_n wl
Xarray_0 vss vdd zero zero zero zero zero zero zero zero wl zero zero zero zero zero zero zero array_0_bl[0] array_0_bl_n[0] SP6TVar18Array_16X1BC
Xarray_1 vss vdd zero zero zero zero zero zero zero zero wl zero zero zero zero zero zero zero array_1_bl[0] array_1_bl_n[0] array_1_bl[1] array_1_bl_n[1] SP6TVar18Array_16X2BC
Xarray_2 vss vdd zero zero zero zero zero zero zero zero wl zero zero zero zero zero zero zero array_2_bl[0] array_2_bl_n[0] array_2_bl[1] array_2_bl_n[1] array_2_bl[2] array_2_bl_n[2] array_2_bl[3] array_2_bl_n[3] SP6TVar18Array_16X4BC
Xcolbc_0 vdd vss bl bl_n SP6TVar18BulkConn
Xcolbc_1 vdd vss bl bl_n SP6TVar18BulkConn
Xcolarray_0 vss vdd zero zero zero zero zero zero zero zero bl bl_n SP6TVar18Array_8X1
Xcolarray_1 vss vdd zero zero zero zero zero zero bl bl_n SP6TVar18Array_6X1
Xbc_noconn zero bl bl_n vdd vss SP6TVar18Cell
Xbc_conn wl bl bl_n vdd vss bit bit_n SP6TVar18CellConnectOut
Xzero vdd vss zero zero_x1
.ends SP6TVar18TestArray_16X8C

.subckt SP6TVar18 vss noco_vdd noco_wl noco_bl noco_bl_n co_vdd co_bl co_bl_n co_bit co_bit_n co_wl
Xframe noco_vdd noco_wl NoConn_PAD0x2 co_vdd co_bl_n co_bit co_bit_n NoConn_PAD0x7 NoConn_PAD0x8 NoConn_PAD0x9 vss noco_bl noco_bl_n vss co_bl co_wl NoConn_PAD1x6 NoConn_PAD1x7 NoConn_PAD1x8 NoConn_PAD1x9 PadFrame_SP18
Xtestarray_noco vss noco_vdd noco_bl noco_bl_n noco_wl SP6TVar18TestArray_16X8
Xtestarray_co vss co_vdd co_bl co_bl_n co_bit co_bit_n co_wl SP6TVar18TestArray_16X8C
.ends SP6TVar18

.subckt PadFrame_SP19 PAD0x0 PAD0x1 PAD0x2 PAD0x3 PAD0x4 PAD0x5 PAD0x6 PAD0x7 PAD0x8 PAD0x9 PAD1x0 PAD1x1 PAD1x2 PAD1x3 PAD1x4 PAD1x5 PAD1x6 PAD1x7 PAD1x8 PAD1x9
XPAD0x0 PAD0x0 BondPad
XPAD0x1 PAD0x1 BondPad
XPAD0x2 PAD0x2 BondPad
XPAD0x3 PAD0x3 BondPad
XPAD0x4 PAD0x4 BondPad
XPAD0x5 PAD0x5 BondPad
XPAD0x6 PAD0x6 BondPad
XPAD0x7 PAD0x7 BondPad
XPAD0x8 PAD0x8 BondPad
XPAD0x9 PAD0x9 BondPad
XPAD1x0 PAD1x0 BondPad
XPAD1x1 PAD1x1 BondPad
XPAD1x2 PAD1x2 BondPad
XPAD1x3 PAD1x3 BondPad
XPAD1x4 PAD1x4 BondPad
XPAD1x5 PAD1x5 BondPad
XPAD1x6 PAD1x6 BondPad
XPAD1x7 PAD1x7 BondPad
XPAD1x8 PAD1x8 BondPad
XPAD1x9 PAD1x9 BondPad
.ends PadFrame_SP19

.subckt SP6TVar19Cell wl bl bl_n vdd vss
Xpu1 vdd bit_n bit vdd sg13_lv_pmos l=1.3e-07 w=2e-07
Xpd1 bit bit_n vss vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpu2 vdd bit bit_n vdd sg13_lv_pmos l=1.3e-07 w=2e-07
Xpd2 bit_n bit vss vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg1 bit wl bl vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg2 bit_n wl bl_n vss sg13_lv_nmos l=1.3e-07 w=2e-07
.ends SP6TVar19Cell

.subckt SP6TVar19Array_2X1 vss vdd wl[0] wl[1] bl[0] bl_n[0]
Xinst0x0 wl[0] bl[0] bl_n[0] vdd vss SP6TVar19Cell
Xinst1x0 wl[1] bl[0] bl_n[0] vdd vss SP6TVar19Cell
.ends SP6TVar19Array_2X1

.subckt SP6TVar19Array_2X2 vss vdd wl[0] wl[1] bl[0] bl_n[0] bl[1] bl_n[1]
Xinst0x0 vss vdd wl[0] wl[1] bl[0] bl_n[0] SP6TVar19Array_2X1
Xinst0x1 vss vdd wl[0] wl[1] bl[1] bl_n[1] SP6TVar19Array_2X1
.ends SP6TVar19Array_2X2

.subckt SP6TVar19Array_4X2 vss vdd wl[0] wl[1] wl[2] wl[3] bl[0] bl_n[0] bl[1] bl_n[1]
Xinst0x0 vss vdd wl[0] wl[1] bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar19Array_2X2
Xinst1x0 vss vdd wl[2] wl[3] bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar19Array_2X2
.ends SP6TVar19Array_4X2

.subckt SP6TVar19Array_4X4 vss vdd wl[0] wl[1] wl[2] wl[3] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar19Array_4X2
Xinst0x1 vss vdd wl[0] wl[1] wl[2] wl[3] bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar19Array_4X2
.ends SP6TVar19Array_4X4

.subckt SP6TVar19Array_8X4 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar19Array_4X4
Xinst1x0 vss vdd wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar19Array_4X4
.ends SP6TVar19Array_8X4

.subckt SP6TVar19Array_8X8 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar19Array_8X4
Xinst0x1 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7] SP6TVar19Array_8X4
.ends SP6TVar19Array_8X8

.subckt SP6TVar19BulkConn vdd vss bl bl_n
.ends SP6TVar19BulkConn

.subckt SP6TVar19BulkConnRow_2 vss vdd bl[0] bl_n[0] bl[1] bl_n[1]
Xinst0 vdd vss bl[0] bl_n[0] SP6TVar19BulkConn
Xinst1 vdd vss bl[1] bl_n[1] SP6TVar19BulkConn
.ends SP6TVar19BulkConnRow_2

.subckt SP6TVar19BulkConnRow_4 vss vdd bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3]
Xinst0 vss vdd bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar19BulkConnRow_2
Xinst1 vss vdd bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar19BulkConnRow_2
.ends SP6TVar19BulkConnRow_4

.subckt SP6TVar19BulkConnRow_8 vss vdd bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7]
Xinst0 vss vdd bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar19BulkConnRow_4
Xinst1 vss vdd bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7] SP6TVar19BulkConnRow_4
.ends SP6TVar19BulkConnRow_8

.subckt SP6TVar19Array_16X8BC vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7] SP6TVar19Array_8X8
Xinst1x0 vss vdd wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7] SP6TVar19Array_8X8
Xbottombcrow vss vdd bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7] SP6TVar19BulkConnRow_8
Xtopbcrow vss vdd bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7] SP6TVar19BulkConnRow_8
.ends SP6TVar19Array_16X8BC

.subckt SP6TVar19TestArray_16X8 vss vdd bl bl_n wl
Xarray vss vdd zero zero zero zero zero zero zero zero wl zero zero zero zero zero zero zero bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl bl_n bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7] SP6TVar19Array_16X8BC
Xzero vdd vss zero zero_x1
.ends SP6TVar19TestArray_16X8

.subckt SP6TVar19Array_4X1 vss vdd wl[0] wl[1] wl[2] wl[3] bl[0] bl_n[0]
Xinst0x0 vss vdd wl[0] wl[1] bl[0] bl_n[0] SP6TVar19Array_2X1
Xinst1x0 vss vdd wl[2] wl[3] bl[0] bl_n[0] SP6TVar19Array_2X1
.ends SP6TVar19Array_4X1

.subckt SP6TVar19Array_8X1 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] bl[0] bl_n[0] SP6TVar19Array_4X1
Xinst1x0 vss vdd wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] SP6TVar19Array_4X1
.ends SP6TVar19Array_8X1

.subckt SP6TVar19Array_16X1BC vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] bl[0] bl_n[0]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] SP6TVar19Array_8X1
Xinst1x0 vss vdd wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] bl[0] bl_n[0] SP6TVar19Array_8X1
Xbottombcrow vdd vss bl[0] bl_n[0] SP6TVar19BulkConn
Xtopbcrow vdd vss bl[0] bl_n[0] SP6TVar19BulkConn
.ends SP6TVar19Array_16X1BC

.subckt SP6TVar19Array_8X2 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar19Array_4X2
Xinst1x0 vss vdd wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar19Array_4X2
.ends SP6TVar19Array_8X2

.subckt SP6TVar19Array_16X2BC vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] bl[0] bl_n[0] bl[1] bl_n[1]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar19Array_8X2
Xinst1x0 vss vdd wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar19Array_8X2
Xbottombcrow vss vdd bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar19BulkConnRow_2
Xtopbcrow vss vdd bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar19BulkConnRow_2
.ends SP6TVar19Array_16X2BC

.subckt SP6TVar19Array_16X4BC vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar19Array_8X4
Xinst1x0 vss vdd wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar19Array_8X4
Xbottombcrow vss vdd bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar19BulkConnRow_4
Xtopbcrow vss vdd bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar19BulkConnRow_4
.ends SP6TVar19Array_16X4BC

.subckt SP6TVar19Array_6X1 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] bl[0] bl_n[0]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] bl[0] bl_n[0] SP6TVar19Array_4X1
Xinst1x0 vss vdd wl[4] wl[5] bl[0] bl_n[0] SP6TVar19Array_2X1
.ends SP6TVar19Array_6X1

.subckt SP6TVar19CellConnectOut wl bl bl_n vdd vss bit bit_n
Xpu1 vdd bit_n bit vdd sg13_lv_pmos l=1.3e-07 w=2e-07
Xpd1 bit bit_n vss vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpu2 vdd bit bit_n vdd sg13_lv_pmos l=1.3e-07 w=2e-07
Xpd2 bit_n bit vss vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg1 bit wl bl vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg2 bit_n wl bl_n vss sg13_lv_nmos l=1.3e-07 w=2e-07
.ends SP6TVar19CellConnectOut

.subckt SP6TVar19TestArray_16X8C vss vdd bl bl_n bit bit_n wl
Xarray_0 vss vdd zero zero zero zero zero zero zero zero wl zero zero zero zero zero zero zero array_0_bl[0] array_0_bl_n[0] SP6TVar19Array_16X1BC
Xarray_1 vss vdd zero zero zero zero zero zero zero zero wl zero zero zero zero zero zero zero array_1_bl[0] array_1_bl_n[0] array_1_bl[1] array_1_bl_n[1] SP6TVar19Array_16X2BC
Xarray_2 vss vdd zero zero zero zero zero zero zero zero wl zero zero zero zero zero zero zero array_2_bl[0] array_2_bl_n[0] array_2_bl[1] array_2_bl_n[1] array_2_bl[2] array_2_bl_n[2] array_2_bl[3] array_2_bl_n[3] SP6TVar19Array_16X4BC
Xcolbc_0 vdd vss bl bl_n SP6TVar19BulkConn
Xcolbc_1 vdd vss bl bl_n SP6TVar19BulkConn
Xcolarray_0 vss vdd zero zero zero zero zero zero zero zero bl bl_n SP6TVar19Array_8X1
Xcolarray_1 vss vdd zero zero zero zero zero zero bl bl_n SP6TVar19Array_6X1
Xbc_noconn zero bl bl_n vdd vss SP6TVar19Cell
Xbc_conn wl bl bl_n vdd vss bit bit_n SP6TVar19CellConnectOut
Xzero vdd vss zero zero_x1
.ends SP6TVar19TestArray_16X8C

.subckt SP6TVar19 vss noco_vdd noco_wl noco_bl noco_bl_n co_vdd co_bl co_bl_n co_bit co_bit_n co_wl
Xframe noco_vdd noco_wl NoConn_PAD0x2 co_vdd co_bl_n co_bit co_bit_n NoConn_PAD0x7 NoConn_PAD0x8 NoConn_PAD0x9 vss noco_bl noco_bl_n vss co_bl co_wl NoConn_PAD1x6 NoConn_PAD1x7 NoConn_PAD1x8 NoConn_PAD1x9 PadFrame_SP19
Xtestarray_noco vss noco_vdd noco_bl noco_bl_n noco_wl SP6TVar19TestArray_16X8
Xtestarray_co vss co_vdd co_bl co_bl_n co_bit co_bit_n co_wl SP6TVar19TestArray_16X8C
.ends SP6TVar19

.subckt PadFrame_SP20 PAD0x0 PAD0x1 PAD0x2 PAD0x3 PAD0x4 PAD0x5 PAD0x6 PAD0x7 PAD0x8 PAD0x9 PAD1x0 PAD1x1 PAD1x2 PAD1x3 PAD1x4 PAD1x5 PAD1x6 PAD1x7 PAD1x8 PAD1x9
XPAD0x0 PAD0x0 BondPad
XPAD0x1 PAD0x1 BondPad
XPAD0x2 PAD0x2 BondPad
XPAD0x3 PAD0x3 BondPad
XPAD0x4 PAD0x4 BondPad
XPAD0x5 PAD0x5 BondPad
XPAD0x6 PAD0x6 BondPad
XPAD0x7 PAD0x7 BondPad
XPAD0x8 PAD0x8 BondPad
XPAD0x9 PAD0x9 BondPad
XPAD1x0 PAD1x0 BondPad
XPAD1x1 PAD1x1 BondPad
XPAD1x2 PAD1x2 BondPad
XPAD1x3 PAD1x3 BondPad
XPAD1x4 PAD1x4 BondPad
XPAD1x5 PAD1x5 BondPad
XPAD1x6 PAD1x6 BondPad
XPAD1x7 PAD1x7 BondPad
XPAD1x8 PAD1x8 BondPad
XPAD1x9 PAD1x9 BondPad
.ends PadFrame_SP20

.subckt SP6TVar20Cell wl bl bl_n vdd vss
Xpu1 vdd bit_n bit vdd sg13_lv_pmos l=1.3e-07 w=1.5e-07
Xpd1 bit bit_n vss vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpu2 vdd bit bit_n vdd sg13_lv_pmos l=1.3e-07 w=1.5e-07
Xpd2 bit_n bit vss vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg1 bit wl bl vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg2 bit_n wl bl_n vss sg13_lv_nmos l=1.3e-07 w=2e-07
.ends SP6TVar20Cell

.subckt SP6TVar20Array_2X1 vss vdd wl[0] wl[1] bl[0] bl_n[0]
Xinst0x0 wl[0] bl[0] bl_n[0] vdd vss SP6TVar20Cell
Xinst1x0 wl[1] bl[0] bl_n[0] vdd vss SP6TVar20Cell
.ends SP6TVar20Array_2X1

.subckt SP6TVar20Array_2X2 vss vdd wl[0] wl[1] bl[0] bl_n[0] bl[1] bl_n[1]
Xinst0x0 vss vdd wl[0] wl[1] bl[0] bl_n[0] SP6TVar20Array_2X1
Xinst0x1 vss vdd wl[0] wl[1] bl[1] bl_n[1] SP6TVar20Array_2X1
.ends SP6TVar20Array_2X2

.subckt SP6TVar20Array_4X2 vss vdd wl[0] wl[1] wl[2] wl[3] bl[0] bl_n[0] bl[1] bl_n[1]
Xinst0x0 vss vdd wl[0] wl[1] bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar20Array_2X2
Xinst1x0 vss vdd wl[2] wl[3] bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar20Array_2X2
.ends SP6TVar20Array_4X2

.subckt SP6TVar20Array_4X4 vss vdd wl[0] wl[1] wl[2] wl[3] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar20Array_4X2
Xinst0x1 vss vdd wl[0] wl[1] wl[2] wl[3] bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar20Array_4X2
.ends SP6TVar20Array_4X4

.subckt SP6TVar20Array_8X4 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar20Array_4X4
Xinst1x0 vss vdd wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar20Array_4X4
.ends SP6TVar20Array_8X4

.subckt SP6TVar20Array_8X8 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar20Array_8X4
Xinst0x1 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7] SP6TVar20Array_8X4
.ends SP6TVar20Array_8X8

.subckt SP6TVar20BulkConn vdd vss bl bl_n
.ends SP6TVar20BulkConn

.subckt SP6TVar20BulkConnRow_2 vss vdd bl[0] bl_n[0] bl[1] bl_n[1]
Xinst0 vdd vss bl[0] bl_n[0] SP6TVar20BulkConn
Xinst1 vdd vss bl[1] bl_n[1] SP6TVar20BulkConn
.ends SP6TVar20BulkConnRow_2

.subckt SP6TVar20BulkConnRow_4 vss vdd bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3]
Xinst0 vss vdd bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar20BulkConnRow_2
Xinst1 vss vdd bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar20BulkConnRow_2
.ends SP6TVar20BulkConnRow_4

.subckt SP6TVar20BulkConnRow_8 vss vdd bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7]
Xinst0 vss vdd bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar20BulkConnRow_4
Xinst1 vss vdd bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7] SP6TVar20BulkConnRow_4
.ends SP6TVar20BulkConnRow_8

.subckt SP6TVar20Array_16X8BC vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7] SP6TVar20Array_8X8
Xinst1x0 vss vdd wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7] SP6TVar20Array_8X8
Xbottombcrow vss vdd bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7] SP6TVar20BulkConnRow_8
Xtopbcrow vss vdd bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7] SP6TVar20BulkConnRow_8
.ends SP6TVar20Array_16X8BC

.subckt SP6TVar20TestArray_16X8 vss vdd bl bl_n wl
Xarray vss vdd zero zero zero zero zero zero zero zero wl zero zero zero zero zero zero zero bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl bl_n bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7] SP6TVar20Array_16X8BC
Xzero vdd vss zero zero_x1
.ends SP6TVar20TestArray_16X8

.subckt SP6TVar20Array_4X1 vss vdd wl[0] wl[1] wl[2] wl[3] bl[0] bl_n[0]
Xinst0x0 vss vdd wl[0] wl[1] bl[0] bl_n[0] SP6TVar20Array_2X1
Xinst1x0 vss vdd wl[2] wl[3] bl[0] bl_n[0] SP6TVar20Array_2X1
.ends SP6TVar20Array_4X1

.subckt SP6TVar20Array_8X1 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] bl[0] bl_n[0] SP6TVar20Array_4X1
Xinst1x0 vss vdd wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] SP6TVar20Array_4X1
.ends SP6TVar20Array_8X1

.subckt SP6TVar20Array_16X1BC vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] bl[0] bl_n[0]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] SP6TVar20Array_8X1
Xinst1x0 vss vdd wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] bl[0] bl_n[0] SP6TVar20Array_8X1
Xbottombcrow vdd vss bl[0] bl_n[0] SP6TVar20BulkConn
Xtopbcrow vdd vss bl[0] bl_n[0] SP6TVar20BulkConn
.ends SP6TVar20Array_16X1BC

.subckt SP6TVar20Array_8X2 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar20Array_4X2
Xinst1x0 vss vdd wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar20Array_4X2
.ends SP6TVar20Array_8X2

.subckt SP6TVar20Array_16X2BC vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] bl[0] bl_n[0] bl[1] bl_n[1]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar20Array_8X2
Xinst1x0 vss vdd wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar20Array_8X2
Xbottombcrow vss vdd bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar20BulkConnRow_2
Xtopbcrow vss vdd bl[0] bl_n[0] bl[1] bl_n[1] SP6TVar20BulkConnRow_2
.ends SP6TVar20Array_16X2BC

.subckt SP6TVar20Array_16X4BC vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar20Array_8X4
Xinst1x0 vss vdd wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar20Array_8X4
Xbottombcrow vss vdd bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar20BulkConnRow_4
Xtopbcrow vss vdd bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] SP6TVar20BulkConnRow_4
.ends SP6TVar20Array_16X4BC

.subckt SP6TVar20Array_6X1 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] bl[0] bl_n[0]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] bl[0] bl_n[0] SP6TVar20Array_4X1
Xinst1x0 vss vdd wl[4] wl[5] bl[0] bl_n[0] SP6TVar20Array_2X1
.ends SP6TVar20Array_6X1

.subckt SP6TVar20CellConnectOut wl bl bl_n vdd vss bit bit_n
Xpu1 vdd bit_n bit vdd sg13_lv_pmos l=1.3e-07 w=1.5e-07
Xpd1 bit bit_n vss vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpu2 vdd bit bit_n vdd sg13_lv_pmos l=1.3e-07 w=1.5e-07
Xpd2 bit_n bit vss vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg1 bit wl bl vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg2 bit_n wl bl_n vss sg13_lv_nmos l=1.3e-07 w=2e-07
.ends SP6TVar20CellConnectOut

.subckt SP6TVar20TestArray_16X8C vss vdd bl bl_n bit bit_n wl
Xarray_0 vss vdd zero zero zero zero zero zero zero zero wl zero zero zero zero zero zero zero array_0_bl[0] array_0_bl_n[0] SP6TVar20Array_16X1BC
Xarray_1 vss vdd zero zero zero zero zero zero zero zero wl zero zero zero zero zero zero zero array_1_bl[0] array_1_bl_n[0] array_1_bl[1] array_1_bl_n[1] SP6TVar20Array_16X2BC
Xarray_2 vss vdd zero zero zero zero zero zero zero zero wl zero zero zero zero zero zero zero array_2_bl[0] array_2_bl_n[0] array_2_bl[1] array_2_bl_n[1] array_2_bl[2] array_2_bl_n[2] array_2_bl[3] array_2_bl_n[3] SP6TVar20Array_16X4BC
Xcolbc_0 vdd vss bl bl_n SP6TVar20BulkConn
Xcolbc_1 vdd vss bl bl_n SP6TVar20BulkConn
Xcolarray_0 vss vdd zero zero zero zero zero zero zero zero bl bl_n SP6TVar20Array_8X1
Xcolarray_1 vss vdd zero zero zero zero zero zero bl bl_n SP6TVar20Array_6X1
Xbc_noconn zero bl bl_n vdd vss SP6TVar20Cell
Xbc_conn wl bl bl_n vdd vss bit bit_n SP6TVar20CellConnectOut
Xzero vdd vss zero zero_x1
.ends SP6TVar20TestArray_16X8C

.subckt SP6TVar20 vss noco_vdd noco_wl noco_bl noco_bl_n co_vdd co_bl co_bl_n co_bit co_bit_n co_wl
Xframe noco_vdd noco_wl NoConn_PAD0x2 co_vdd co_bl_n co_bit co_bit_n NoConn_PAD0x7 NoConn_PAD0x8 NoConn_PAD0x9 vss noco_bl noco_bl_n vss co_bl co_wl NoConn_PAD1x6 NoConn_PAD1x7 NoConn_PAD1x8 NoConn_PAD1x9 PadFrame_SP20
Xtestarray_noco vss noco_vdd noco_bl noco_bl_n noco_wl SP6TVar20TestArray_16X8
Xtestarray_co vss co_vdd co_bl co_bl_n co_bit co_bit_n co_wl SP6TVar20TestArray_16X8C
.ends SP6TVar20

.subckt PadFrame_SP21 PAD0x0 PAD0x1 PAD0x2 PAD0x3 PAD0x4 PAD0x5 PAD0x6 PAD0x7 PAD0x8 PAD0x9 PAD1x0 PAD1x1 PAD1x2 PAD1x3 PAD1x4 PAD1x5 PAD1x6 PAD1x7 PAD1x8 PAD1x9
XPAD0x0 PAD0x0 BondPad
XPAD0x1 PAD0x1 BondPad
XPAD0x2 PAD0x2 BondPad
XPAD0x3 PAD0x3 BondPad
XPAD0x4 PAD0x4 BondPad
XPAD0x5 PAD0x5 BondPad
XPAD0x6 PAD0x6 BondPad
XPAD0x7 PAD0x7 BondPad
XPAD0x8 PAD0x8 BondPad
XPAD0x9 PAD0x9 BondPad
XPAD1x0 PAD1x0 BondPad
XPAD1x1 PAD1x1 BondPad
XPAD1x2 PAD1x2 BondPad
XPAD1x3 PAD1x3 BondPad
XPAD1x4 PAD1x4 BondPad
XPAD1x5 PAD1x5 BondPad
XPAD1x6 PAD1x6 BondPad
XPAD1x7 PAD1x7 BondPad
XPAD1x8 PAD1x8 BondPad
XPAD1x9 PAD1x9 BondPad
.ends PadFrame_SP21

.subckt OldSP6TCell wl bl bl_n vdd vss
Xpu1 vdd bit_n bit vdd sg13_lv_pmos l=1.3e-07 w=1.5e-07
Xpd1 bit bit_n vss vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpu2 vdd bit bit_n vdd sg13_lv_pmos l=1.3e-07 w=1.5e-07
Xpd2 bit_n bit vss vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg1 bit wl bl vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg2 bit_n wl bl_n vss sg13_lv_nmos l=1.3e-07 w=3e-07
.ends OldSP6TCell

.subckt OldSP6TArray_2X1 vss vdd wl[0] wl[1] bl[0] bl_n[0]
Xinst0x0 wl[0] bl[0] bl_n[0] vdd vss OldSP6TCell
Xinst1x0 wl[1] bl[0] bl_n[0] vdd vss OldSP6TCell
.ends OldSP6TArray_2X1

.subckt OldSP6TArray_2X2 vss vdd wl[0] wl[1] bl[0] bl_n[0] bl[1] bl_n[1]
Xinst0x0 vss vdd wl[0] wl[1] bl[0] bl_n[0] OldSP6TArray_2X1
Xinst0x1 vss vdd wl[0] wl[1] bl[1] bl_n[1] OldSP6TArray_2X1
.ends OldSP6TArray_2X2

.subckt OldSP6TArray_4X2 vss vdd wl[0] wl[1] wl[2] wl[3] bl[0] bl_n[0] bl[1] bl_n[1]
Xinst0x0 vss vdd wl[0] wl[1] bl[0] bl_n[0] bl[1] bl_n[1] OldSP6TArray_2X2
Xinst1x0 vss vdd wl[2] wl[3] bl[0] bl_n[0] bl[1] bl_n[1] OldSP6TArray_2X2
.ends OldSP6TArray_4X2

.subckt OldSP6TArray_4X4 vss vdd wl[0] wl[1] wl[2] wl[3] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] bl[0] bl_n[0] bl[1] bl_n[1] OldSP6TArray_4X2
Xinst0x1 vss vdd wl[0] wl[1] wl[2] wl[3] bl[2] bl_n[2] bl[3] bl_n[3] OldSP6TArray_4X2
.ends OldSP6TArray_4X4

.subckt OldSP6TArray_8X4 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] OldSP6TArray_4X4
Xinst1x0 vss vdd wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] OldSP6TArray_4X4
.ends OldSP6TArray_8X4

.subckt OldSP6TArray_8X8 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] OldSP6TArray_8X4
Xinst0x1 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7] OldSP6TArray_8X4
.ends OldSP6TArray_8X8

.subckt OldSP6TBulkConn vdd vss bl bl_n
.ends OldSP6TBulkConn

.subckt OldSP6TBulkConnRow_2 vss vdd bl[0] bl_n[0] bl[1] bl_n[1]
Xinst0 vdd vss bl[0] bl_n[0] OldSP6TBulkConn
Xinst1 vdd vss bl[1] bl_n[1] OldSP6TBulkConn
.ends OldSP6TBulkConnRow_2

.subckt OldSP6TBulkConnRow_4 vss vdd bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3]
Xinst0 vss vdd bl[0] bl_n[0] bl[1] bl_n[1] OldSP6TBulkConnRow_2
Xinst1 vss vdd bl[2] bl_n[2] bl[3] bl_n[3] OldSP6TBulkConnRow_2
.ends OldSP6TBulkConnRow_4

.subckt OldSP6TBulkConnRow_8 vss vdd bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7]
Xinst0 vss vdd bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] OldSP6TBulkConnRow_4
Xinst1 vss vdd bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7] OldSP6TBulkConnRow_4
.ends OldSP6TBulkConnRow_8

.subckt OldSP6TArray_16X8BC vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7] OldSP6TArray_8X8
Xinst1x0 vss vdd wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7] OldSP6TArray_8X8
Xbottombcrow vss vdd bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7] OldSP6TBulkConnRow_8
Xtopbcrow vss vdd bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7] OldSP6TBulkConnRow_8
.ends OldSP6TArray_16X8BC

.subckt OldSP6TTestArray_16X8 vss vdd bl bl_n wl
Xarray vss vdd zero zero zero zero zero zero zero zero wl zero zero zero zero zero zero zero bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] bl bl_n bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7] OldSP6TArray_16X8BC
Xzero vdd vss zero zero_x1
.ends OldSP6TTestArray_16X8

.subckt OldSP6TArray_4X1 vss vdd wl[0] wl[1] wl[2] wl[3] bl[0] bl_n[0]
Xinst0x0 vss vdd wl[0] wl[1] bl[0] bl_n[0] OldSP6TArray_2X1
Xinst1x0 vss vdd wl[2] wl[3] bl[0] bl_n[0] OldSP6TArray_2X1
.ends OldSP6TArray_4X1

.subckt OldSP6TArray_8X1 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] bl[0] bl_n[0] OldSP6TArray_4X1
Xinst1x0 vss vdd wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] OldSP6TArray_4X1
.ends OldSP6TArray_8X1

.subckt OldSP6TArray_16X1BC vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] bl[0] bl_n[0]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] OldSP6TArray_8X1
Xinst1x0 vss vdd wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] bl[0] bl_n[0] OldSP6TArray_8X1
Xbottombcrow vdd vss bl[0] bl_n[0] OldSP6TBulkConn
Xtopbcrow vdd vss bl[0] bl_n[0] OldSP6TBulkConn
.ends OldSP6TArray_16X1BC

.subckt OldSP6TArray_8X2 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] bl[0] bl_n[0] bl[1] bl_n[1] OldSP6TArray_4X2
Xinst1x0 vss vdd wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1] OldSP6TArray_4X2
.ends OldSP6TArray_8X2

.subckt OldSP6TArray_16X2BC vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] bl[0] bl_n[0] bl[1] bl_n[1]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1] OldSP6TArray_8X2
Xinst1x0 vss vdd wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] bl[0] bl_n[0] bl[1] bl_n[1] OldSP6TArray_8X2
Xbottombcrow vss vdd bl[0] bl_n[0] bl[1] bl_n[1] OldSP6TBulkConnRow_2
Xtopbcrow vss vdd bl[0] bl_n[0] bl[1] bl_n[1] OldSP6TBulkConnRow_2
.ends OldSP6TArray_16X2BC

.subckt OldSP6TArray_16X4BC vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] OldSP6TArray_8X4
Xinst1x0 vss vdd wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] OldSP6TArray_8X4
Xbottombcrow vss vdd bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] OldSP6TBulkConnRow_4
Xtopbcrow vss vdd bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] OldSP6TBulkConnRow_4
.ends OldSP6TArray_16X4BC

.subckt OldSP6TArray_6X1 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] bl[0] bl_n[0]
Xinst0x0 vss vdd wl[0] wl[1] wl[2] wl[3] bl[0] bl_n[0] OldSP6TArray_4X1
Xinst1x0 vss vdd wl[4] wl[5] bl[0] bl_n[0] OldSP6TArray_2X1
.ends OldSP6TArray_6X1

.subckt OldSP6TCellConnectOut wl bl bl_n vdd vss bit bit_n
Xpu1 vdd bit_n bit vdd sg13_lv_pmos l=1.3e-07 w=1.5e-07
Xpd1 bit bit_n vss vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpu2 vdd bit bit_n vdd sg13_lv_pmos l=1.3e-07 w=1.5e-07
Xpd2 bit_n bit vss vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg1 bit wl bl vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg2 bit_n wl bl_n vss sg13_lv_nmos l=1.3e-07 w=3e-07
.ends OldSP6TCellConnectOut

.subckt OldSP6TTestArray_16X8C vss vdd bl bl_n bit bit_n wl
Xarray_0 vss vdd zero zero zero zero zero zero zero zero wl zero zero zero zero zero zero zero array_0_bl[0] array_0_bl_n[0] OldSP6TArray_16X1BC
Xarray_1 vss vdd zero zero zero zero zero zero zero zero wl zero zero zero zero zero zero zero array_1_bl[0] array_1_bl_n[0] array_1_bl[1] array_1_bl_n[1] OldSP6TArray_16X2BC
Xarray_2 vss vdd zero zero zero zero zero zero zero zero wl zero zero zero zero zero zero zero array_2_bl[0] array_2_bl_n[0] array_2_bl[1] array_2_bl_n[1] array_2_bl[2] array_2_bl_n[2] array_2_bl[3] array_2_bl_n[3] OldSP6TArray_16X4BC
Xcolbc_0 vdd vss bl bl_n OldSP6TBulkConn
Xcolbc_1 vdd vss bl bl_n OldSP6TBulkConn
Xcolarray_0 vss vdd zero zero zero zero zero zero zero zero bl bl_n OldSP6TArray_8X1
Xcolarray_1 vss vdd zero zero zero zero zero zero bl bl_n OldSP6TArray_6X1
Xbc_noconn zero bl bl_n vdd vss OldSP6TCell
Xbc_conn wl bl bl_n vdd vss bit bit_n OldSP6TCellConnectOut
Xzero vdd vss zero zero_x1
.ends OldSP6TTestArray_16X8C

.subckt SP6TVar21 vss noco_vdd noco_wl noco_bl noco_bl_n co_vdd co_bl co_bl_n co_bit co_bit_n co_wl
Xframe noco_vdd noco_wl NoConn_PAD0x2 co_vdd co_bl_n co_bit co_bit_n NoConn_PAD0x7 NoConn_PAD0x8 NoConn_PAD0x9 vss noco_bl noco_bl_n vss co_bl co_wl NoConn_PAD1x6 NoConn_PAD1x7 NoConn_PAD1x8 NoConn_PAD1x9 PadFrame_SP21
Xtestarray_noco vss noco_vdd noco_bl noco_bl_n noco_wl OldSP6TTestArray_16X8
Xtestarray_co vss co_vdd co_bl co_bl_n co_bit co_bit_n co_wl OldSP6TTestArray_16X8C
.ends SP6TVar21

.subckt PadFrame_DP07 PAD0x0 PAD0x1 PAD0x2 PAD0x3 PAD0x4 PAD0x5 PAD0x6 PAD0x7 PAD0x8 PAD0x9 PAD1x0 PAD1x1 PAD1x2 PAD1x3 PAD1x4 PAD1x5 PAD1x6 PAD1x7 PAD1x8 PAD1x9
XPAD0x0 PAD0x0 BondPad
XPAD0x1 PAD0x1 BondPad
XPAD0x2 PAD0x2 BondPad
XPAD0x3 PAD0x3 BondPad
XPAD0x4 PAD0x4 BondPad
XPAD0x5 PAD0x5 BondPad
XPAD0x6 PAD0x6 BondPad
XPAD0x7 PAD0x7 BondPad
XPAD0x8 PAD0x8 BondPad
XPAD0x9 PAD0x9 BondPad
XPAD1x0 PAD1x0 BondPad
XPAD1x1 PAD1x1 BondPad
XPAD1x2 PAD1x2 BondPad
XPAD1x3 PAD1x3 BondPad
XPAD1x4 PAD1x4 BondPad
XPAD1x5 PAD1x5 BondPad
XPAD1x6 PAD1x6 BondPad
XPAD1x7 PAD1x7 BondPad
XPAD1x8 PAD1x8 BondPad
XPAD1x9 PAD1x9 BondPad
.ends PadFrame_DP07

.subckt DP8TVar7Cell wl1 wl2 bl1 bl1_n bl2 bl2_n vdd vss
Xpu1 vdd bit_n bit vdd sg13_lv_pmos l=1.3e-07 w=3e-07
Xpd1 bit bit_n vss vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpu2 vdd bit bit_n vdd sg13_lv_pmos l=1.3e-07 w=3e-07
Xpd2 bit_n bit vss vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg1 bit wl1 bl1 vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg1n bit_n wl1 bl1_n vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg2 bit wl2 bl2 vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg2n bit_n wl2 bl2_n vss sg13_lv_nmos l=1.3e-07 w=3e-07
.ends DP8TVar7Cell

.subckt DP8TVar7Array_2X1 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0]
Xinst0x0 wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] vdd vss DP8TVar7Cell
Xinst1x0 wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0] vdd vss DP8TVar7Cell
.ends DP8TVar7Array_2X1

.subckt DP8TVar7Array_2X2 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0] DP8TVar7Array_2X1
Xinst0x1 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TVar7Array_2X1
.ends DP8TVar7Array_2X2

.subckt DP8TVar7Array_4X2 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TVar7Array_2X2
Xinst1x0 vss vdd wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TVar7Array_2X2
.ends DP8TVar7Array_4X2

.subckt DP8TVar7Array_4X4 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TVar7Array_4X2
Xinst0x1 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar7Array_4X2
.ends DP8TVar7Array_4X4

.subckt DP8TVar7Array_8X4 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar7Array_4X4
Xinst1x0 vss vdd wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar7Array_4X4
.ends DP8TVar7Array_8X4

.subckt DP8TVar7Array_8X8 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar7Array_8X4
Xinst0x1 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar7Array_8X4
.ends DP8TVar7Array_8X8

.subckt DP8TVar7BulkConn vdd vss bl1 bl2 bl1_n bl2_n
.ends DP8TVar7BulkConn

.subckt DP8TVar7BulkConnRow_2 vss vdd bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1]
Xinst0 vdd vss bl1[0] bl2[0] bl1_n[0] bl2_n[0] DP8TVar7BulkConn
Xinst1 vdd vss bl1[1] bl2[1] bl1_n[1] bl2_n[1] DP8TVar7BulkConn
.ends DP8TVar7BulkConnRow_2

.subckt DP8TVar7BulkConnRow_4 vss vdd bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3]
Xinst0 vss vdd bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TVar7BulkConnRow_2
Xinst1 vss vdd bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar7BulkConnRow_2
.ends DP8TVar7BulkConnRow_4

.subckt DP8TVar7BulkConnRow_8 vss vdd bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0 vss vdd bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar7BulkConnRow_4
Xinst1 vss vdd bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar7BulkConnRow_4
.ends DP8TVar7BulkConnRow_8

.subckt DP8TVar7Array_16X8BC vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] wl1[8] wl2[8] wl1[9] wl2[9] wl1[10] wl2[10] wl1[11] wl2[11] wl1[12] wl2[12] wl1[13] wl2[13] wl1[14] wl2[14] wl1[15] wl2[15] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar7Array_8X8
Xinst1x0 vss vdd wl1[8] wl2[8] wl1[9] wl2[9] wl1[10] wl2[10] wl1[11] wl2[11] wl1[12] wl2[12] wl1[13] wl2[13] wl1[14] wl2[14] wl1[15] wl2[15] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar7Array_8X8
Xbottombcrow vss vdd bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar7BulkConnRow_8
Xtopbcrow vss vdd bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar7BulkConnRow_8
.ends DP8TVar7Array_16X8BC

.subckt DP8TVar7TestArray_16X8 vss vdd wl1 wl2 bl1 bl1_n bl2 bl2_n
Xarray vss vdd zero zero zero zero zero zero zero zero zero zero zero zero zero zero zero zero wl1 wl2 zero zero zero zero zero zero zero zero zero zero zero zero zero zero bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1 bl1_n bl2 bl2_n bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar7Array_16X8BC
Xzero vdd vss zero zero_x1
.ends DP8TVar7TestArray_16X8

.subckt DP8TVar7Array_4X8 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar7Array_4X4
Xinst0x1 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar7Array_4X4
.ends DP8TVar7Array_4X8

.subckt DP8TVar7Array_2X4 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TVar7Array_2X2
Xinst0x1 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar7Array_2X2
.ends DP8TVar7Array_2X4

.subckt DP8TVar7Array_2X8 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar7Array_2X4
Xinst0x1 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar7Array_2X4
.ends DP8TVar7Array_2X8

.subckt DP8TVar7Array_1X2 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1]
Xinst0x0 wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] vdd vss DP8TVar7Cell
Xinst0x1 wl1[0] wl2[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] vdd vss DP8TVar7Cell
.ends DP8TVar7Array_1X2

.subckt DP8TVar7Array_1X4 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3]
Xinst0x0 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TVar7Array_1X2
Xinst0x1 vss vdd wl1[0] wl2[0] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar7Array_1X2
.ends DP8TVar7Array_1X4

.subckt DP8TVar7Array_1X8 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar7Array_1X4
Xinst0x1 vss vdd wl1[0] wl2[0] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar7Array_1X4
.ends DP8TVar7Array_1X8

.subckt DP8TVar7Array_7X8 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar7Array_4X8
Xinst1x0 vss vdd wl1[4] wl2[4] wl1[5] wl2[5] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar7Array_2X8
Xinst2x0 vss vdd wl1[6] wl2[6] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar7Array_1X8
.ends DP8TVar7Array_7X8

.subckt DP8TVar7CellShWL1 wl1 wl2 bl1 bl1_n bl2 bl2_n vdd vss
Xpu1 vdd bit_n bit vdd sg13_lv_pmos l=1.3e-07 w=3e-07
Xpd1 bit bit_n vss vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpu2 vdd bit bit_n vdd sg13_lv_pmos l=1.3e-07 w=3e-07
Xpd2 bit_n bit vss vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg1 bit wl1 bl1 vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg1n bit_n wl1 bl1_n vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg2 bit wl1 bl2 vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg2n bit_n wl1 bl2_n vss sg13_lv_nmos l=1.3e-07 w=3e-07
.ends DP8TVar7CellShWL1

.subckt DP8TVar7ArrayShWL1_1X2 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1]
Xinst0x0 wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] vdd vss DP8TVar7CellShWL1
Xinst0x1 wl1[0] wl2[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] vdd vss DP8TVar7CellShWL1
.ends DP8TVar7ArrayShWL1_1X2

.subckt DP8TVar7ArrayShWL1_1X4 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3]
Xinst0x0 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TVar7ArrayShWL1_1X2
Xinst0x1 vss vdd wl1[0] wl2[0] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar7ArrayShWL1_1X2
.ends DP8TVar7ArrayShWL1_1X4

.subckt DP8TVar7ArrayShWL1_1X8 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar7ArrayShWL1_1X4
Xinst0x1 vss vdd wl1[0] wl2[0] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar7ArrayShWL1_1X4
.ends DP8TVar7ArrayShWL1_1X8

.subckt DP8TVar7CellConnectOut wl1 wl2 bl1 bl1_n bl2 bl2_n vdd vss bit bit_n
Xpu1 vdd bit_n bit vdd sg13_lv_pmos l=1.3e-07 w=3e-07
Xpd1 bit bit_n vss vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpu2 vdd bit bit_n vdd sg13_lv_pmos l=1.3e-07 w=3e-07
Xpd2 bit_n bit vss vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg1 bit wl1 bl1 vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg1n bit_n wl1 bl1_n vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg2 bit wl2 bl2 vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg2n bit_n wl2 bl2_n vss sg13_lv_nmos l=1.3e-07 w=3e-07
.ends DP8TVar7CellConnectOut

.subckt DP8TVar7CellShWL2 wl1 wl2 bl1 bl1_n bl2 bl2_n vdd vss
Xpu1 vdd bit_n bit vdd sg13_lv_pmos l=1.3e-07 w=3e-07
Xpd1 bit bit_n vss vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpu2 vdd bit bit_n vdd sg13_lv_pmos l=1.3e-07 w=3e-07
Xpd2 bit_n bit vss vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg1 bit wl2 bl1 vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg1n bit_n wl2 bl1_n vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg2 bit wl2 bl2 vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg2n bit_n wl2 bl2_n vss sg13_lv_nmos l=1.3e-07 w=3e-07
.ends DP8TVar7CellShWL2

.subckt DP8TVar7ArrayShWL2_1X2 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1]
Xinst0x0 wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] vdd vss DP8TVar7CellShWL2
Xinst0x1 wl1[0] wl2[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] vdd vss DP8TVar7CellShWL2
.ends DP8TVar7ArrayShWL2_1X2

.subckt DP8TVar7ArrayShWL2_1X4 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3]
Xinst0x0 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TVar7ArrayShWL2_1X2
Xinst0x1 vss vdd wl1[0] wl2[0] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar7ArrayShWL2_1X2
.ends DP8TVar7ArrayShWL2_1X4

.subckt DP8TVar7ArrayShWL2_1X8 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar7ArrayShWL2_1X4
Xinst0x1 vss vdd wl1[0] wl2[0] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar7ArrayShWL2_1X4
.ends DP8TVar7ArrayShWL2_1X8

.subckt DP8TVar7Array_6X8 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar7Array_4X8
Xinst1x0 vss vdd wl1[4] wl2[4] wl1[5] wl2[5] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar7Array_2X8
.ends DP8TVar7Array_6X8

.subckt DP8TVar7TestArray_16X8C vss vdd wl1 wl2 bl1 bl1_n bl2 bl2_n bit bit_n
Xbcconn_bot vss vdd bcconn_bot_bl1[0] bcconn_bot_bl1_n[0] bcconn_bot_bl2[0] bcconn_bot_bl2_n[0] bcconn_bot_bl1[1] bcconn_bot_bl1_n[1] bcconn_bot_bl2[1] bcconn_bot_bl2_n[1] bcconn_bot_bl1[2] bcconn_bot_bl1_n[2] bcconn_bot_bl2[2] bcconn_bot_bl2_n[2] bcconn_bot_bl1[3] bcconn_bot_bl1_n[3] bcconn_bot_bl2[3] bcconn_bot_bl2_n[3] bl1 bl1_n bl2 bl2_n bcconn_bot_bl1[5] bcconn_bot_bl1_n[5] bcconn_bot_bl2[5] bcconn_bot_bl2_n[5] bcconn_bot_bl1[6] bcconn_bot_bl1_n[6] bcconn_bot_bl2[6] bcconn_bot_bl2_n[6] bcconn_bot_bl1[7] bcconn_bot_bl1_n[7] bcconn_bot_bl2[7] bcconn_bot_bl2_n[7] DP8TVar7BulkConnRow_8
Xbcconn_top vss vdd bcconn_top_bl1[0] bcconn_top_bl1_n[0] bcconn_top_bl2[0] bcconn_top_bl2_n[0] bcconn_top_bl1[1] bcconn_top_bl1_n[1] bcconn_top_bl2[1] bcconn_top_bl2_n[1] bcconn_top_bl1[2] bcconn_top_bl1_n[2] bcconn_top_bl2[2] bcconn_top_bl2_n[2] bcconn_top_bl1[3] bcconn_top_bl1_n[3] bcconn_top_bl2[3] bcconn_top_bl2_n[3] bl1 bl1_n bl2 bl2_n bcconn_top_bl1[5] bcconn_top_bl1_n[5] bcconn_top_bl2[5] bcconn_top_bl2_n[5] bcconn_top_bl1[6] bcconn_top_bl1_n[6] bcconn_top_bl2[6] bcconn_top_bl2_n[6] bcconn_top_bl1[7] bcconn_top_bl1_n[7] bcconn_top_bl2[7] bcconn_top_bl2_n[7] DP8TVar7BulkConnRow_8
Xarray_bot vss vdd zero zero zero zero zero zero zero zero zero zero zero zero zero zero array_bot_bl1[0] array_bot_bl1_n[0] array_bot_bl2[0] array_bot_bl2_n[0] array_bot_bl1[1] array_bot_bl1_n[1] array_bot_bl2[1] array_bot_bl2_n[1] array_bot_bl1[2] array_bot_bl1_n[2] array_bot_bl2[2] array_bot_bl2_n[2] array_bot_bl1[3] array_bot_bl1_n[3] array_bot_bl2[3] array_bot_bl2_n[3] bl1 bl1_n bl2 bl2_n array_bot_bl1[5] array_bot_bl1_n[5] array_bot_bl2[5] array_bot_bl2_n[5] array_bot_bl1[6] array_bot_bl1_n[6] array_bot_bl2[6] array_bot_bl2_n[6] array_bot_bl1[7] array_bot_bl1_n[7] array_bot_bl2[7] array_bot_bl2_n[7] DP8TVar7Array_7X8
Xshwl1_row vss vdd zero bit shwl1_row_bl1[0] shwl1_row_bl1_n[0] shwl1_row_bl2[0] shwl1_row_bl2_n[0] shwl1_row_bl1[1] shwl1_row_bl1_n[1] shwl1_row_bl2[1] shwl1_row_bl2_n[1] shwl1_row_bl1[2] shwl1_row_bl1_n[2] shwl1_row_bl2[2] shwl1_row_bl2_n[2] shwl1_row_bl1[3] shwl1_row_bl1_n[3] shwl1_row_bl2[3] shwl1_row_bl2_n[3] bl1 bl1_n bl2 bl2_n shwl1_row_bl1[5] shwl1_row_bl1_n[5] shwl1_row_bl2[5] shwl1_row_bl2_n[5] shwl1_row_bl1[6] shwl1_row_bl1_n[6] shwl1_row_bl2[6] shwl1_row_bl2_n[6] shwl1_row_bl1[7] shwl1_row_bl1_n[7] shwl1_row_bl2[7] shwl1_row_bl2_n[7] DP8TVar7ArrayShWL1_1X8
Xcell_cols_left vss vdd wl1 wl2 cell_cols_left_bl1[0] cell_cols_left_bl1_n[0] cell_cols_left_bl2[0] cell_cols_left_bl2_n[0] cell_cols_left_bl1[1] cell_cols_left_bl1_n[1] cell_cols_left_bl2[1] cell_cols_left_bl2_n[1] cell_cols_left_bl1[2] cell_cols_left_bl1_n[2] cell_cols_left_bl2[2] cell_cols_left_bl2_n[2] cell_cols_left_bl1[3] cell_cols_left_bl1_n[3] cell_cols_left_bl2[3] cell_cols_left_bl2_n[3] DP8TVar7Array_1X4
Xconncell wl1 wl2 bl1 bl1_n bl2 bl2_n vdd vss bit bit_n DP8TVar7CellConnectOut
Xfillcell wl1 wl2 fillcell_bl1 fillcell_bl1_n fillcell_bl2 fillcell_bl2_n vdd vss DP8TVar7Cell
Xcell_cols_right vss vdd wl1 wl2 cell_cols_right_bl1[0] cell_cols_right_bl1_n[0] cell_cols_right_bl2[0] cell_cols_right_bl2_n[0] cell_cols_right_bl1[1] cell_cols_right_bl1_n[1] cell_cols_right_bl2[1] cell_cols_right_bl2_n[1] DP8TVar7Array_1X2
Xshwl2_row vss vdd bit_n zero shwl2_row_bl1[0] shwl2_row_bl1_n[0] shwl2_row_bl2[0] shwl2_row_bl2_n[0] shwl2_row_bl1[1] shwl2_row_bl1_n[1] shwl2_row_bl2[1] shwl2_row_bl2_n[1] shwl2_row_bl1[2] shwl2_row_bl1_n[2] shwl2_row_bl2[2] shwl2_row_bl2_n[2] shwl2_row_bl1[3] shwl2_row_bl1_n[3] shwl2_row_bl2[3] shwl2_row_bl2_n[3] bl1 bl1_n bl2 bl2_n shwl2_row_bl1[5] shwl2_row_bl1_n[5] shwl2_row_bl2[5] shwl2_row_bl2_n[5] shwl2_row_bl1[6] shwl2_row_bl1_n[6] shwl2_row_bl2[6] shwl2_row_bl2_n[6] shwl2_row_bl1[7] shwl2_row_bl1_n[7] shwl2_row_bl2[7] shwl2_row_bl2_n[7] DP8TVar7ArrayShWL2_1X8
Xarray_top vss vdd zero zero zero zero zero zero zero zero zero zero zero zero array_top_bl1[0] array_top_bl1_n[0] array_top_bl2[0] array_top_bl2_n[0] array_top_bl1[1] array_top_bl1_n[1] array_top_bl2[1] array_top_bl2_n[1] array_top_bl1[2] array_top_bl1_n[2] array_top_bl2[2] array_top_bl2_n[2] array_top_bl1[3] array_top_bl1_n[3] array_top_bl2[3] array_top_bl2_n[3] bl1 bl1_n bl2 bl2_n array_top_bl1[5] array_top_bl1_n[5] array_top_bl2[5] array_top_bl2_n[5] array_top_bl1[6] array_top_bl1_n[6] array_top_bl2[6] array_top_bl2_n[6] array_top_bl1[7] array_top_bl1_n[7] array_top_bl2[7] array_top_bl2_n[7] DP8TVar7Array_6X8
Xzero vdd vss zero zero_x1
.ends DP8TVar7TestArray_16X8C

.subckt DP8TVar7 vss noco_vdd noco_wl1 noco_wl2 noco_bl1 noco_bl1_n noco_bl2 noco_bl2_n co_vdd co_bit co_bit_n co_wl1 co_wl2 co_bl1 co_bl1_n co_bl2_n co_bl2
Xframe noco_vdd noco_wl1 noco_wl2 noco_bl2 co_vdd co_bit co_bit_n co_wl1 co_wl2 NoConn_PAD0x9 vss noco_bl1 noco_bl1_n noco_bl2_n vss co_bl1 co_bl1_n co_bl2_n co_bl2 NoConn_PAD1x9 PadFrame_DP07
Xtestarray_noco vss noco_vdd noco_wl1 noco_wl2 noco_bl1 noco_bl1_n noco_bl2 noco_bl2_n DP8TVar7TestArray_16X8
Xtestarray_co vss co_vdd co_wl1 co_wl2 co_bl1 co_bl1_n co_bl2 co_bl2_n co_bit co_bit_n DP8TVar7TestArray_16X8C
.ends DP8TVar7

.subckt PadFrame_DP08 PAD0x0 PAD0x1 PAD0x2 PAD0x3 PAD0x4 PAD0x5 PAD0x6 PAD0x7 PAD0x8 PAD0x9 PAD1x0 PAD1x1 PAD1x2 PAD1x3 PAD1x4 PAD1x5 PAD1x6 PAD1x7 PAD1x8 PAD1x9
XPAD0x0 PAD0x0 BondPad
XPAD0x1 PAD0x1 BondPad
XPAD0x2 PAD0x2 BondPad
XPAD0x3 PAD0x3 BondPad
XPAD0x4 PAD0x4 BondPad
XPAD0x5 PAD0x5 BondPad
XPAD0x6 PAD0x6 BondPad
XPAD0x7 PAD0x7 BondPad
XPAD0x8 PAD0x8 BondPad
XPAD0x9 PAD0x9 BondPad
XPAD1x0 PAD1x0 BondPad
XPAD1x1 PAD1x1 BondPad
XPAD1x2 PAD1x2 BondPad
XPAD1x3 PAD1x3 BondPad
XPAD1x4 PAD1x4 BondPad
XPAD1x5 PAD1x5 BondPad
XPAD1x6 PAD1x6 BondPad
XPAD1x7 PAD1x7 BondPad
XPAD1x8 PAD1x8 BondPad
XPAD1x9 PAD1x9 BondPad
.ends PadFrame_DP08

.subckt DP8TVar8Cell wl1 wl2 bl1 bl1_n bl2 bl2_n vdd vss
Xpu1 vdd bit_n bit vdd sg13_lv_pmos l=1.3e-07 w=2e-07
Xpd1 bit bit_n vss vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpu2 vdd bit bit_n vdd sg13_lv_pmos l=1.3e-07 w=2e-07
Xpd2 bit_n bit vss vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg1 bit wl1 bl1 vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg1n bit_n wl1 bl1_n vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg2 bit wl2 bl2 vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg2n bit_n wl2 bl2_n vss sg13_lv_nmos l=1.3e-07 w=3e-07
.ends DP8TVar8Cell

.subckt DP8TVar8Array_2X1 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0]
Xinst0x0 wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] vdd vss DP8TVar8Cell
Xinst1x0 wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0] vdd vss DP8TVar8Cell
.ends DP8TVar8Array_2X1

.subckt DP8TVar8Array_2X2 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0] DP8TVar8Array_2X1
Xinst0x1 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TVar8Array_2X1
.ends DP8TVar8Array_2X2

.subckt DP8TVar8Array_4X2 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TVar8Array_2X2
Xinst1x0 vss vdd wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TVar8Array_2X2
.ends DP8TVar8Array_4X2

.subckt DP8TVar8Array_4X4 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TVar8Array_4X2
Xinst0x1 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar8Array_4X2
.ends DP8TVar8Array_4X4

.subckt DP8TVar8Array_8X4 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar8Array_4X4
Xinst1x0 vss vdd wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar8Array_4X4
.ends DP8TVar8Array_8X4

.subckt DP8TVar8Array_8X8 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar8Array_8X4
Xinst0x1 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar8Array_8X4
.ends DP8TVar8Array_8X8

.subckt DP8TVar8BulkConn vdd vss bl1 bl2 bl1_n bl2_n
.ends DP8TVar8BulkConn

.subckt DP8TVar8BulkConnRow_2 vss vdd bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1]
Xinst0 vdd vss bl1[0] bl2[0] bl1_n[0] bl2_n[0] DP8TVar8BulkConn
Xinst1 vdd vss bl1[1] bl2[1] bl1_n[1] bl2_n[1] DP8TVar8BulkConn
.ends DP8TVar8BulkConnRow_2

.subckt DP8TVar8BulkConnRow_4 vss vdd bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3]
Xinst0 vss vdd bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TVar8BulkConnRow_2
Xinst1 vss vdd bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar8BulkConnRow_2
.ends DP8TVar8BulkConnRow_4

.subckt DP8TVar8BulkConnRow_8 vss vdd bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0 vss vdd bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar8BulkConnRow_4
Xinst1 vss vdd bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar8BulkConnRow_4
.ends DP8TVar8BulkConnRow_8

.subckt DP8TVar8Array_16X8BC vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] wl1[8] wl2[8] wl1[9] wl2[9] wl1[10] wl2[10] wl1[11] wl2[11] wl1[12] wl2[12] wl1[13] wl2[13] wl1[14] wl2[14] wl1[15] wl2[15] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar8Array_8X8
Xinst1x0 vss vdd wl1[8] wl2[8] wl1[9] wl2[9] wl1[10] wl2[10] wl1[11] wl2[11] wl1[12] wl2[12] wl1[13] wl2[13] wl1[14] wl2[14] wl1[15] wl2[15] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar8Array_8X8
Xbottombcrow vss vdd bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar8BulkConnRow_8
Xtopbcrow vss vdd bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar8BulkConnRow_8
.ends DP8TVar8Array_16X8BC

.subckt DP8TVar8TestArray_16X8 vss vdd wl1 wl2 bl1 bl1_n bl2 bl2_n
Xarray vss vdd zero zero zero zero zero zero zero zero zero zero zero zero zero zero zero zero wl1 wl2 zero zero zero zero zero zero zero zero zero zero zero zero zero zero bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1 bl1_n bl2 bl2_n bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar8Array_16X8BC
Xzero vdd vss zero zero_x1
.ends DP8TVar8TestArray_16X8

.subckt DP8TVar8Array_4X8 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar8Array_4X4
Xinst0x1 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar8Array_4X4
.ends DP8TVar8Array_4X8

.subckt DP8TVar8Array_2X4 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TVar8Array_2X2
Xinst0x1 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar8Array_2X2
.ends DP8TVar8Array_2X4

.subckt DP8TVar8Array_2X8 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar8Array_2X4
Xinst0x1 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar8Array_2X4
.ends DP8TVar8Array_2X8

.subckt DP8TVar8Array_1X2 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1]
Xinst0x0 wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] vdd vss DP8TVar8Cell
Xinst0x1 wl1[0] wl2[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] vdd vss DP8TVar8Cell
.ends DP8TVar8Array_1X2

.subckt DP8TVar8Array_1X4 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3]
Xinst0x0 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TVar8Array_1X2
Xinst0x1 vss vdd wl1[0] wl2[0] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar8Array_1X2
.ends DP8TVar8Array_1X4

.subckt DP8TVar8Array_1X8 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar8Array_1X4
Xinst0x1 vss vdd wl1[0] wl2[0] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar8Array_1X4
.ends DP8TVar8Array_1X8

.subckt DP8TVar8Array_7X8 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar8Array_4X8
Xinst1x0 vss vdd wl1[4] wl2[4] wl1[5] wl2[5] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar8Array_2X8
Xinst2x0 vss vdd wl1[6] wl2[6] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar8Array_1X8
.ends DP8TVar8Array_7X8

.subckt DP8TVar8CellShWL1 wl1 wl2 bl1 bl1_n bl2 bl2_n vdd vss
Xpu1 vdd bit_n bit vdd sg13_lv_pmos l=1.3e-07 w=2e-07
Xpd1 bit bit_n vss vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpu2 vdd bit bit_n vdd sg13_lv_pmos l=1.3e-07 w=2e-07
Xpd2 bit_n bit vss vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg1 bit wl1 bl1 vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg1n bit_n wl1 bl1_n vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg2 bit wl1 bl2 vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg2n bit_n wl1 bl2_n vss sg13_lv_nmos l=1.3e-07 w=3e-07
.ends DP8TVar8CellShWL1

.subckt DP8TVar8ArrayShWL1_1X2 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1]
Xinst0x0 wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] vdd vss DP8TVar8CellShWL1
Xinst0x1 wl1[0] wl2[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] vdd vss DP8TVar8CellShWL1
.ends DP8TVar8ArrayShWL1_1X2

.subckt DP8TVar8ArrayShWL1_1X4 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3]
Xinst0x0 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TVar8ArrayShWL1_1X2
Xinst0x1 vss vdd wl1[0] wl2[0] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar8ArrayShWL1_1X2
.ends DP8TVar8ArrayShWL1_1X4

.subckt DP8TVar8ArrayShWL1_1X8 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar8ArrayShWL1_1X4
Xinst0x1 vss vdd wl1[0] wl2[0] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar8ArrayShWL1_1X4
.ends DP8TVar8ArrayShWL1_1X8

.subckt DP8TVar8CellConnectOut wl1 wl2 bl1 bl1_n bl2 bl2_n vdd vss bit bit_n
Xpu1 vdd bit_n bit vdd sg13_lv_pmos l=1.3e-07 w=2e-07
Xpd1 bit bit_n vss vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpu2 vdd bit bit_n vdd sg13_lv_pmos l=1.3e-07 w=2e-07
Xpd2 bit_n bit vss vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg1 bit wl1 bl1 vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg1n bit_n wl1 bl1_n vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg2 bit wl2 bl2 vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg2n bit_n wl2 bl2_n vss sg13_lv_nmos l=1.3e-07 w=3e-07
.ends DP8TVar8CellConnectOut

.subckt DP8TVar8CellShWL2 wl1 wl2 bl1 bl1_n bl2 bl2_n vdd vss
Xpu1 vdd bit_n bit vdd sg13_lv_pmos l=1.3e-07 w=2e-07
Xpd1 bit bit_n vss vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpu2 vdd bit bit_n vdd sg13_lv_pmos l=1.3e-07 w=2e-07
Xpd2 bit_n bit vss vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg1 bit wl2 bl1 vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg1n bit_n wl2 bl1_n vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg2 bit wl2 bl2 vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg2n bit_n wl2 bl2_n vss sg13_lv_nmos l=1.3e-07 w=3e-07
.ends DP8TVar8CellShWL2

.subckt DP8TVar8ArrayShWL2_1X2 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1]
Xinst0x0 wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] vdd vss DP8TVar8CellShWL2
Xinst0x1 wl1[0] wl2[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] vdd vss DP8TVar8CellShWL2
.ends DP8TVar8ArrayShWL2_1X2

.subckt DP8TVar8ArrayShWL2_1X4 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3]
Xinst0x0 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TVar8ArrayShWL2_1X2
Xinst0x1 vss vdd wl1[0] wl2[0] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar8ArrayShWL2_1X2
.ends DP8TVar8ArrayShWL2_1X4

.subckt DP8TVar8ArrayShWL2_1X8 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar8ArrayShWL2_1X4
Xinst0x1 vss vdd wl1[0] wl2[0] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar8ArrayShWL2_1X4
.ends DP8TVar8ArrayShWL2_1X8

.subckt DP8TVar8Array_6X8 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar8Array_4X8
Xinst1x0 vss vdd wl1[4] wl2[4] wl1[5] wl2[5] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar8Array_2X8
.ends DP8TVar8Array_6X8

.subckt DP8TVar8TestArray_16X8C vss vdd wl1 wl2 bl1 bl1_n bl2 bl2_n bit bit_n
Xbcconn_bot vss vdd bcconn_bot_bl1[0] bcconn_bot_bl1_n[0] bcconn_bot_bl2[0] bcconn_bot_bl2_n[0] bcconn_bot_bl1[1] bcconn_bot_bl1_n[1] bcconn_bot_bl2[1] bcconn_bot_bl2_n[1] bcconn_bot_bl1[2] bcconn_bot_bl1_n[2] bcconn_bot_bl2[2] bcconn_bot_bl2_n[2] bcconn_bot_bl1[3] bcconn_bot_bl1_n[3] bcconn_bot_bl2[3] bcconn_bot_bl2_n[3] bl1 bl1_n bl2 bl2_n bcconn_bot_bl1[5] bcconn_bot_bl1_n[5] bcconn_bot_bl2[5] bcconn_bot_bl2_n[5] bcconn_bot_bl1[6] bcconn_bot_bl1_n[6] bcconn_bot_bl2[6] bcconn_bot_bl2_n[6] bcconn_bot_bl1[7] bcconn_bot_bl1_n[7] bcconn_bot_bl2[7] bcconn_bot_bl2_n[7] DP8TVar8BulkConnRow_8
Xbcconn_top vss vdd bcconn_top_bl1[0] bcconn_top_bl1_n[0] bcconn_top_bl2[0] bcconn_top_bl2_n[0] bcconn_top_bl1[1] bcconn_top_bl1_n[1] bcconn_top_bl2[1] bcconn_top_bl2_n[1] bcconn_top_bl1[2] bcconn_top_bl1_n[2] bcconn_top_bl2[2] bcconn_top_bl2_n[2] bcconn_top_bl1[3] bcconn_top_bl1_n[3] bcconn_top_bl2[3] bcconn_top_bl2_n[3] bl1 bl1_n bl2 bl2_n bcconn_top_bl1[5] bcconn_top_bl1_n[5] bcconn_top_bl2[5] bcconn_top_bl2_n[5] bcconn_top_bl1[6] bcconn_top_bl1_n[6] bcconn_top_bl2[6] bcconn_top_bl2_n[6] bcconn_top_bl1[7] bcconn_top_bl1_n[7] bcconn_top_bl2[7] bcconn_top_bl2_n[7] DP8TVar8BulkConnRow_8
Xarray_bot vss vdd zero zero zero zero zero zero zero zero zero zero zero zero zero zero array_bot_bl1[0] array_bot_bl1_n[0] array_bot_bl2[0] array_bot_bl2_n[0] array_bot_bl1[1] array_bot_bl1_n[1] array_bot_bl2[1] array_bot_bl2_n[1] array_bot_bl1[2] array_bot_bl1_n[2] array_bot_bl2[2] array_bot_bl2_n[2] array_bot_bl1[3] array_bot_bl1_n[3] array_bot_bl2[3] array_bot_bl2_n[3] bl1 bl1_n bl2 bl2_n array_bot_bl1[5] array_bot_bl1_n[5] array_bot_bl2[5] array_bot_bl2_n[5] array_bot_bl1[6] array_bot_bl1_n[6] array_bot_bl2[6] array_bot_bl2_n[6] array_bot_bl1[7] array_bot_bl1_n[7] array_bot_bl2[7] array_bot_bl2_n[7] DP8TVar8Array_7X8
Xshwl1_row vss vdd zero bit shwl1_row_bl1[0] shwl1_row_bl1_n[0] shwl1_row_bl2[0] shwl1_row_bl2_n[0] shwl1_row_bl1[1] shwl1_row_bl1_n[1] shwl1_row_bl2[1] shwl1_row_bl2_n[1] shwl1_row_bl1[2] shwl1_row_bl1_n[2] shwl1_row_bl2[2] shwl1_row_bl2_n[2] shwl1_row_bl1[3] shwl1_row_bl1_n[3] shwl1_row_bl2[3] shwl1_row_bl2_n[3] bl1 bl1_n bl2 bl2_n shwl1_row_bl1[5] shwl1_row_bl1_n[5] shwl1_row_bl2[5] shwl1_row_bl2_n[5] shwl1_row_bl1[6] shwl1_row_bl1_n[6] shwl1_row_bl2[6] shwl1_row_bl2_n[6] shwl1_row_bl1[7] shwl1_row_bl1_n[7] shwl1_row_bl2[7] shwl1_row_bl2_n[7] DP8TVar8ArrayShWL1_1X8
Xcell_cols_left vss vdd wl1 wl2 cell_cols_left_bl1[0] cell_cols_left_bl1_n[0] cell_cols_left_bl2[0] cell_cols_left_bl2_n[0] cell_cols_left_bl1[1] cell_cols_left_bl1_n[1] cell_cols_left_bl2[1] cell_cols_left_bl2_n[1] cell_cols_left_bl1[2] cell_cols_left_bl1_n[2] cell_cols_left_bl2[2] cell_cols_left_bl2_n[2] cell_cols_left_bl1[3] cell_cols_left_bl1_n[3] cell_cols_left_bl2[3] cell_cols_left_bl2_n[3] DP8TVar8Array_1X4
Xconncell wl1 wl2 bl1 bl1_n bl2 bl2_n vdd vss bit bit_n DP8TVar8CellConnectOut
Xfillcell wl1 wl2 fillcell_bl1 fillcell_bl1_n fillcell_bl2 fillcell_bl2_n vdd vss DP8TVar8Cell
Xcell_cols_right vss vdd wl1 wl2 cell_cols_right_bl1[0] cell_cols_right_bl1_n[0] cell_cols_right_bl2[0] cell_cols_right_bl2_n[0] cell_cols_right_bl1[1] cell_cols_right_bl1_n[1] cell_cols_right_bl2[1] cell_cols_right_bl2_n[1] DP8TVar8Array_1X2
Xshwl2_row vss vdd bit_n zero shwl2_row_bl1[0] shwl2_row_bl1_n[0] shwl2_row_bl2[0] shwl2_row_bl2_n[0] shwl2_row_bl1[1] shwl2_row_bl1_n[1] shwl2_row_bl2[1] shwl2_row_bl2_n[1] shwl2_row_bl1[2] shwl2_row_bl1_n[2] shwl2_row_bl2[2] shwl2_row_bl2_n[2] shwl2_row_bl1[3] shwl2_row_bl1_n[3] shwl2_row_bl2[3] shwl2_row_bl2_n[3] bl1 bl1_n bl2 bl2_n shwl2_row_bl1[5] shwl2_row_bl1_n[5] shwl2_row_bl2[5] shwl2_row_bl2_n[5] shwl2_row_bl1[6] shwl2_row_bl1_n[6] shwl2_row_bl2[6] shwl2_row_bl2_n[6] shwl2_row_bl1[7] shwl2_row_bl1_n[7] shwl2_row_bl2[7] shwl2_row_bl2_n[7] DP8TVar8ArrayShWL2_1X8
Xarray_top vss vdd zero zero zero zero zero zero zero zero zero zero zero zero array_top_bl1[0] array_top_bl1_n[0] array_top_bl2[0] array_top_bl2_n[0] array_top_bl1[1] array_top_bl1_n[1] array_top_bl2[1] array_top_bl2_n[1] array_top_bl1[2] array_top_bl1_n[2] array_top_bl2[2] array_top_bl2_n[2] array_top_bl1[3] array_top_bl1_n[3] array_top_bl2[3] array_top_bl2_n[3] bl1 bl1_n bl2 bl2_n array_top_bl1[5] array_top_bl1_n[5] array_top_bl2[5] array_top_bl2_n[5] array_top_bl1[6] array_top_bl1_n[6] array_top_bl2[6] array_top_bl2_n[6] array_top_bl1[7] array_top_bl1_n[7] array_top_bl2[7] array_top_bl2_n[7] DP8TVar8Array_6X8
Xzero vdd vss zero zero_x1
.ends DP8TVar8TestArray_16X8C

.subckt DP8TVar8 vss noco_vdd noco_wl1 noco_wl2 noco_bl1 noco_bl1_n noco_bl2 noco_bl2_n co_vdd co_bit co_bit_n co_wl1 co_wl2 co_bl1 co_bl1_n co_bl2_n co_bl2
Xframe noco_vdd noco_wl1 noco_wl2 noco_bl2 co_vdd co_bit co_bit_n co_wl1 co_wl2 NoConn_PAD0x9 vss noco_bl1 noco_bl1_n noco_bl2_n vss co_bl1 co_bl1_n co_bl2_n co_bl2 NoConn_PAD1x9 PadFrame_DP08
Xtestarray_noco vss noco_vdd noco_wl1 noco_wl2 noco_bl1 noco_bl1_n noco_bl2 noco_bl2_n DP8TVar8TestArray_16X8
Xtestarray_co vss co_vdd co_wl1 co_wl2 co_bl1 co_bl1_n co_bl2 co_bl2_n co_bit co_bit_n DP8TVar8TestArray_16X8C
.ends DP8TVar8

.subckt PadFrame_DP09 PAD0x0 PAD0x1 PAD0x2 PAD0x3 PAD0x4 PAD0x5 PAD0x6 PAD0x7 PAD0x8 PAD0x9 PAD1x0 PAD1x1 PAD1x2 PAD1x3 PAD1x4 PAD1x5 PAD1x6 PAD1x7 PAD1x8 PAD1x9
XPAD0x0 PAD0x0 BondPad
XPAD0x1 PAD0x1 BondPad
XPAD0x2 PAD0x2 BondPad
XPAD0x3 PAD0x3 BondPad
XPAD0x4 PAD0x4 BondPad
XPAD0x5 PAD0x5 BondPad
XPAD0x6 PAD0x6 BondPad
XPAD0x7 PAD0x7 BondPad
XPAD0x8 PAD0x8 BondPad
XPAD0x9 PAD0x9 BondPad
XPAD1x0 PAD1x0 BondPad
XPAD1x1 PAD1x1 BondPad
XPAD1x2 PAD1x2 BondPad
XPAD1x3 PAD1x3 BondPad
XPAD1x4 PAD1x4 BondPad
XPAD1x5 PAD1x5 BondPad
XPAD1x6 PAD1x6 BondPad
XPAD1x7 PAD1x7 BondPad
XPAD1x8 PAD1x8 BondPad
XPAD1x9 PAD1x9 BondPad
.ends PadFrame_DP09

.subckt DP8TVar9Cell wl1 wl2 bl1 bl1_n bl2 bl2_n vdd vss
Xpu1 vdd bit_n bit vdd sg13_lv_pmos l=1.3e-07 w=1.5e-07
Xpd1 bit bit_n vss vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpu2 vdd bit bit_n vdd sg13_lv_pmos l=1.3e-07 w=1.5e-07
Xpd2 bit_n bit vss vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg1 bit wl1 bl1 vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg1n bit_n wl1 bl1_n vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg2 bit wl2 bl2 vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg2n bit_n wl2 bl2_n vss sg13_lv_nmos l=1.3e-07 w=3e-07
.ends DP8TVar9Cell

.subckt DP8TVar9Array_2X1 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0]
Xinst0x0 wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] vdd vss DP8TVar9Cell
Xinst1x0 wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0] vdd vss DP8TVar9Cell
.ends DP8TVar9Array_2X1

.subckt DP8TVar9Array_2X2 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0] DP8TVar9Array_2X1
Xinst0x1 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TVar9Array_2X1
.ends DP8TVar9Array_2X2

.subckt DP8TVar9Array_4X2 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TVar9Array_2X2
Xinst1x0 vss vdd wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TVar9Array_2X2
.ends DP8TVar9Array_4X2

.subckt DP8TVar9Array_4X4 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TVar9Array_4X2
Xinst0x1 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar9Array_4X2
.ends DP8TVar9Array_4X4

.subckt DP8TVar9Array_8X4 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar9Array_4X4
Xinst1x0 vss vdd wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar9Array_4X4
.ends DP8TVar9Array_8X4

.subckt DP8TVar9Array_8X8 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar9Array_8X4
Xinst0x1 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar9Array_8X4
.ends DP8TVar9Array_8X8

.subckt DP8TVar9BulkConn vdd vss bl1 bl2 bl1_n bl2_n
.ends DP8TVar9BulkConn

.subckt DP8TVar9BulkConnRow_2 vss vdd bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1]
Xinst0 vdd vss bl1[0] bl2[0] bl1_n[0] bl2_n[0] DP8TVar9BulkConn
Xinst1 vdd vss bl1[1] bl2[1] bl1_n[1] bl2_n[1] DP8TVar9BulkConn
.ends DP8TVar9BulkConnRow_2

.subckt DP8TVar9BulkConnRow_4 vss vdd bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3]
Xinst0 vss vdd bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TVar9BulkConnRow_2
Xinst1 vss vdd bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar9BulkConnRow_2
.ends DP8TVar9BulkConnRow_4

.subckt DP8TVar9BulkConnRow_8 vss vdd bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0 vss vdd bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar9BulkConnRow_4
Xinst1 vss vdd bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar9BulkConnRow_4
.ends DP8TVar9BulkConnRow_8

.subckt DP8TVar9Array_16X8BC vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] wl1[8] wl2[8] wl1[9] wl2[9] wl1[10] wl2[10] wl1[11] wl2[11] wl1[12] wl2[12] wl1[13] wl2[13] wl1[14] wl2[14] wl1[15] wl2[15] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar9Array_8X8
Xinst1x0 vss vdd wl1[8] wl2[8] wl1[9] wl2[9] wl1[10] wl2[10] wl1[11] wl2[11] wl1[12] wl2[12] wl1[13] wl2[13] wl1[14] wl2[14] wl1[15] wl2[15] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar9Array_8X8
Xbottombcrow vss vdd bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar9BulkConnRow_8
Xtopbcrow vss vdd bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar9BulkConnRow_8
.ends DP8TVar9Array_16X8BC

.subckt DP8TVar9TestArray_16X8 vss vdd wl1 wl2 bl1 bl1_n bl2 bl2_n
Xarray vss vdd zero zero zero zero zero zero zero zero zero zero zero zero zero zero zero zero wl1 wl2 zero zero zero zero zero zero zero zero zero zero zero zero zero zero bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1 bl1_n bl2 bl2_n bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar9Array_16X8BC
Xzero vdd vss zero zero_x1
.ends DP8TVar9TestArray_16X8

.subckt DP8TVar9Array_4X8 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar9Array_4X4
Xinst0x1 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar9Array_4X4
.ends DP8TVar9Array_4X8

.subckt DP8TVar9Array_2X4 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TVar9Array_2X2
Xinst0x1 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar9Array_2X2
.ends DP8TVar9Array_2X4

.subckt DP8TVar9Array_2X8 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar9Array_2X4
Xinst0x1 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar9Array_2X4
.ends DP8TVar9Array_2X8

.subckt DP8TVar9Array_1X2 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1]
Xinst0x0 wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] vdd vss DP8TVar9Cell
Xinst0x1 wl1[0] wl2[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] vdd vss DP8TVar9Cell
.ends DP8TVar9Array_1X2

.subckt DP8TVar9Array_1X4 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3]
Xinst0x0 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TVar9Array_1X2
Xinst0x1 vss vdd wl1[0] wl2[0] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar9Array_1X2
.ends DP8TVar9Array_1X4

.subckt DP8TVar9Array_1X8 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar9Array_1X4
Xinst0x1 vss vdd wl1[0] wl2[0] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar9Array_1X4
.ends DP8TVar9Array_1X8

.subckt DP8TVar9Array_7X8 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar9Array_4X8
Xinst1x0 vss vdd wl1[4] wl2[4] wl1[5] wl2[5] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar9Array_2X8
Xinst2x0 vss vdd wl1[6] wl2[6] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar9Array_1X8
.ends DP8TVar9Array_7X8

.subckt DP8TVar9CellShWL1 wl1 wl2 bl1 bl1_n bl2 bl2_n vdd vss
Xpu1 vdd bit_n bit vdd sg13_lv_pmos l=1.3e-07 w=1.5e-07
Xpd1 bit bit_n vss vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpu2 vdd bit bit_n vdd sg13_lv_pmos l=1.3e-07 w=1.5e-07
Xpd2 bit_n bit vss vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg1 bit wl1 bl1 vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg1n bit_n wl1 bl1_n vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg2 bit wl1 bl2 vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg2n bit_n wl1 bl2_n vss sg13_lv_nmos l=1.3e-07 w=3e-07
.ends DP8TVar9CellShWL1

.subckt DP8TVar9ArrayShWL1_1X2 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1]
Xinst0x0 wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] vdd vss DP8TVar9CellShWL1
Xinst0x1 wl1[0] wl2[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] vdd vss DP8TVar9CellShWL1
.ends DP8TVar9ArrayShWL1_1X2

.subckt DP8TVar9ArrayShWL1_1X4 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3]
Xinst0x0 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TVar9ArrayShWL1_1X2
Xinst0x1 vss vdd wl1[0] wl2[0] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar9ArrayShWL1_1X2
.ends DP8TVar9ArrayShWL1_1X4

.subckt DP8TVar9ArrayShWL1_1X8 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar9ArrayShWL1_1X4
Xinst0x1 vss vdd wl1[0] wl2[0] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar9ArrayShWL1_1X4
.ends DP8TVar9ArrayShWL1_1X8

.subckt DP8TVar9CellConnectOut wl1 wl2 bl1 bl1_n bl2 bl2_n vdd vss bit bit_n
Xpu1 vdd bit_n bit vdd sg13_lv_pmos l=1.3e-07 w=1.5e-07
Xpd1 bit bit_n vss vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpu2 vdd bit bit_n vdd sg13_lv_pmos l=1.3e-07 w=1.5e-07
Xpd2 bit_n bit vss vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg1 bit wl1 bl1 vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg1n bit_n wl1 bl1_n vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg2 bit wl2 bl2 vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg2n bit_n wl2 bl2_n vss sg13_lv_nmos l=1.3e-07 w=3e-07
.ends DP8TVar9CellConnectOut

.subckt DP8TVar9CellShWL2 wl1 wl2 bl1 bl1_n bl2 bl2_n vdd vss
Xpu1 vdd bit_n bit vdd sg13_lv_pmos l=1.3e-07 w=1.5e-07
Xpd1 bit bit_n vss vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpu2 vdd bit bit_n vdd sg13_lv_pmos l=1.3e-07 w=1.5e-07
Xpd2 bit_n bit vss vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg1 bit wl2 bl1 vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg1n bit_n wl2 bl1_n vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg2 bit wl2 bl2 vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg2n bit_n wl2 bl2_n vss sg13_lv_nmos l=1.3e-07 w=3e-07
.ends DP8TVar9CellShWL2

.subckt DP8TVar9ArrayShWL2_1X2 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1]
Xinst0x0 wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] vdd vss DP8TVar9CellShWL2
Xinst0x1 wl1[0] wl2[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] vdd vss DP8TVar9CellShWL2
.ends DP8TVar9ArrayShWL2_1X2

.subckt DP8TVar9ArrayShWL2_1X4 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3]
Xinst0x0 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TVar9ArrayShWL2_1X2
Xinst0x1 vss vdd wl1[0] wl2[0] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar9ArrayShWL2_1X2
.ends DP8TVar9ArrayShWL2_1X4

.subckt DP8TVar9ArrayShWL2_1X8 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar9ArrayShWL2_1X4
Xinst0x1 vss vdd wl1[0] wl2[0] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar9ArrayShWL2_1X4
.ends DP8TVar9ArrayShWL2_1X8

.subckt DP8TVar9Array_6X8 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar9Array_4X8
Xinst1x0 vss vdd wl1[4] wl2[4] wl1[5] wl2[5] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar9Array_2X8
.ends DP8TVar9Array_6X8

.subckt DP8TVar9TestArray_16X8C vss vdd wl1 wl2 bl1 bl1_n bl2 bl2_n bit bit_n
Xbcconn_bot vss vdd bcconn_bot_bl1[0] bcconn_bot_bl1_n[0] bcconn_bot_bl2[0] bcconn_bot_bl2_n[0] bcconn_bot_bl1[1] bcconn_bot_bl1_n[1] bcconn_bot_bl2[1] bcconn_bot_bl2_n[1] bcconn_bot_bl1[2] bcconn_bot_bl1_n[2] bcconn_bot_bl2[2] bcconn_bot_bl2_n[2] bcconn_bot_bl1[3] bcconn_bot_bl1_n[3] bcconn_bot_bl2[3] bcconn_bot_bl2_n[3] bl1 bl1_n bl2 bl2_n bcconn_bot_bl1[5] bcconn_bot_bl1_n[5] bcconn_bot_bl2[5] bcconn_bot_bl2_n[5] bcconn_bot_bl1[6] bcconn_bot_bl1_n[6] bcconn_bot_bl2[6] bcconn_bot_bl2_n[6] bcconn_bot_bl1[7] bcconn_bot_bl1_n[7] bcconn_bot_bl2[7] bcconn_bot_bl2_n[7] DP8TVar9BulkConnRow_8
Xbcconn_top vss vdd bcconn_top_bl1[0] bcconn_top_bl1_n[0] bcconn_top_bl2[0] bcconn_top_bl2_n[0] bcconn_top_bl1[1] bcconn_top_bl1_n[1] bcconn_top_bl2[1] bcconn_top_bl2_n[1] bcconn_top_bl1[2] bcconn_top_bl1_n[2] bcconn_top_bl2[2] bcconn_top_bl2_n[2] bcconn_top_bl1[3] bcconn_top_bl1_n[3] bcconn_top_bl2[3] bcconn_top_bl2_n[3] bl1 bl1_n bl2 bl2_n bcconn_top_bl1[5] bcconn_top_bl1_n[5] bcconn_top_bl2[5] bcconn_top_bl2_n[5] bcconn_top_bl1[6] bcconn_top_bl1_n[6] bcconn_top_bl2[6] bcconn_top_bl2_n[6] bcconn_top_bl1[7] bcconn_top_bl1_n[7] bcconn_top_bl2[7] bcconn_top_bl2_n[7] DP8TVar9BulkConnRow_8
Xarray_bot vss vdd zero zero zero zero zero zero zero zero zero zero zero zero zero zero array_bot_bl1[0] array_bot_bl1_n[0] array_bot_bl2[0] array_bot_bl2_n[0] array_bot_bl1[1] array_bot_bl1_n[1] array_bot_bl2[1] array_bot_bl2_n[1] array_bot_bl1[2] array_bot_bl1_n[2] array_bot_bl2[2] array_bot_bl2_n[2] array_bot_bl1[3] array_bot_bl1_n[3] array_bot_bl2[3] array_bot_bl2_n[3] bl1 bl1_n bl2 bl2_n array_bot_bl1[5] array_bot_bl1_n[5] array_bot_bl2[5] array_bot_bl2_n[5] array_bot_bl1[6] array_bot_bl1_n[6] array_bot_bl2[6] array_bot_bl2_n[6] array_bot_bl1[7] array_bot_bl1_n[7] array_bot_bl2[7] array_bot_bl2_n[7] DP8TVar9Array_7X8
Xshwl1_row vss vdd zero bit shwl1_row_bl1[0] shwl1_row_bl1_n[0] shwl1_row_bl2[0] shwl1_row_bl2_n[0] shwl1_row_bl1[1] shwl1_row_bl1_n[1] shwl1_row_bl2[1] shwl1_row_bl2_n[1] shwl1_row_bl1[2] shwl1_row_bl1_n[2] shwl1_row_bl2[2] shwl1_row_bl2_n[2] shwl1_row_bl1[3] shwl1_row_bl1_n[3] shwl1_row_bl2[3] shwl1_row_bl2_n[3] bl1 bl1_n bl2 bl2_n shwl1_row_bl1[5] shwl1_row_bl1_n[5] shwl1_row_bl2[5] shwl1_row_bl2_n[5] shwl1_row_bl1[6] shwl1_row_bl1_n[6] shwl1_row_bl2[6] shwl1_row_bl2_n[6] shwl1_row_bl1[7] shwl1_row_bl1_n[7] shwl1_row_bl2[7] shwl1_row_bl2_n[7] DP8TVar9ArrayShWL1_1X8
Xcell_cols_left vss vdd wl1 wl2 cell_cols_left_bl1[0] cell_cols_left_bl1_n[0] cell_cols_left_bl2[0] cell_cols_left_bl2_n[0] cell_cols_left_bl1[1] cell_cols_left_bl1_n[1] cell_cols_left_bl2[1] cell_cols_left_bl2_n[1] cell_cols_left_bl1[2] cell_cols_left_bl1_n[2] cell_cols_left_bl2[2] cell_cols_left_bl2_n[2] cell_cols_left_bl1[3] cell_cols_left_bl1_n[3] cell_cols_left_bl2[3] cell_cols_left_bl2_n[3] DP8TVar9Array_1X4
Xconncell wl1 wl2 bl1 bl1_n bl2 bl2_n vdd vss bit bit_n DP8TVar9CellConnectOut
Xfillcell wl1 wl2 fillcell_bl1 fillcell_bl1_n fillcell_bl2 fillcell_bl2_n vdd vss DP8TVar9Cell
Xcell_cols_right vss vdd wl1 wl2 cell_cols_right_bl1[0] cell_cols_right_bl1_n[0] cell_cols_right_bl2[0] cell_cols_right_bl2_n[0] cell_cols_right_bl1[1] cell_cols_right_bl1_n[1] cell_cols_right_bl2[1] cell_cols_right_bl2_n[1] DP8TVar9Array_1X2
Xshwl2_row vss vdd bit_n zero shwl2_row_bl1[0] shwl2_row_bl1_n[0] shwl2_row_bl2[0] shwl2_row_bl2_n[0] shwl2_row_bl1[1] shwl2_row_bl1_n[1] shwl2_row_bl2[1] shwl2_row_bl2_n[1] shwl2_row_bl1[2] shwl2_row_bl1_n[2] shwl2_row_bl2[2] shwl2_row_bl2_n[2] shwl2_row_bl1[3] shwl2_row_bl1_n[3] shwl2_row_bl2[3] shwl2_row_bl2_n[3] bl1 bl1_n bl2 bl2_n shwl2_row_bl1[5] shwl2_row_bl1_n[5] shwl2_row_bl2[5] shwl2_row_bl2_n[5] shwl2_row_bl1[6] shwl2_row_bl1_n[6] shwl2_row_bl2[6] shwl2_row_bl2_n[6] shwl2_row_bl1[7] shwl2_row_bl1_n[7] shwl2_row_bl2[7] shwl2_row_bl2_n[7] DP8TVar9ArrayShWL2_1X8
Xarray_top vss vdd zero zero zero zero zero zero zero zero zero zero zero zero array_top_bl1[0] array_top_bl1_n[0] array_top_bl2[0] array_top_bl2_n[0] array_top_bl1[1] array_top_bl1_n[1] array_top_bl2[1] array_top_bl2_n[1] array_top_bl1[2] array_top_bl1_n[2] array_top_bl2[2] array_top_bl2_n[2] array_top_bl1[3] array_top_bl1_n[3] array_top_bl2[3] array_top_bl2_n[3] bl1 bl1_n bl2 bl2_n array_top_bl1[5] array_top_bl1_n[5] array_top_bl2[5] array_top_bl2_n[5] array_top_bl1[6] array_top_bl1_n[6] array_top_bl2[6] array_top_bl2_n[6] array_top_bl1[7] array_top_bl1_n[7] array_top_bl2[7] array_top_bl2_n[7] DP8TVar9Array_6X8
Xzero vdd vss zero zero_x1
.ends DP8TVar9TestArray_16X8C

.subckt DP8TVar9 vss noco_vdd noco_wl1 noco_wl2 noco_bl1 noco_bl1_n noco_bl2 noco_bl2_n co_vdd co_bit co_bit_n co_wl1 co_wl2 co_bl1 co_bl1_n co_bl2_n co_bl2
Xframe noco_vdd noco_wl1 noco_wl2 noco_bl2 co_vdd co_bit co_bit_n co_wl1 co_wl2 NoConn_PAD0x9 vss noco_bl1 noco_bl1_n noco_bl2_n vss co_bl1 co_bl1_n co_bl2_n co_bl2 NoConn_PAD1x9 PadFrame_DP09
Xtestarray_noco vss noco_vdd noco_wl1 noco_wl2 noco_bl1 noco_bl1_n noco_bl2 noco_bl2_n DP8TVar9TestArray_16X8
Xtestarray_co vss co_vdd co_wl1 co_wl2 co_bl1 co_bl1_n co_bl2 co_bl2_n co_bit co_bit_n DP8TVar9TestArray_16X8C
.ends DP8TVar9

.subckt PadFrame_DP10 PAD0x0 PAD0x1 PAD0x2 PAD0x3 PAD0x4 PAD0x5 PAD0x6 PAD0x7 PAD0x8 PAD0x9 PAD1x0 PAD1x1 PAD1x2 PAD1x3 PAD1x4 PAD1x5 PAD1x6 PAD1x7 PAD1x8 PAD1x9
XPAD0x0 PAD0x0 BondPad
XPAD0x1 PAD0x1 BondPad
XPAD0x2 PAD0x2 BondPad
XPAD0x3 PAD0x3 BondPad
XPAD0x4 PAD0x4 BondPad
XPAD0x5 PAD0x5 BondPad
XPAD0x6 PAD0x6 BondPad
XPAD0x7 PAD0x7 BondPad
XPAD0x8 PAD0x8 BondPad
XPAD0x9 PAD0x9 BondPad
XPAD1x0 PAD1x0 BondPad
XPAD1x1 PAD1x1 BondPad
XPAD1x2 PAD1x2 BondPad
XPAD1x3 PAD1x3 BondPad
XPAD1x4 PAD1x4 BondPad
XPAD1x5 PAD1x5 BondPad
XPAD1x6 PAD1x6 BondPad
XPAD1x7 PAD1x7 BondPad
XPAD1x8 PAD1x8 BondPad
XPAD1x9 PAD1x9 BondPad
.ends PadFrame_DP10

.subckt DP8TVar10Cell wl1 wl2 bl1 bl1_n bl2 bl2_n vdd vss
Xpu1 vdd bit_n bit vdd sg13_lv_pmos l=1.3e-07 w=2e-07
Xpd1 bit bit_n vss vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpu2 vdd bit bit_n vdd sg13_lv_pmos l=1.3e-07 w=2e-07
Xpd2 bit_n bit vss vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg1 bit wl1 bl1 vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg1n bit_n wl1 bl1_n vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg2 bit wl2 bl2 vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg2n bit_n wl2 bl2_n vss sg13_lv_nmos l=1.3e-07 w=2e-07
.ends DP8TVar10Cell

.subckt DP8TVar10Array_2X1 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0]
Xinst0x0 wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] vdd vss DP8TVar10Cell
Xinst1x0 wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0] vdd vss DP8TVar10Cell
.ends DP8TVar10Array_2X1

.subckt DP8TVar10Array_2X2 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0] DP8TVar10Array_2X1
Xinst0x1 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TVar10Array_2X1
.ends DP8TVar10Array_2X2

.subckt DP8TVar10Array_4X2 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TVar10Array_2X2
Xinst1x0 vss vdd wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TVar10Array_2X2
.ends DP8TVar10Array_4X2

.subckt DP8TVar10Array_4X4 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TVar10Array_4X2
Xinst0x1 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar10Array_4X2
.ends DP8TVar10Array_4X4

.subckt DP8TVar10Array_8X4 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar10Array_4X4
Xinst1x0 vss vdd wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar10Array_4X4
.ends DP8TVar10Array_8X4

.subckt DP8TVar10Array_8X8 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar10Array_8X4
Xinst0x1 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar10Array_8X4
.ends DP8TVar10Array_8X8

.subckt DP8TVar10BulkConn vdd vss bl1 bl2 bl1_n bl2_n
.ends DP8TVar10BulkConn

.subckt DP8TVar10BulkConnRow_2 vss vdd bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1]
Xinst0 vdd vss bl1[0] bl2[0] bl1_n[0] bl2_n[0] DP8TVar10BulkConn
Xinst1 vdd vss bl1[1] bl2[1] bl1_n[1] bl2_n[1] DP8TVar10BulkConn
.ends DP8TVar10BulkConnRow_2

.subckt DP8TVar10BulkConnRow_4 vss vdd bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3]
Xinst0 vss vdd bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TVar10BulkConnRow_2
Xinst1 vss vdd bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar10BulkConnRow_2
.ends DP8TVar10BulkConnRow_4

.subckt DP8TVar10BulkConnRow_8 vss vdd bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0 vss vdd bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar10BulkConnRow_4
Xinst1 vss vdd bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar10BulkConnRow_4
.ends DP8TVar10BulkConnRow_8

.subckt DP8TVar10Array_16X8BC vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] wl1[8] wl2[8] wl1[9] wl2[9] wl1[10] wl2[10] wl1[11] wl2[11] wl1[12] wl2[12] wl1[13] wl2[13] wl1[14] wl2[14] wl1[15] wl2[15] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar10Array_8X8
Xinst1x0 vss vdd wl1[8] wl2[8] wl1[9] wl2[9] wl1[10] wl2[10] wl1[11] wl2[11] wl1[12] wl2[12] wl1[13] wl2[13] wl1[14] wl2[14] wl1[15] wl2[15] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar10Array_8X8
Xbottombcrow vss vdd bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar10BulkConnRow_8
Xtopbcrow vss vdd bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar10BulkConnRow_8
.ends DP8TVar10Array_16X8BC

.subckt DP8TVar10TestArray_16X8 vss vdd wl1 wl2 bl1 bl1_n bl2 bl2_n
Xarray vss vdd zero zero zero zero zero zero zero zero zero zero zero zero zero zero zero zero wl1 wl2 zero zero zero zero zero zero zero zero zero zero zero zero zero zero bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1 bl1_n bl2 bl2_n bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar10Array_16X8BC
Xzero vdd vss zero zero_x1
.ends DP8TVar10TestArray_16X8

.subckt DP8TVar10Array_4X8 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar10Array_4X4
Xinst0x1 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar10Array_4X4
.ends DP8TVar10Array_4X8

.subckt DP8TVar10Array_2X4 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TVar10Array_2X2
Xinst0x1 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar10Array_2X2
.ends DP8TVar10Array_2X4

.subckt DP8TVar10Array_2X8 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar10Array_2X4
Xinst0x1 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar10Array_2X4
.ends DP8TVar10Array_2X8

.subckt DP8TVar10Array_1X2 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1]
Xinst0x0 wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] vdd vss DP8TVar10Cell
Xinst0x1 wl1[0] wl2[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] vdd vss DP8TVar10Cell
.ends DP8TVar10Array_1X2

.subckt DP8TVar10Array_1X4 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3]
Xinst0x0 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TVar10Array_1X2
Xinst0x1 vss vdd wl1[0] wl2[0] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar10Array_1X2
.ends DP8TVar10Array_1X4

.subckt DP8TVar10Array_1X8 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar10Array_1X4
Xinst0x1 vss vdd wl1[0] wl2[0] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar10Array_1X4
.ends DP8TVar10Array_1X8

.subckt DP8TVar10Array_7X8 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar10Array_4X8
Xinst1x0 vss vdd wl1[4] wl2[4] wl1[5] wl2[5] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar10Array_2X8
Xinst2x0 vss vdd wl1[6] wl2[6] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar10Array_1X8
.ends DP8TVar10Array_7X8

.subckt DP8TVar10CellShWL1 wl1 wl2 bl1 bl1_n bl2 bl2_n vdd vss
Xpu1 vdd bit_n bit vdd sg13_lv_pmos l=1.3e-07 w=2e-07
Xpd1 bit bit_n vss vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpu2 vdd bit bit_n vdd sg13_lv_pmos l=1.3e-07 w=2e-07
Xpd2 bit_n bit vss vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg1 bit wl1 bl1 vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg1n bit_n wl1 bl1_n vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg2 bit wl1 bl2 vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg2n bit_n wl1 bl2_n vss sg13_lv_nmos l=1.3e-07 w=2e-07
.ends DP8TVar10CellShWL1

.subckt DP8TVar10ArrayShWL1_1X2 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1]
Xinst0x0 wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] vdd vss DP8TVar10CellShWL1
Xinst0x1 wl1[0] wl2[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] vdd vss DP8TVar10CellShWL1
.ends DP8TVar10ArrayShWL1_1X2

.subckt DP8TVar10ArrayShWL1_1X4 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3]
Xinst0x0 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TVar10ArrayShWL1_1X2
Xinst0x1 vss vdd wl1[0] wl2[0] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar10ArrayShWL1_1X2
.ends DP8TVar10ArrayShWL1_1X4

.subckt DP8TVar10ArrayShWL1_1X8 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar10ArrayShWL1_1X4
Xinst0x1 vss vdd wl1[0] wl2[0] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar10ArrayShWL1_1X4
.ends DP8TVar10ArrayShWL1_1X8

.subckt DP8TVar10CellConnectOut wl1 wl2 bl1 bl1_n bl2 bl2_n vdd vss bit bit_n
Xpu1 vdd bit_n bit vdd sg13_lv_pmos l=1.3e-07 w=2e-07
Xpd1 bit bit_n vss vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpu2 vdd bit bit_n vdd sg13_lv_pmos l=1.3e-07 w=2e-07
Xpd2 bit_n bit vss vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg1 bit wl1 bl1 vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg1n bit_n wl1 bl1_n vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg2 bit wl2 bl2 vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg2n bit_n wl2 bl2_n vss sg13_lv_nmos l=1.3e-07 w=2e-07
.ends DP8TVar10CellConnectOut

.subckt DP8TVar10CellShWL2 wl1 wl2 bl1 bl1_n bl2 bl2_n vdd vss
Xpu1 vdd bit_n bit vdd sg13_lv_pmos l=1.3e-07 w=2e-07
Xpd1 bit bit_n vss vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpu2 vdd bit bit_n vdd sg13_lv_pmos l=1.3e-07 w=2e-07
Xpd2 bit_n bit vss vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg1 bit wl2 bl1 vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg1n bit_n wl2 bl1_n vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg2 bit wl2 bl2 vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg2n bit_n wl2 bl2_n vss sg13_lv_nmos l=1.3e-07 w=2e-07
.ends DP8TVar10CellShWL2

.subckt DP8TVar10ArrayShWL2_1X2 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1]
Xinst0x0 wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] vdd vss DP8TVar10CellShWL2
Xinst0x1 wl1[0] wl2[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] vdd vss DP8TVar10CellShWL2
.ends DP8TVar10ArrayShWL2_1X2

.subckt DP8TVar10ArrayShWL2_1X4 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3]
Xinst0x0 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TVar10ArrayShWL2_1X2
Xinst0x1 vss vdd wl1[0] wl2[0] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar10ArrayShWL2_1X2
.ends DP8TVar10ArrayShWL2_1X4

.subckt DP8TVar10ArrayShWL2_1X8 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar10ArrayShWL2_1X4
Xinst0x1 vss vdd wl1[0] wl2[0] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar10ArrayShWL2_1X4
.ends DP8TVar10ArrayShWL2_1X8

.subckt DP8TVar10Array_6X8 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar10Array_4X8
Xinst1x0 vss vdd wl1[4] wl2[4] wl1[5] wl2[5] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar10Array_2X8
.ends DP8TVar10Array_6X8

.subckt DP8TVar10TestArray_16X8C vss vdd wl1 wl2 bl1 bl1_n bl2 bl2_n bit bit_n
Xbcconn_bot vss vdd bcconn_bot_bl1[0] bcconn_bot_bl1_n[0] bcconn_bot_bl2[0] bcconn_bot_bl2_n[0] bcconn_bot_bl1[1] bcconn_bot_bl1_n[1] bcconn_bot_bl2[1] bcconn_bot_bl2_n[1] bcconn_bot_bl1[2] bcconn_bot_bl1_n[2] bcconn_bot_bl2[2] bcconn_bot_bl2_n[2] bcconn_bot_bl1[3] bcconn_bot_bl1_n[3] bcconn_bot_bl2[3] bcconn_bot_bl2_n[3] bl1 bl1_n bl2 bl2_n bcconn_bot_bl1[5] bcconn_bot_bl1_n[5] bcconn_bot_bl2[5] bcconn_bot_bl2_n[5] bcconn_bot_bl1[6] bcconn_bot_bl1_n[6] bcconn_bot_bl2[6] bcconn_bot_bl2_n[6] bcconn_bot_bl1[7] bcconn_bot_bl1_n[7] bcconn_bot_bl2[7] bcconn_bot_bl2_n[7] DP8TVar10BulkConnRow_8
Xbcconn_top vss vdd bcconn_top_bl1[0] bcconn_top_bl1_n[0] bcconn_top_bl2[0] bcconn_top_bl2_n[0] bcconn_top_bl1[1] bcconn_top_bl1_n[1] bcconn_top_bl2[1] bcconn_top_bl2_n[1] bcconn_top_bl1[2] bcconn_top_bl1_n[2] bcconn_top_bl2[2] bcconn_top_bl2_n[2] bcconn_top_bl1[3] bcconn_top_bl1_n[3] bcconn_top_bl2[3] bcconn_top_bl2_n[3] bl1 bl1_n bl2 bl2_n bcconn_top_bl1[5] bcconn_top_bl1_n[5] bcconn_top_bl2[5] bcconn_top_bl2_n[5] bcconn_top_bl1[6] bcconn_top_bl1_n[6] bcconn_top_bl2[6] bcconn_top_bl2_n[6] bcconn_top_bl1[7] bcconn_top_bl1_n[7] bcconn_top_bl2[7] bcconn_top_bl2_n[7] DP8TVar10BulkConnRow_8
Xarray_bot vss vdd zero zero zero zero zero zero zero zero zero zero zero zero zero zero array_bot_bl1[0] array_bot_bl1_n[0] array_bot_bl2[0] array_bot_bl2_n[0] array_bot_bl1[1] array_bot_bl1_n[1] array_bot_bl2[1] array_bot_bl2_n[1] array_bot_bl1[2] array_bot_bl1_n[2] array_bot_bl2[2] array_bot_bl2_n[2] array_bot_bl1[3] array_bot_bl1_n[3] array_bot_bl2[3] array_bot_bl2_n[3] bl1 bl1_n bl2 bl2_n array_bot_bl1[5] array_bot_bl1_n[5] array_bot_bl2[5] array_bot_bl2_n[5] array_bot_bl1[6] array_bot_bl1_n[6] array_bot_bl2[6] array_bot_bl2_n[6] array_bot_bl1[7] array_bot_bl1_n[7] array_bot_bl2[7] array_bot_bl2_n[7] DP8TVar10Array_7X8
Xshwl1_row vss vdd zero bit shwl1_row_bl1[0] shwl1_row_bl1_n[0] shwl1_row_bl2[0] shwl1_row_bl2_n[0] shwl1_row_bl1[1] shwl1_row_bl1_n[1] shwl1_row_bl2[1] shwl1_row_bl2_n[1] shwl1_row_bl1[2] shwl1_row_bl1_n[2] shwl1_row_bl2[2] shwl1_row_bl2_n[2] shwl1_row_bl1[3] shwl1_row_bl1_n[3] shwl1_row_bl2[3] shwl1_row_bl2_n[3] bl1 bl1_n bl2 bl2_n shwl1_row_bl1[5] shwl1_row_bl1_n[5] shwl1_row_bl2[5] shwl1_row_bl2_n[5] shwl1_row_bl1[6] shwl1_row_bl1_n[6] shwl1_row_bl2[6] shwl1_row_bl2_n[6] shwl1_row_bl1[7] shwl1_row_bl1_n[7] shwl1_row_bl2[7] shwl1_row_bl2_n[7] DP8TVar10ArrayShWL1_1X8
Xcell_cols_left vss vdd wl1 wl2 cell_cols_left_bl1[0] cell_cols_left_bl1_n[0] cell_cols_left_bl2[0] cell_cols_left_bl2_n[0] cell_cols_left_bl1[1] cell_cols_left_bl1_n[1] cell_cols_left_bl2[1] cell_cols_left_bl2_n[1] cell_cols_left_bl1[2] cell_cols_left_bl1_n[2] cell_cols_left_bl2[2] cell_cols_left_bl2_n[2] cell_cols_left_bl1[3] cell_cols_left_bl1_n[3] cell_cols_left_bl2[3] cell_cols_left_bl2_n[3] DP8TVar10Array_1X4
Xconncell wl1 wl2 bl1 bl1_n bl2 bl2_n vdd vss bit bit_n DP8TVar10CellConnectOut
Xfillcell wl1 wl2 fillcell_bl1 fillcell_bl1_n fillcell_bl2 fillcell_bl2_n vdd vss DP8TVar10Cell
Xcell_cols_right vss vdd wl1 wl2 cell_cols_right_bl1[0] cell_cols_right_bl1_n[0] cell_cols_right_bl2[0] cell_cols_right_bl2_n[0] cell_cols_right_bl1[1] cell_cols_right_bl1_n[1] cell_cols_right_bl2[1] cell_cols_right_bl2_n[1] DP8TVar10Array_1X2
Xshwl2_row vss vdd bit_n zero shwl2_row_bl1[0] shwl2_row_bl1_n[0] shwl2_row_bl2[0] shwl2_row_bl2_n[0] shwl2_row_bl1[1] shwl2_row_bl1_n[1] shwl2_row_bl2[1] shwl2_row_bl2_n[1] shwl2_row_bl1[2] shwl2_row_bl1_n[2] shwl2_row_bl2[2] shwl2_row_bl2_n[2] shwl2_row_bl1[3] shwl2_row_bl1_n[3] shwl2_row_bl2[3] shwl2_row_bl2_n[3] bl1 bl1_n bl2 bl2_n shwl2_row_bl1[5] shwl2_row_bl1_n[5] shwl2_row_bl2[5] shwl2_row_bl2_n[5] shwl2_row_bl1[6] shwl2_row_bl1_n[6] shwl2_row_bl2[6] shwl2_row_bl2_n[6] shwl2_row_bl1[7] shwl2_row_bl1_n[7] shwl2_row_bl2[7] shwl2_row_bl2_n[7] DP8TVar10ArrayShWL2_1X8
Xarray_top vss vdd zero zero zero zero zero zero zero zero zero zero zero zero array_top_bl1[0] array_top_bl1_n[0] array_top_bl2[0] array_top_bl2_n[0] array_top_bl1[1] array_top_bl1_n[1] array_top_bl2[1] array_top_bl2_n[1] array_top_bl1[2] array_top_bl1_n[2] array_top_bl2[2] array_top_bl2_n[2] array_top_bl1[3] array_top_bl1_n[3] array_top_bl2[3] array_top_bl2_n[3] bl1 bl1_n bl2 bl2_n array_top_bl1[5] array_top_bl1_n[5] array_top_bl2[5] array_top_bl2_n[5] array_top_bl1[6] array_top_bl1_n[6] array_top_bl2[6] array_top_bl2_n[6] array_top_bl1[7] array_top_bl1_n[7] array_top_bl2[7] array_top_bl2_n[7] DP8TVar10Array_6X8
Xzero vdd vss zero zero_x1
.ends DP8TVar10TestArray_16X8C

.subckt DP8TVar10 vss noco_vdd noco_wl1 noco_wl2 noco_bl1 noco_bl1_n noco_bl2 noco_bl2_n co_vdd co_bit co_bit_n co_wl1 co_wl2 co_bl1 co_bl1_n co_bl2_n co_bl2
Xframe noco_vdd noco_wl1 noco_wl2 noco_bl2 co_vdd co_bit co_bit_n co_wl1 co_wl2 NoConn_PAD0x9 vss noco_bl1 noco_bl1_n noco_bl2_n vss co_bl1 co_bl1_n co_bl2_n co_bl2 NoConn_PAD1x9 PadFrame_DP10
Xtestarray_noco vss noco_vdd noco_wl1 noco_wl2 noco_bl1 noco_bl1_n noco_bl2 noco_bl2_n DP8TVar10TestArray_16X8
Xtestarray_co vss co_vdd co_wl1 co_wl2 co_bl1 co_bl1_n co_bl2 co_bl2_n co_bit co_bit_n DP8TVar10TestArray_16X8C
.ends DP8TVar10

.subckt PadFrame_DP11 PAD0x0 PAD0x1 PAD0x2 PAD0x3 PAD0x4 PAD0x5 PAD0x6 PAD0x7 PAD0x8 PAD0x9 PAD1x0 PAD1x1 PAD1x2 PAD1x3 PAD1x4 PAD1x5 PAD1x6 PAD1x7 PAD1x8 PAD1x9
XPAD0x0 PAD0x0 BondPad
XPAD0x1 PAD0x1 BondPad
XPAD0x2 PAD0x2 BondPad
XPAD0x3 PAD0x3 BondPad
XPAD0x4 PAD0x4 BondPad
XPAD0x5 PAD0x5 BondPad
XPAD0x6 PAD0x6 BondPad
XPAD0x7 PAD0x7 BondPad
XPAD0x8 PAD0x8 BondPad
XPAD0x9 PAD0x9 BondPad
XPAD1x0 PAD1x0 BondPad
XPAD1x1 PAD1x1 BondPad
XPAD1x2 PAD1x2 BondPad
XPAD1x3 PAD1x3 BondPad
XPAD1x4 PAD1x4 BondPad
XPAD1x5 PAD1x5 BondPad
XPAD1x6 PAD1x6 BondPad
XPAD1x7 PAD1x7 BondPad
XPAD1x8 PAD1x8 BondPad
XPAD1x9 PAD1x9 BondPad
.ends PadFrame_DP11

.subckt DP8TVar11Cell wl1 wl2 bl1 bl1_n bl2 bl2_n vdd vss
Xpu1 vdd bit_n bit vdd sg13_lv_pmos l=1.3e-07 w=1.5e-07
Xpd1 bit bit_n vss vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpu2 vdd bit bit_n vdd sg13_lv_pmos l=1.3e-07 w=1.5e-07
Xpd2 bit_n bit vss vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg1 bit wl1 bl1 vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg1n bit_n wl1 bl1_n vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg2 bit wl2 bl2 vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg2n bit_n wl2 bl2_n vss sg13_lv_nmos l=1.3e-07 w=2e-07
.ends DP8TVar11Cell

.subckt DP8TVar11Array_2X1 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0]
Xinst0x0 wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] vdd vss DP8TVar11Cell
Xinst1x0 wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0] vdd vss DP8TVar11Cell
.ends DP8TVar11Array_2X1

.subckt DP8TVar11Array_2X2 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0] DP8TVar11Array_2X1
Xinst0x1 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TVar11Array_2X1
.ends DP8TVar11Array_2X2

.subckt DP8TVar11Array_4X2 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TVar11Array_2X2
Xinst1x0 vss vdd wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TVar11Array_2X2
.ends DP8TVar11Array_4X2

.subckt DP8TVar11Array_4X4 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TVar11Array_4X2
Xinst0x1 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar11Array_4X2
.ends DP8TVar11Array_4X4

.subckt DP8TVar11Array_8X4 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar11Array_4X4
Xinst1x0 vss vdd wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar11Array_4X4
.ends DP8TVar11Array_8X4

.subckt DP8TVar11Array_8X8 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar11Array_8X4
Xinst0x1 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar11Array_8X4
.ends DP8TVar11Array_8X8

.subckt DP8TVar11BulkConn vdd vss bl1 bl2 bl1_n bl2_n
.ends DP8TVar11BulkConn

.subckt DP8TVar11BulkConnRow_2 vss vdd bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1]
Xinst0 vdd vss bl1[0] bl2[0] bl1_n[0] bl2_n[0] DP8TVar11BulkConn
Xinst1 vdd vss bl1[1] bl2[1] bl1_n[1] bl2_n[1] DP8TVar11BulkConn
.ends DP8TVar11BulkConnRow_2

.subckt DP8TVar11BulkConnRow_4 vss vdd bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3]
Xinst0 vss vdd bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TVar11BulkConnRow_2
Xinst1 vss vdd bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar11BulkConnRow_2
.ends DP8TVar11BulkConnRow_4

.subckt DP8TVar11BulkConnRow_8 vss vdd bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0 vss vdd bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar11BulkConnRow_4
Xinst1 vss vdd bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar11BulkConnRow_4
.ends DP8TVar11BulkConnRow_8

.subckt DP8TVar11Array_16X8BC vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] wl1[8] wl2[8] wl1[9] wl2[9] wl1[10] wl2[10] wl1[11] wl2[11] wl1[12] wl2[12] wl1[13] wl2[13] wl1[14] wl2[14] wl1[15] wl2[15] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar11Array_8X8
Xinst1x0 vss vdd wl1[8] wl2[8] wl1[9] wl2[9] wl1[10] wl2[10] wl1[11] wl2[11] wl1[12] wl2[12] wl1[13] wl2[13] wl1[14] wl2[14] wl1[15] wl2[15] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar11Array_8X8
Xbottombcrow vss vdd bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar11BulkConnRow_8
Xtopbcrow vss vdd bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar11BulkConnRow_8
.ends DP8TVar11Array_16X8BC

.subckt DP8TVar11TestArray_16X8 vss vdd wl1 wl2 bl1 bl1_n bl2 bl2_n
Xarray vss vdd zero zero zero zero zero zero zero zero zero zero zero zero zero zero zero zero wl1 wl2 zero zero zero zero zero zero zero zero zero zero zero zero zero zero bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1 bl1_n bl2 bl2_n bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar11Array_16X8BC
Xzero vdd vss zero zero_x1
.ends DP8TVar11TestArray_16X8

.subckt DP8TVar11Array_4X8 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar11Array_4X4
Xinst0x1 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar11Array_4X4
.ends DP8TVar11Array_4X8

.subckt DP8TVar11Array_2X4 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TVar11Array_2X2
Xinst0x1 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar11Array_2X2
.ends DP8TVar11Array_2X4

.subckt DP8TVar11Array_2X8 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar11Array_2X4
Xinst0x1 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar11Array_2X4
.ends DP8TVar11Array_2X8

.subckt DP8TVar11Array_1X2 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1]
Xinst0x0 wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] vdd vss DP8TVar11Cell
Xinst0x1 wl1[0] wl2[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] vdd vss DP8TVar11Cell
.ends DP8TVar11Array_1X2

.subckt DP8TVar11Array_1X4 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3]
Xinst0x0 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TVar11Array_1X2
Xinst0x1 vss vdd wl1[0] wl2[0] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar11Array_1X2
.ends DP8TVar11Array_1X4

.subckt DP8TVar11Array_1X8 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar11Array_1X4
Xinst0x1 vss vdd wl1[0] wl2[0] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar11Array_1X4
.ends DP8TVar11Array_1X8

.subckt DP8TVar11Array_7X8 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar11Array_4X8
Xinst1x0 vss vdd wl1[4] wl2[4] wl1[5] wl2[5] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar11Array_2X8
Xinst2x0 vss vdd wl1[6] wl2[6] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar11Array_1X8
.ends DP8TVar11Array_7X8

.subckt DP8TVar11CellShWL1 wl1 wl2 bl1 bl1_n bl2 bl2_n vdd vss
Xpu1 vdd bit_n bit vdd sg13_lv_pmos l=1.3e-07 w=1.5e-07
Xpd1 bit bit_n vss vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpu2 vdd bit bit_n vdd sg13_lv_pmos l=1.3e-07 w=1.5e-07
Xpd2 bit_n bit vss vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg1 bit wl1 bl1 vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg1n bit_n wl1 bl1_n vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg2 bit wl1 bl2 vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg2n bit_n wl1 bl2_n vss sg13_lv_nmos l=1.3e-07 w=2e-07
.ends DP8TVar11CellShWL1

.subckt DP8TVar11ArrayShWL1_1X2 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1]
Xinst0x0 wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] vdd vss DP8TVar11CellShWL1
Xinst0x1 wl1[0] wl2[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] vdd vss DP8TVar11CellShWL1
.ends DP8TVar11ArrayShWL1_1X2

.subckt DP8TVar11ArrayShWL1_1X4 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3]
Xinst0x0 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TVar11ArrayShWL1_1X2
Xinst0x1 vss vdd wl1[0] wl2[0] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar11ArrayShWL1_1X2
.ends DP8TVar11ArrayShWL1_1X4

.subckt DP8TVar11ArrayShWL1_1X8 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar11ArrayShWL1_1X4
Xinst0x1 vss vdd wl1[0] wl2[0] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar11ArrayShWL1_1X4
.ends DP8TVar11ArrayShWL1_1X8

.subckt DP8TVar11CellConnectOut wl1 wl2 bl1 bl1_n bl2 bl2_n vdd vss bit bit_n
Xpu1 vdd bit_n bit vdd sg13_lv_pmos l=1.3e-07 w=1.5e-07
Xpd1 bit bit_n vss vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpu2 vdd bit bit_n vdd sg13_lv_pmos l=1.3e-07 w=1.5e-07
Xpd2 bit_n bit vss vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg1 bit wl1 bl1 vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg1n bit_n wl1 bl1_n vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg2 bit wl2 bl2 vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg2n bit_n wl2 bl2_n vss sg13_lv_nmos l=1.3e-07 w=2e-07
.ends DP8TVar11CellConnectOut

.subckt DP8TVar11CellShWL2 wl1 wl2 bl1 bl1_n bl2 bl2_n vdd vss
Xpu1 vdd bit_n bit vdd sg13_lv_pmos l=1.3e-07 w=1.5e-07
Xpd1 bit bit_n vss vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpu2 vdd bit bit_n vdd sg13_lv_pmos l=1.3e-07 w=1.5e-07
Xpd2 bit_n bit vss vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg1 bit wl2 bl1 vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg1n bit_n wl2 bl1_n vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg2 bit wl2 bl2 vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg2n bit_n wl2 bl2_n vss sg13_lv_nmos l=1.3e-07 w=2e-07
.ends DP8TVar11CellShWL2

.subckt DP8TVar11ArrayShWL2_1X2 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1]
Xinst0x0 wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] vdd vss DP8TVar11CellShWL2
Xinst0x1 wl1[0] wl2[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] vdd vss DP8TVar11CellShWL2
.ends DP8TVar11ArrayShWL2_1X2

.subckt DP8TVar11ArrayShWL2_1X4 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3]
Xinst0x0 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TVar11ArrayShWL2_1X2
Xinst0x1 vss vdd wl1[0] wl2[0] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar11ArrayShWL2_1X2
.ends DP8TVar11ArrayShWL2_1X4

.subckt DP8TVar11ArrayShWL2_1X8 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar11ArrayShWL2_1X4
Xinst0x1 vss vdd wl1[0] wl2[0] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar11ArrayShWL2_1X4
.ends DP8TVar11ArrayShWL2_1X8

.subckt DP8TVar11Array_6X8 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar11Array_4X8
Xinst1x0 vss vdd wl1[4] wl2[4] wl1[5] wl2[5] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar11Array_2X8
.ends DP8TVar11Array_6X8

.subckt DP8TVar11TestArray_16X8C vss vdd wl1 wl2 bl1 bl1_n bl2 bl2_n bit bit_n
Xbcconn_bot vss vdd bcconn_bot_bl1[0] bcconn_bot_bl1_n[0] bcconn_bot_bl2[0] bcconn_bot_bl2_n[0] bcconn_bot_bl1[1] bcconn_bot_bl1_n[1] bcconn_bot_bl2[1] bcconn_bot_bl2_n[1] bcconn_bot_bl1[2] bcconn_bot_bl1_n[2] bcconn_bot_bl2[2] bcconn_bot_bl2_n[2] bcconn_bot_bl1[3] bcconn_bot_bl1_n[3] bcconn_bot_bl2[3] bcconn_bot_bl2_n[3] bl1 bl1_n bl2 bl2_n bcconn_bot_bl1[5] bcconn_bot_bl1_n[5] bcconn_bot_bl2[5] bcconn_bot_bl2_n[5] bcconn_bot_bl1[6] bcconn_bot_bl1_n[6] bcconn_bot_bl2[6] bcconn_bot_bl2_n[6] bcconn_bot_bl1[7] bcconn_bot_bl1_n[7] bcconn_bot_bl2[7] bcconn_bot_bl2_n[7] DP8TVar11BulkConnRow_8
Xbcconn_top vss vdd bcconn_top_bl1[0] bcconn_top_bl1_n[0] bcconn_top_bl2[0] bcconn_top_bl2_n[0] bcconn_top_bl1[1] bcconn_top_bl1_n[1] bcconn_top_bl2[1] bcconn_top_bl2_n[1] bcconn_top_bl1[2] bcconn_top_bl1_n[2] bcconn_top_bl2[2] bcconn_top_bl2_n[2] bcconn_top_bl1[3] bcconn_top_bl1_n[3] bcconn_top_bl2[3] bcconn_top_bl2_n[3] bl1 bl1_n bl2 bl2_n bcconn_top_bl1[5] bcconn_top_bl1_n[5] bcconn_top_bl2[5] bcconn_top_bl2_n[5] bcconn_top_bl1[6] bcconn_top_bl1_n[6] bcconn_top_bl2[6] bcconn_top_bl2_n[6] bcconn_top_bl1[7] bcconn_top_bl1_n[7] bcconn_top_bl2[7] bcconn_top_bl2_n[7] DP8TVar11BulkConnRow_8
Xarray_bot vss vdd zero zero zero zero zero zero zero zero zero zero zero zero zero zero array_bot_bl1[0] array_bot_bl1_n[0] array_bot_bl2[0] array_bot_bl2_n[0] array_bot_bl1[1] array_bot_bl1_n[1] array_bot_bl2[1] array_bot_bl2_n[1] array_bot_bl1[2] array_bot_bl1_n[2] array_bot_bl2[2] array_bot_bl2_n[2] array_bot_bl1[3] array_bot_bl1_n[3] array_bot_bl2[3] array_bot_bl2_n[3] bl1 bl1_n bl2 bl2_n array_bot_bl1[5] array_bot_bl1_n[5] array_bot_bl2[5] array_bot_bl2_n[5] array_bot_bl1[6] array_bot_bl1_n[6] array_bot_bl2[6] array_bot_bl2_n[6] array_bot_bl1[7] array_bot_bl1_n[7] array_bot_bl2[7] array_bot_bl2_n[7] DP8TVar11Array_7X8
Xshwl1_row vss vdd zero bit shwl1_row_bl1[0] shwl1_row_bl1_n[0] shwl1_row_bl2[0] shwl1_row_bl2_n[0] shwl1_row_bl1[1] shwl1_row_bl1_n[1] shwl1_row_bl2[1] shwl1_row_bl2_n[1] shwl1_row_bl1[2] shwl1_row_bl1_n[2] shwl1_row_bl2[2] shwl1_row_bl2_n[2] shwl1_row_bl1[3] shwl1_row_bl1_n[3] shwl1_row_bl2[3] shwl1_row_bl2_n[3] bl1 bl1_n bl2 bl2_n shwl1_row_bl1[5] shwl1_row_bl1_n[5] shwl1_row_bl2[5] shwl1_row_bl2_n[5] shwl1_row_bl1[6] shwl1_row_bl1_n[6] shwl1_row_bl2[6] shwl1_row_bl2_n[6] shwl1_row_bl1[7] shwl1_row_bl1_n[7] shwl1_row_bl2[7] shwl1_row_bl2_n[7] DP8TVar11ArrayShWL1_1X8
Xcell_cols_left vss vdd wl1 wl2 cell_cols_left_bl1[0] cell_cols_left_bl1_n[0] cell_cols_left_bl2[0] cell_cols_left_bl2_n[0] cell_cols_left_bl1[1] cell_cols_left_bl1_n[1] cell_cols_left_bl2[1] cell_cols_left_bl2_n[1] cell_cols_left_bl1[2] cell_cols_left_bl1_n[2] cell_cols_left_bl2[2] cell_cols_left_bl2_n[2] cell_cols_left_bl1[3] cell_cols_left_bl1_n[3] cell_cols_left_bl2[3] cell_cols_left_bl2_n[3] DP8TVar11Array_1X4
Xconncell wl1 wl2 bl1 bl1_n bl2 bl2_n vdd vss bit bit_n DP8TVar11CellConnectOut
Xfillcell wl1 wl2 fillcell_bl1 fillcell_bl1_n fillcell_bl2 fillcell_bl2_n vdd vss DP8TVar11Cell
Xcell_cols_right vss vdd wl1 wl2 cell_cols_right_bl1[0] cell_cols_right_bl1_n[0] cell_cols_right_bl2[0] cell_cols_right_bl2_n[0] cell_cols_right_bl1[1] cell_cols_right_bl1_n[1] cell_cols_right_bl2[1] cell_cols_right_bl2_n[1] DP8TVar11Array_1X2
Xshwl2_row vss vdd bit_n zero shwl2_row_bl1[0] shwl2_row_bl1_n[0] shwl2_row_bl2[0] shwl2_row_bl2_n[0] shwl2_row_bl1[1] shwl2_row_bl1_n[1] shwl2_row_bl2[1] shwl2_row_bl2_n[1] shwl2_row_bl1[2] shwl2_row_bl1_n[2] shwl2_row_bl2[2] shwl2_row_bl2_n[2] shwl2_row_bl1[3] shwl2_row_bl1_n[3] shwl2_row_bl2[3] shwl2_row_bl2_n[3] bl1 bl1_n bl2 bl2_n shwl2_row_bl1[5] shwl2_row_bl1_n[5] shwl2_row_bl2[5] shwl2_row_bl2_n[5] shwl2_row_bl1[6] shwl2_row_bl1_n[6] shwl2_row_bl2[6] shwl2_row_bl2_n[6] shwl2_row_bl1[7] shwl2_row_bl1_n[7] shwl2_row_bl2[7] shwl2_row_bl2_n[7] DP8TVar11ArrayShWL2_1X8
Xarray_top vss vdd zero zero zero zero zero zero zero zero zero zero zero zero array_top_bl1[0] array_top_bl1_n[0] array_top_bl2[0] array_top_bl2_n[0] array_top_bl1[1] array_top_bl1_n[1] array_top_bl2[1] array_top_bl2_n[1] array_top_bl1[2] array_top_bl1_n[2] array_top_bl2[2] array_top_bl2_n[2] array_top_bl1[3] array_top_bl1_n[3] array_top_bl2[3] array_top_bl2_n[3] bl1 bl1_n bl2 bl2_n array_top_bl1[5] array_top_bl1_n[5] array_top_bl2[5] array_top_bl2_n[5] array_top_bl1[6] array_top_bl1_n[6] array_top_bl2[6] array_top_bl2_n[6] array_top_bl1[7] array_top_bl1_n[7] array_top_bl2[7] array_top_bl2_n[7] DP8TVar11Array_6X8
Xzero vdd vss zero zero_x1
.ends DP8TVar11TestArray_16X8C

.subckt DP8TVar11 vss noco_vdd noco_wl1 noco_wl2 noco_bl1 noco_bl1_n noco_bl2 noco_bl2_n co_vdd co_bit co_bit_n co_wl1 co_wl2 co_bl1 co_bl1_n co_bl2_n co_bl2
Xframe noco_vdd noco_wl1 noco_wl2 noco_bl2 co_vdd co_bit co_bit_n co_wl1 co_wl2 NoConn_PAD0x9 vss noco_bl1 noco_bl1_n noco_bl2_n vss co_bl1 co_bl1_n co_bl2_n co_bl2 NoConn_PAD1x9 PadFrame_DP11
Xtestarray_noco vss noco_vdd noco_wl1 noco_wl2 noco_bl1 noco_bl1_n noco_bl2 noco_bl2_n DP8TVar11TestArray_16X8
Xtestarray_co vss co_vdd co_wl1 co_wl2 co_bl1 co_bl1_n co_bl2 co_bl2_n co_bit co_bit_n DP8TVar11TestArray_16X8C
.ends DP8TVar11

.subckt PadFrame_DP12 PAD0x0 PAD0x1 PAD0x2 PAD0x3 PAD0x4 PAD0x5 PAD0x6 PAD0x7 PAD0x8 PAD0x9 PAD1x0 PAD1x1 PAD1x2 PAD1x3 PAD1x4 PAD1x5 PAD1x6 PAD1x7 PAD1x8 PAD1x9
XPAD0x0 PAD0x0 BondPad
XPAD0x1 PAD0x1 BondPad
XPAD0x2 PAD0x2 BondPad
XPAD0x3 PAD0x3 BondPad
XPAD0x4 PAD0x4 BondPad
XPAD0x5 PAD0x5 BondPad
XPAD0x6 PAD0x6 BondPad
XPAD0x7 PAD0x7 BondPad
XPAD0x8 PAD0x8 BondPad
XPAD0x9 PAD0x9 BondPad
XPAD1x0 PAD1x0 BondPad
XPAD1x1 PAD1x1 BondPad
XPAD1x2 PAD1x2 BondPad
XPAD1x3 PAD1x3 BondPad
XPAD1x4 PAD1x4 BondPad
XPAD1x5 PAD1x5 BondPad
XPAD1x6 PAD1x6 BondPad
XPAD1x7 PAD1x7 BondPad
XPAD1x8 PAD1x8 BondPad
XPAD1x9 PAD1x9 BondPad
.ends PadFrame_DP12

.subckt DP8TVar12Cell wl1 wl2 bl1 bl1_n bl2 bl2_n vdd vss
Xpu1 vdd bit_n bit vdd sg13_lv_pmos l=1.3e-07 w=2e-07
Xpd1 bit bit_n vss vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpu2 vdd bit bit_n vdd sg13_lv_pmos l=1.3e-07 w=2e-07
Xpd2 bit_n bit vss vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg1 bit wl1 bl1 vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg1n bit_n wl1 bl1_n vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg2 bit wl2 bl2 vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg2n bit_n wl2 bl2_n vss sg13_lv_nmos l=1.3e-07 w=2e-07
.ends DP8TVar12Cell

.subckt DP8TVar12Array_2X1 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0]
Xinst0x0 wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] vdd vss DP8TVar12Cell
Xinst1x0 wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0] vdd vss DP8TVar12Cell
.ends DP8TVar12Array_2X1

.subckt DP8TVar12Array_2X2 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0] DP8TVar12Array_2X1
Xinst0x1 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TVar12Array_2X1
.ends DP8TVar12Array_2X2

.subckt DP8TVar12Array_4X2 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TVar12Array_2X2
Xinst1x0 vss vdd wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TVar12Array_2X2
.ends DP8TVar12Array_4X2

.subckt DP8TVar12Array_4X4 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TVar12Array_4X2
Xinst0x1 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar12Array_4X2
.ends DP8TVar12Array_4X4

.subckt DP8TVar12Array_8X4 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar12Array_4X4
Xinst1x0 vss vdd wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar12Array_4X4
.ends DP8TVar12Array_8X4

.subckt DP8TVar12Array_8X8 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar12Array_8X4
Xinst0x1 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar12Array_8X4
.ends DP8TVar12Array_8X8

.subckt DP8TVar12BulkConn vdd vss bl1 bl2 bl1_n bl2_n
.ends DP8TVar12BulkConn

.subckt DP8TVar12BulkConnRow_2 vss vdd bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1]
Xinst0 vdd vss bl1[0] bl2[0] bl1_n[0] bl2_n[0] DP8TVar12BulkConn
Xinst1 vdd vss bl1[1] bl2[1] bl1_n[1] bl2_n[1] DP8TVar12BulkConn
.ends DP8TVar12BulkConnRow_2

.subckt DP8TVar12BulkConnRow_4 vss vdd bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3]
Xinst0 vss vdd bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TVar12BulkConnRow_2
Xinst1 vss vdd bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar12BulkConnRow_2
.ends DP8TVar12BulkConnRow_4

.subckt DP8TVar12BulkConnRow_8 vss vdd bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0 vss vdd bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar12BulkConnRow_4
Xinst1 vss vdd bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar12BulkConnRow_4
.ends DP8TVar12BulkConnRow_8

.subckt DP8TVar12Array_16X8BC vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] wl1[8] wl2[8] wl1[9] wl2[9] wl1[10] wl2[10] wl1[11] wl2[11] wl1[12] wl2[12] wl1[13] wl2[13] wl1[14] wl2[14] wl1[15] wl2[15] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar12Array_8X8
Xinst1x0 vss vdd wl1[8] wl2[8] wl1[9] wl2[9] wl1[10] wl2[10] wl1[11] wl2[11] wl1[12] wl2[12] wl1[13] wl2[13] wl1[14] wl2[14] wl1[15] wl2[15] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar12Array_8X8
Xbottombcrow vss vdd bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar12BulkConnRow_8
Xtopbcrow vss vdd bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar12BulkConnRow_8
.ends DP8TVar12Array_16X8BC

.subckt DP8TVar12TestArray_16X8 vss vdd wl1 wl2 bl1 bl1_n bl2 bl2_n
Xarray vss vdd zero zero zero zero zero zero zero zero zero zero zero zero zero zero zero zero wl1 wl2 zero zero zero zero zero zero zero zero zero zero zero zero zero zero bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1 bl1_n bl2 bl2_n bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar12Array_16X8BC
Xzero vdd vss zero zero_x1
.ends DP8TVar12TestArray_16X8

.subckt DP8TVar12Array_4X8 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar12Array_4X4
Xinst0x1 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar12Array_4X4
.ends DP8TVar12Array_4X8

.subckt DP8TVar12Array_2X4 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TVar12Array_2X2
Xinst0x1 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar12Array_2X2
.ends DP8TVar12Array_2X4

.subckt DP8TVar12Array_2X8 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar12Array_2X4
Xinst0x1 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar12Array_2X4
.ends DP8TVar12Array_2X8

.subckt DP8TVar12Array_1X2 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1]
Xinst0x0 wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] vdd vss DP8TVar12Cell
Xinst0x1 wl1[0] wl2[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] vdd vss DP8TVar12Cell
.ends DP8TVar12Array_1X2

.subckt DP8TVar12Array_1X4 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3]
Xinst0x0 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TVar12Array_1X2
Xinst0x1 vss vdd wl1[0] wl2[0] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar12Array_1X2
.ends DP8TVar12Array_1X4

.subckt DP8TVar12Array_1X8 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar12Array_1X4
Xinst0x1 vss vdd wl1[0] wl2[0] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar12Array_1X4
.ends DP8TVar12Array_1X8

.subckt DP8TVar12Array_7X8 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar12Array_4X8
Xinst1x0 vss vdd wl1[4] wl2[4] wl1[5] wl2[5] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar12Array_2X8
Xinst2x0 vss vdd wl1[6] wl2[6] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar12Array_1X8
.ends DP8TVar12Array_7X8

.subckt DP8TVar12CellShWL1 wl1 wl2 bl1 bl1_n bl2 bl2_n vdd vss
Xpu1 vdd bit_n bit vdd sg13_lv_pmos l=1.3e-07 w=2e-07
Xpd1 bit bit_n vss vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpu2 vdd bit bit_n vdd sg13_lv_pmos l=1.3e-07 w=2e-07
Xpd2 bit_n bit vss vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg1 bit wl1 bl1 vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg1n bit_n wl1 bl1_n vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg2 bit wl1 bl2 vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg2n bit_n wl1 bl2_n vss sg13_lv_nmos l=1.3e-07 w=2e-07
.ends DP8TVar12CellShWL1

.subckt DP8TVar12ArrayShWL1_1X2 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1]
Xinst0x0 wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] vdd vss DP8TVar12CellShWL1
Xinst0x1 wl1[0] wl2[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] vdd vss DP8TVar12CellShWL1
.ends DP8TVar12ArrayShWL1_1X2

.subckt DP8TVar12ArrayShWL1_1X4 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3]
Xinst0x0 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TVar12ArrayShWL1_1X2
Xinst0x1 vss vdd wl1[0] wl2[0] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar12ArrayShWL1_1X2
.ends DP8TVar12ArrayShWL1_1X4

.subckt DP8TVar12ArrayShWL1_1X8 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar12ArrayShWL1_1X4
Xinst0x1 vss vdd wl1[0] wl2[0] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar12ArrayShWL1_1X4
.ends DP8TVar12ArrayShWL1_1X8

.subckt DP8TVar12CellConnectOut wl1 wl2 bl1 bl1_n bl2 bl2_n vdd vss bit bit_n
Xpu1 vdd bit_n bit vdd sg13_lv_pmos l=1.3e-07 w=2e-07
Xpd1 bit bit_n vss vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpu2 vdd bit bit_n vdd sg13_lv_pmos l=1.3e-07 w=2e-07
Xpd2 bit_n bit vss vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg1 bit wl1 bl1 vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg1n bit_n wl1 bl1_n vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg2 bit wl2 bl2 vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg2n bit_n wl2 bl2_n vss sg13_lv_nmos l=1.3e-07 w=2e-07
.ends DP8TVar12CellConnectOut

.subckt DP8TVar12CellShWL2 wl1 wl2 bl1 bl1_n bl2 bl2_n vdd vss
Xpu1 vdd bit_n bit vdd sg13_lv_pmos l=1.3e-07 w=2e-07
Xpd1 bit bit_n vss vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpu2 vdd bit bit_n vdd sg13_lv_pmos l=1.3e-07 w=2e-07
Xpd2 bit_n bit vss vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg1 bit wl2 bl1 vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg1n bit_n wl2 bl1_n vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg2 bit wl2 bl2 vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg2n bit_n wl2 bl2_n vss sg13_lv_nmos l=1.3e-07 w=2e-07
.ends DP8TVar12CellShWL2

.subckt DP8TVar12ArrayShWL2_1X2 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1]
Xinst0x0 wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] vdd vss DP8TVar12CellShWL2
Xinst0x1 wl1[0] wl2[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] vdd vss DP8TVar12CellShWL2
.ends DP8TVar12ArrayShWL2_1X2

.subckt DP8TVar12ArrayShWL2_1X4 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3]
Xinst0x0 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TVar12ArrayShWL2_1X2
Xinst0x1 vss vdd wl1[0] wl2[0] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar12ArrayShWL2_1X2
.ends DP8TVar12ArrayShWL2_1X4

.subckt DP8TVar12ArrayShWL2_1X8 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar12ArrayShWL2_1X4
Xinst0x1 vss vdd wl1[0] wl2[0] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar12ArrayShWL2_1X4
.ends DP8TVar12ArrayShWL2_1X8

.subckt DP8TVar12Array_6X8 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar12Array_4X8
Xinst1x0 vss vdd wl1[4] wl2[4] wl1[5] wl2[5] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar12Array_2X8
.ends DP8TVar12Array_6X8

.subckt DP8TVar12TestArray_16X8C vss vdd wl1 wl2 bl1 bl1_n bl2 bl2_n bit bit_n
Xbcconn_bot vss vdd bcconn_bot_bl1[0] bcconn_bot_bl1_n[0] bcconn_bot_bl2[0] bcconn_bot_bl2_n[0] bcconn_bot_bl1[1] bcconn_bot_bl1_n[1] bcconn_bot_bl2[1] bcconn_bot_bl2_n[1] bcconn_bot_bl1[2] bcconn_bot_bl1_n[2] bcconn_bot_bl2[2] bcconn_bot_bl2_n[2] bcconn_bot_bl1[3] bcconn_bot_bl1_n[3] bcconn_bot_bl2[3] bcconn_bot_bl2_n[3] bl1 bl1_n bl2 bl2_n bcconn_bot_bl1[5] bcconn_bot_bl1_n[5] bcconn_bot_bl2[5] bcconn_bot_bl2_n[5] bcconn_bot_bl1[6] bcconn_bot_bl1_n[6] bcconn_bot_bl2[6] bcconn_bot_bl2_n[6] bcconn_bot_bl1[7] bcconn_bot_bl1_n[7] bcconn_bot_bl2[7] bcconn_bot_bl2_n[7] DP8TVar12BulkConnRow_8
Xbcconn_top vss vdd bcconn_top_bl1[0] bcconn_top_bl1_n[0] bcconn_top_bl2[0] bcconn_top_bl2_n[0] bcconn_top_bl1[1] bcconn_top_bl1_n[1] bcconn_top_bl2[1] bcconn_top_bl2_n[1] bcconn_top_bl1[2] bcconn_top_bl1_n[2] bcconn_top_bl2[2] bcconn_top_bl2_n[2] bcconn_top_bl1[3] bcconn_top_bl1_n[3] bcconn_top_bl2[3] bcconn_top_bl2_n[3] bl1 bl1_n bl2 bl2_n bcconn_top_bl1[5] bcconn_top_bl1_n[5] bcconn_top_bl2[5] bcconn_top_bl2_n[5] bcconn_top_bl1[6] bcconn_top_bl1_n[6] bcconn_top_bl2[6] bcconn_top_bl2_n[6] bcconn_top_bl1[7] bcconn_top_bl1_n[7] bcconn_top_bl2[7] bcconn_top_bl2_n[7] DP8TVar12BulkConnRow_8
Xarray_bot vss vdd zero zero zero zero zero zero zero zero zero zero zero zero zero zero array_bot_bl1[0] array_bot_bl1_n[0] array_bot_bl2[0] array_bot_bl2_n[0] array_bot_bl1[1] array_bot_bl1_n[1] array_bot_bl2[1] array_bot_bl2_n[1] array_bot_bl1[2] array_bot_bl1_n[2] array_bot_bl2[2] array_bot_bl2_n[2] array_bot_bl1[3] array_bot_bl1_n[3] array_bot_bl2[3] array_bot_bl2_n[3] bl1 bl1_n bl2 bl2_n array_bot_bl1[5] array_bot_bl1_n[5] array_bot_bl2[5] array_bot_bl2_n[5] array_bot_bl1[6] array_bot_bl1_n[6] array_bot_bl2[6] array_bot_bl2_n[6] array_bot_bl1[7] array_bot_bl1_n[7] array_bot_bl2[7] array_bot_bl2_n[7] DP8TVar12Array_7X8
Xshwl1_row vss vdd zero bit shwl1_row_bl1[0] shwl1_row_bl1_n[0] shwl1_row_bl2[0] shwl1_row_bl2_n[0] shwl1_row_bl1[1] shwl1_row_bl1_n[1] shwl1_row_bl2[1] shwl1_row_bl2_n[1] shwl1_row_bl1[2] shwl1_row_bl1_n[2] shwl1_row_bl2[2] shwl1_row_bl2_n[2] shwl1_row_bl1[3] shwl1_row_bl1_n[3] shwl1_row_bl2[3] shwl1_row_bl2_n[3] bl1 bl1_n bl2 bl2_n shwl1_row_bl1[5] shwl1_row_bl1_n[5] shwl1_row_bl2[5] shwl1_row_bl2_n[5] shwl1_row_bl1[6] shwl1_row_bl1_n[6] shwl1_row_bl2[6] shwl1_row_bl2_n[6] shwl1_row_bl1[7] shwl1_row_bl1_n[7] shwl1_row_bl2[7] shwl1_row_bl2_n[7] DP8TVar12ArrayShWL1_1X8
Xcell_cols_left vss vdd wl1 wl2 cell_cols_left_bl1[0] cell_cols_left_bl1_n[0] cell_cols_left_bl2[0] cell_cols_left_bl2_n[0] cell_cols_left_bl1[1] cell_cols_left_bl1_n[1] cell_cols_left_bl2[1] cell_cols_left_bl2_n[1] cell_cols_left_bl1[2] cell_cols_left_bl1_n[2] cell_cols_left_bl2[2] cell_cols_left_bl2_n[2] cell_cols_left_bl1[3] cell_cols_left_bl1_n[3] cell_cols_left_bl2[3] cell_cols_left_bl2_n[3] DP8TVar12Array_1X4
Xconncell wl1 wl2 bl1 bl1_n bl2 bl2_n vdd vss bit bit_n DP8TVar12CellConnectOut
Xfillcell wl1 wl2 fillcell_bl1 fillcell_bl1_n fillcell_bl2 fillcell_bl2_n vdd vss DP8TVar12Cell
Xcell_cols_right vss vdd wl1 wl2 cell_cols_right_bl1[0] cell_cols_right_bl1_n[0] cell_cols_right_bl2[0] cell_cols_right_bl2_n[0] cell_cols_right_bl1[1] cell_cols_right_bl1_n[1] cell_cols_right_bl2[1] cell_cols_right_bl2_n[1] DP8TVar12Array_1X2
Xshwl2_row vss vdd bit_n zero shwl2_row_bl1[0] shwl2_row_bl1_n[0] shwl2_row_bl2[0] shwl2_row_bl2_n[0] shwl2_row_bl1[1] shwl2_row_bl1_n[1] shwl2_row_bl2[1] shwl2_row_bl2_n[1] shwl2_row_bl1[2] shwl2_row_bl1_n[2] shwl2_row_bl2[2] shwl2_row_bl2_n[2] shwl2_row_bl1[3] shwl2_row_bl1_n[3] shwl2_row_bl2[3] shwl2_row_bl2_n[3] bl1 bl1_n bl2 bl2_n shwl2_row_bl1[5] shwl2_row_bl1_n[5] shwl2_row_bl2[5] shwl2_row_bl2_n[5] shwl2_row_bl1[6] shwl2_row_bl1_n[6] shwl2_row_bl2[6] shwl2_row_bl2_n[6] shwl2_row_bl1[7] shwl2_row_bl1_n[7] shwl2_row_bl2[7] shwl2_row_bl2_n[7] DP8TVar12ArrayShWL2_1X8
Xarray_top vss vdd zero zero zero zero zero zero zero zero zero zero zero zero array_top_bl1[0] array_top_bl1_n[0] array_top_bl2[0] array_top_bl2_n[0] array_top_bl1[1] array_top_bl1_n[1] array_top_bl2[1] array_top_bl2_n[1] array_top_bl1[2] array_top_bl1_n[2] array_top_bl2[2] array_top_bl2_n[2] array_top_bl1[3] array_top_bl1_n[3] array_top_bl2[3] array_top_bl2_n[3] bl1 bl1_n bl2 bl2_n array_top_bl1[5] array_top_bl1_n[5] array_top_bl2[5] array_top_bl2_n[5] array_top_bl1[6] array_top_bl1_n[6] array_top_bl2[6] array_top_bl2_n[6] array_top_bl1[7] array_top_bl1_n[7] array_top_bl2[7] array_top_bl2_n[7] DP8TVar12Array_6X8
Xzero vdd vss zero zero_x1
.ends DP8TVar12TestArray_16X8C

.subckt DP8TVar12 vss noco_vdd noco_wl1 noco_wl2 noco_bl1 noco_bl1_n noco_bl2 noco_bl2_n co_vdd co_bit co_bit_n co_wl1 co_wl2 co_bl1 co_bl1_n co_bl2_n co_bl2
Xframe noco_vdd noco_wl1 noco_wl2 noco_bl2 co_vdd co_bit co_bit_n co_wl1 co_wl2 NoConn_PAD0x9 vss noco_bl1 noco_bl1_n noco_bl2_n vss co_bl1 co_bl1_n co_bl2_n co_bl2 NoConn_PAD1x9 PadFrame_DP12
Xtestarray_noco vss noco_vdd noco_wl1 noco_wl2 noco_bl1 noco_bl1_n noco_bl2 noco_bl2_n DP8TVar12TestArray_16X8
Xtestarray_co vss co_vdd co_wl1 co_wl2 co_bl1 co_bl1_n co_bl2 co_bl2_n co_bit co_bit_n DP8TVar12TestArray_16X8C
.ends DP8TVar12

.subckt PadFrame_DP13 PAD0x0 PAD0x1 PAD0x2 PAD0x3 PAD0x4 PAD0x5 PAD0x6 PAD0x7 PAD0x8 PAD0x9 PAD1x0 PAD1x1 PAD1x2 PAD1x3 PAD1x4 PAD1x5 PAD1x6 PAD1x7 PAD1x8 PAD1x9
XPAD0x0 PAD0x0 BondPad
XPAD0x1 PAD0x1 BondPad
XPAD0x2 PAD0x2 BondPad
XPAD0x3 PAD0x3 BondPad
XPAD0x4 PAD0x4 BondPad
XPAD0x5 PAD0x5 BondPad
XPAD0x6 PAD0x6 BondPad
XPAD0x7 PAD0x7 BondPad
XPAD0x8 PAD0x8 BondPad
XPAD0x9 PAD0x9 BondPad
XPAD1x0 PAD1x0 BondPad
XPAD1x1 PAD1x1 BondPad
XPAD1x2 PAD1x2 BondPad
XPAD1x3 PAD1x3 BondPad
XPAD1x4 PAD1x4 BondPad
XPAD1x5 PAD1x5 BondPad
XPAD1x6 PAD1x6 BondPad
XPAD1x7 PAD1x7 BondPad
XPAD1x8 PAD1x8 BondPad
XPAD1x9 PAD1x9 BondPad
.ends PadFrame_DP13

.subckt DP8TVar13Cell wl1 wl2 bl1 bl1_n bl2 bl2_n vdd vss
Xpu1 vdd bit_n bit vdd sg13_lv_pmos l=1.3e-07 w=1.5e-07
Xpd1 bit bit_n vss vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpu2 vdd bit bit_n vdd sg13_lv_pmos l=1.3e-07 w=1.5e-07
Xpd2 bit_n bit vss vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg1 bit wl1 bl1 vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg1n bit_n wl1 bl1_n vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg2 bit wl2 bl2 vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg2n bit_n wl2 bl2_n vss sg13_lv_nmos l=1.3e-07 w=2e-07
.ends DP8TVar13Cell

.subckt DP8TVar13Array_2X1 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0]
Xinst0x0 wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] vdd vss DP8TVar13Cell
Xinst1x0 wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0] vdd vss DP8TVar13Cell
.ends DP8TVar13Array_2X1

.subckt DP8TVar13Array_2X2 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0] DP8TVar13Array_2X1
Xinst0x1 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TVar13Array_2X1
.ends DP8TVar13Array_2X2

.subckt DP8TVar13Array_4X2 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TVar13Array_2X2
Xinst1x0 vss vdd wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TVar13Array_2X2
.ends DP8TVar13Array_4X2

.subckt DP8TVar13Array_4X4 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TVar13Array_4X2
Xinst0x1 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar13Array_4X2
.ends DP8TVar13Array_4X4

.subckt DP8TVar13Array_8X4 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar13Array_4X4
Xinst1x0 vss vdd wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar13Array_4X4
.ends DP8TVar13Array_8X4

.subckt DP8TVar13Array_8X8 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar13Array_8X4
Xinst0x1 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar13Array_8X4
.ends DP8TVar13Array_8X8

.subckt DP8TVar13BulkConn vdd vss bl1 bl2 bl1_n bl2_n
.ends DP8TVar13BulkConn

.subckt DP8TVar13BulkConnRow_2 vss vdd bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1]
Xinst0 vdd vss bl1[0] bl2[0] bl1_n[0] bl2_n[0] DP8TVar13BulkConn
Xinst1 vdd vss bl1[1] bl2[1] bl1_n[1] bl2_n[1] DP8TVar13BulkConn
.ends DP8TVar13BulkConnRow_2

.subckt DP8TVar13BulkConnRow_4 vss vdd bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3]
Xinst0 vss vdd bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TVar13BulkConnRow_2
Xinst1 vss vdd bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar13BulkConnRow_2
.ends DP8TVar13BulkConnRow_4

.subckt DP8TVar13BulkConnRow_8 vss vdd bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0 vss vdd bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar13BulkConnRow_4
Xinst1 vss vdd bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar13BulkConnRow_4
.ends DP8TVar13BulkConnRow_8

.subckt DP8TVar13Array_16X8BC vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] wl1[8] wl2[8] wl1[9] wl2[9] wl1[10] wl2[10] wl1[11] wl2[11] wl1[12] wl2[12] wl1[13] wl2[13] wl1[14] wl2[14] wl1[15] wl2[15] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar13Array_8X8
Xinst1x0 vss vdd wl1[8] wl2[8] wl1[9] wl2[9] wl1[10] wl2[10] wl1[11] wl2[11] wl1[12] wl2[12] wl1[13] wl2[13] wl1[14] wl2[14] wl1[15] wl2[15] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar13Array_8X8
Xbottombcrow vss vdd bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar13BulkConnRow_8
Xtopbcrow vss vdd bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar13BulkConnRow_8
.ends DP8TVar13Array_16X8BC

.subckt DP8TVar13TestArray_16X8 vss vdd wl1 wl2 bl1 bl1_n bl2 bl2_n
Xarray vss vdd zero zero zero zero zero zero zero zero zero zero zero zero zero zero zero zero wl1 wl2 zero zero zero zero zero zero zero zero zero zero zero zero zero zero bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1 bl1_n bl2 bl2_n bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar13Array_16X8BC
Xzero vdd vss zero zero_x1
.ends DP8TVar13TestArray_16X8

.subckt DP8TVar13Array_4X8 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar13Array_4X4
Xinst0x1 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar13Array_4X4
.ends DP8TVar13Array_4X8

.subckt DP8TVar13Array_2X4 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TVar13Array_2X2
Xinst0x1 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar13Array_2X2
.ends DP8TVar13Array_2X4

.subckt DP8TVar13Array_2X8 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar13Array_2X4
Xinst0x1 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar13Array_2X4
.ends DP8TVar13Array_2X8

.subckt DP8TVar13Array_1X2 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1]
Xinst0x0 wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] vdd vss DP8TVar13Cell
Xinst0x1 wl1[0] wl2[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] vdd vss DP8TVar13Cell
.ends DP8TVar13Array_1X2

.subckt DP8TVar13Array_1X4 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3]
Xinst0x0 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TVar13Array_1X2
Xinst0x1 vss vdd wl1[0] wl2[0] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar13Array_1X2
.ends DP8TVar13Array_1X4

.subckt DP8TVar13Array_1X8 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar13Array_1X4
Xinst0x1 vss vdd wl1[0] wl2[0] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar13Array_1X4
.ends DP8TVar13Array_1X8

.subckt DP8TVar13Array_7X8 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar13Array_4X8
Xinst1x0 vss vdd wl1[4] wl2[4] wl1[5] wl2[5] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar13Array_2X8
Xinst2x0 vss vdd wl1[6] wl2[6] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar13Array_1X8
.ends DP8TVar13Array_7X8

.subckt DP8TVar13CellShWL1 wl1 wl2 bl1 bl1_n bl2 bl2_n vdd vss
Xpu1 vdd bit_n bit vdd sg13_lv_pmos l=1.3e-07 w=1.5e-07
Xpd1 bit bit_n vss vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpu2 vdd bit bit_n vdd sg13_lv_pmos l=1.3e-07 w=1.5e-07
Xpd2 bit_n bit vss vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg1 bit wl1 bl1 vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg1n bit_n wl1 bl1_n vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg2 bit wl1 bl2 vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg2n bit_n wl1 bl2_n vss sg13_lv_nmos l=1.3e-07 w=2e-07
.ends DP8TVar13CellShWL1

.subckt DP8TVar13ArrayShWL1_1X2 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1]
Xinst0x0 wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] vdd vss DP8TVar13CellShWL1
Xinst0x1 wl1[0] wl2[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] vdd vss DP8TVar13CellShWL1
.ends DP8TVar13ArrayShWL1_1X2

.subckt DP8TVar13ArrayShWL1_1X4 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3]
Xinst0x0 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TVar13ArrayShWL1_1X2
Xinst0x1 vss vdd wl1[0] wl2[0] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar13ArrayShWL1_1X2
.ends DP8TVar13ArrayShWL1_1X4

.subckt DP8TVar13ArrayShWL1_1X8 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar13ArrayShWL1_1X4
Xinst0x1 vss vdd wl1[0] wl2[0] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar13ArrayShWL1_1X4
.ends DP8TVar13ArrayShWL1_1X8

.subckt DP8TVar13CellConnectOut wl1 wl2 bl1 bl1_n bl2 bl2_n vdd vss bit bit_n
Xpu1 vdd bit_n bit vdd sg13_lv_pmos l=1.3e-07 w=1.5e-07
Xpd1 bit bit_n vss vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpu2 vdd bit bit_n vdd sg13_lv_pmos l=1.3e-07 w=1.5e-07
Xpd2 bit_n bit vss vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg1 bit wl1 bl1 vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg1n bit_n wl1 bl1_n vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg2 bit wl2 bl2 vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg2n bit_n wl2 bl2_n vss sg13_lv_nmos l=1.3e-07 w=2e-07
.ends DP8TVar13CellConnectOut

.subckt DP8TVar13CellShWL2 wl1 wl2 bl1 bl1_n bl2 bl2_n vdd vss
Xpu1 vdd bit_n bit vdd sg13_lv_pmos l=1.3e-07 w=1.5e-07
Xpd1 bit bit_n vss vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpu2 vdd bit bit_n vdd sg13_lv_pmos l=1.3e-07 w=1.5e-07
Xpd2 bit_n bit vss vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg1 bit wl2 bl1 vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg1n bit_n wl2 bl1_n vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg2 bit wl2 bl2 vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg2n bit_n wl2 bl2_n vss sg13_lv_nmos l=1.3e-07 w=2e-07
.ends DP8TVar13CellShWL2

.subckt DP8TVar13ArrayShWL2_1X2 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1]
Xinst0x0 wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] vdd vss DP8TVar13CellShWL2
Xinst0x1 wl1[0] wl2[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] vdd vss DP8TVar13CellShWL2
.ends DP8TVar13ArrayShWL2_1X2

.subckt DP8TVar13ArrayShWL2_1X4 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3]
Xinst0x0 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TVar13ArrayShWL2_1X2
Xinst0x1 vss vdd wl1[0] wl2[0] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar13ArrayShWL2_1X2
.ends DP8TVar13ArrayShWL2_1X4

.subckt DP8TVar13ArrayShWL2_1X8 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar13ArrayShWL2_1X4
Xinst0x1 vss vdd wl1[0] wl2[0] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar13ArrayShWL2_1X4
.ends DP8TVar13ArrayShWL2_1X8

.subckt DP8TVar13Array_6X8 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar13Array_4X8
Xinst1x0 vss vdd wl1[4] wl2[4] wl1[5] wl2[5] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar13Array_2X8
.ends DP8TVar13Array_6X8

.subckt DP8TVar13TestArray_16X8C vss vdd wl1 wl2 bl1 bl1_n bl2 bl2_n bit bit_n
Xbcconn_bot vss vdd bcconn_bot_bl1[0] bcconn_bot_bl1_n[0] bcconn_bot_bl2[0] bcconn_bot_bl2_n[0] bcconn_bot_bl1[1] bcconn_bot_bl1_n[1] bcconn_bot_bl2[1] bcconn_bot_bl2_n[1] bcconn_bot_bl1[2] bcconn_bot_bl1_n[2] bcconn_bot_bl2[2] bcconn_bot_bl2_n[2] bcconn_bot_bl1[3] bcconn_bot_bl1_n[3] bcconn_bot_bl2[3] bcconn_bot_bl2_n[3] bl1 bl1_n bl2 bl2_n bcconn_bot_bl1[5] bcconn_bot_bl1_n[5] bcconn_bot_bl2[5] bcconn_bot_bl2_n[5] bcconn_bot_bl1[6] bcconn_bot_bl1_n[6] bcconn_bot_bl2[6] bcconn_bot_bl2_n[6] bcconn_bot_bl1[7] bcconn_bot_bl1_n[7] bcconn_bot_bl2[7] bcconn_bot_bl2_n[7] DP8TVar13BulkConnRow_8
Xbcconn_top vss vdd bcconn_top_bl1[0] bcconn_top_bl1_n[0] bcconn_top_bl2[0] bcconn_top_bl2_n[0] bcconn_top_bl1[1] bcconn_top_bl1_n[1] bcconn_top_bl2[1] bcconn_top_bl2_n[1] bcconn_top_bl1[2] bcconn_top_bl1_n[2] bcconn_top_bl2[2] bcconn_top_bl2_n[2] bcconn_top_bl1[3] bcconn_top_bl1_n[3] bcconn_top_bl2[3] bcconn_top_bl2_n[3] bl1 bl1_n bl2 bl2_n bcconn_top_bl1[5] bcconn_top_bl1_n[5] bcconn_top_bl2[5] bcconn_top_bl2_n[5] bcconn_top_bl1[6] bcconn_top_bl1_n[6] bcconn_top_bl2[6] bcconn_top_bl2_n[6] bcconn_top_bl1[7] bcconn_top_bl1_n[7] bcconn_top_bl2[7] bcconn_top_bl2_n[7] DP8TVar13BulkConnRow_8
Xarray_bot vss vdd zero zero zero zero zero zero zero zero zero zero zero zero zero zero array_bot_bl1[0] array_bot_bl1_n[0] array_bot_bl2[0] array_bot_bl2_n[0] array_bot_bl1[1] array_bot_bl1_n[1] array_bot_bl2[1] array_bot_bl2_n[1] array_bot_bl1[2] array_bot_bl1_n[2] array_bot_bl2[2] array_bot_bl2_n[2] array_bot_bl1[3] array_bot_bl1_n[3] array_bot_bl2[3] array_bot_bl2_n[3] bl1 bl1_n bl2 bl2_n array_bot_bl1[5] array_bot_bl1_n[5] array_bot_bl2[5] array_bot_bl2_n[5] array_bot_bl1[6] array_bot_bl1_n[6] array_bot_bl2[6] array_bot_bl2_n[6] array_bot_bl1[7] array_bot_bl1_n[7] array_bot_bl2[7] array_bot_bl2_n[7] DP8TVar13Array_7X8
Xshwl1_row vss vdd zero bit shwl1_row_bl1[0] shwl1_row_bl1_n[0] shwl1_row_bl2[0] shwl1_row_bl2_n[0] shwl1_row_bl1[1] shwl1_row_bl1_n[1] shwl1_row_bl2[1] shwl1_row_bl2_n[1] shwl1_row_bl1[2] shwl1_row_bl1_n[2] shwl1_row_bl2[2] shwl1_row_bl2_n[2] shwl1_row_bl1[3] shwl1_row_bl1_n[3] shwl1_row_bl2[3] shwl1_row_bl2_n[3] bl1 bl1_n bl2 bl2_n shwl1_row_bl1[5] shwl1_row_bl1_n[5] shwl1_row_bl2[5] shwl1_row_bl2_n[5] shwl1_row_bl1[6] shwl1_row_bl1_n[6] shwl1_row_bl2[6] shwl1_row_bl2_n[6] shwl1_row_bl1[7] shwl1_row_bl1_n[7] shwl1_row_bl2[7] shwl1_row_bl2_n[7] DP8TVar13ArrayShWL1_1X8
Xcell_cols_left vss vdd wl1 wl2 cell_cols_left_bl1[0] cell_cols_left_bl1_n[0] cell_cols_left_bl2[0] cell_cols_left_bl2_n[0] cell_cols_left_bl1[1] cell_cols_left_bl1_n[1] cell_cols_left_bl2[1] cell_cols_left_bl2_n[1] cell_cols_left_bl1[2] cell_cols_left_bl1_n[2] cell_cols_left_bl2[2] cell_cols_left_bl2_n[2] cell_cols_left_bl1[3] cell_cols_left_bl1_n[3] cell_cols_left_bl2[3] cell_cols_left_bl2_n[3] DP8TVar13Array_1X4
Xconncell wl1 wl2 bl1 bl1_n bl2 bl2_n vdd vss bit bit_n DP8TVar13CellConnectOut
Xfillcell wl1 wl2 fillcell_bl1 fillcell_bl1_n fillcell_bl2 fillcell_bl2_n vdd vss DP8TVar13Cell
Xcell_cols_right vss vdd wl1 wl2 cell_cols_right_bl1[0] cell_cols_right_bl1_n[0] cell_cols_right_bl2[0] cell_cols_right_bl2_n[0] cell_cols_right_bl1[1] cell_cols_right_bl1_n[1] cell_cols_right_bl2[1] cell_cols_right_bl2_n[1] DP8TVar13Array_1X2
Xshwl2_row vss vdd bit_n zero shwl2_row_bl1[0] shwl2_row_bl1_n[0] shwl2_row_bl2[0] shwl2_row_bl2_n[0] shwl2_row_bl1[1] shwl2_row_bl1_n[1] shwl2_row_bl2[1] shwl2_row_bl2_n[1] shwl2_row_bl1[2] shwl2_row_bl1_n[2] shwl2_row_bl2[2] shwl2_row_bl2_n[2] shwl2_row_bl1[3] shwl2_row_bl1_n[3] shwl2_row_bl2[3] shwl2_row_bl2_n[3] bl1 bl1_n bl2 bl2_n shwl2_row_bl1[5] shwl2_row_bl1_n[5] shwl2_row_bl2[5] shwl2_row_bl2_n[5] shwl2_row_bl1[6] shwl2_row_bl1_n[6] shwl2_row_bl2[6] shwl2_row_bl2_n[6] shwl2_row_bl1[7] shwl2_row_bl1_n[7] shwl2_row_bl2[7] shwl2_row_bl2_n[7] DP8TVar13ArrayShWL2_1X8
Xarray_top vss vdd zero zero zero zero zero zero zero zero zero zero zero zero array_top_bl1[0] array_top_bl1_n[0] array_top_bl2[0] array_top_bl2_n[0] array_top_bl1[1] array_top_bl1_n[1] array_top_bl2[1] array_top_bl2_n[1] array_top_bl1[2] array_top_bl1_n[2] array_top_bl2[2] array_top_bl2_n[2] array_top_bl1[3] array_top_bl1_n[3] array_top_bl2[3] array_top_bl2_n[3] bl1 bl1_n bl2 bl2_n array_top_bl1[5] array_top_bl1_n[5] array_top_bl2[5] array_top_bl2_n[5] array_top_bl1[6] array_top_bl1_n[6] array_top_bl2[6] array_top_bl2_n[6] array_top_bl1[7] array_top_bl1_n[7] array_top_bl2[7] array_top_bl2_n[7] DP8TVar13Array_6X8
Xzero vdd vss zero zero_x1
.ends DP8TVar13TestArray_16X8C

.subckt DP8TVar13 vss noco_vdd noco_wl1 noco_wl2 noco_bl1 noco_bl1_n noco_bl2 noco_bl2_n co_vdd co_bit co_bit_n co_wl1 co_wl2 co_bl1 co_bl1_n co_bl2_n co_bl2
Xframe noco_vdd noco_wl1 noco_wl2 noco_bl2 co_vdd co_bit co_bit_n co_wl1 co_wl2 NoConn_PAD0x9 vss noco_bl1 noco_bl1_n noco_bl2_n vss co_bl1 co_bl1_n co_bl2_n co_bl2 NoConn_PAD1x9 PadFrame_DP13
Xtestarray_noco vss noco_vdd noco_wl1 noco_wl2 noco_bl1 noco_bl1_n noco_bl2 noco_bl2_n DP8TVar13TestArray_16X8
Xtestarray_co vss co_vdd co_wl1 co_wl2 co_bl1 co_bl1_n co_bl2 co_bl2_n co_bit co_bit_n DP8TVar13TestArray_16X8C
.ends DP8TVar13

.subckt PadFrame_DP14 PAD0x0 PAD0x1 PAD0x2 PAD0x3 PAD0x4 PAD0x5 PAD0x6 PAD0x7 PAD0x8 PAD0x9 PAD1x0 PAD1x1 PAD1x2 PAD1x3 PAD1x4 PAD1x5 PAD1x6 PAD1x7 PAD1x8 PAD1x9
XPAD0x0 PAD0x0 BondPad
XPAD0x1 PAD0x1 BondPad
XPAD0x2 PAD0x2 BondPad
XPAD0x3 PAD0x3 BondPad
XPAD0x4 PAD0x4 BondPad
XPAD0x5 PAD0x5 BondPad
XPAD0x6 PAD0x6 BondPad
XPAD0x7 PAD0x7 BondPad
XPAD0x8 PAD0x8 BondPad
XPAD0x9 PAD0x9 BondPad
XPAD1x0 PAD1x0 BondPad
XPAD1x1 PAD1x1 BondPad
XPAD1x2 PAD1x2 BondPad
XPAD1x3 PAD1x3 BondPad
XPAD1x4 PAD1x4 BondPad
XPAD1x5 PAD1x5 BondPad
XPAD1x6 PAD1x6 BondPad
XPAD1x7 PAD1x7 BondPad
XPAD1x8 PAD1x8 BondPad
XPAD1x9 PAD1x9 BondPad
.ends PadFrame_DP14

.subckt DP8TVar14Cell wl1 wl2 bl1 bl1_n bl2 bl2_n vdd vss
Xpu1 vdd bit_n bit vdd sg13_lv_pmos l=1.3e-07 w=3e-07
Xpd1 bit bit_n vss vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpu2 vdd bit bit_n vdd sg13_lv_pmos l=1.3e-07 w=3e-07
Xpd2 bit_n bit vss vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg1 bit wl1 bl1 vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg1n bit_n wl1 bl1_n vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg2 bit wl2 bl2 vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg2n bit_n wl2 bl2_n vss sg13_lv_nmos l=1.3e-07 w=3e-07
.ends DP8TVar14Cell

.subckt DP8TVar14Array_2X1 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0]
Xinst0x0 wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] vdd vss DP8TVar14Cell
Xinst1x0 wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0] vdd vss DP8TVar14Cell
.ends DP8TVar14Array_2X1

.subckt DP8TVar14Array_2X2 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0] DP8TVar14Array_2X1
Xinst0x1 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TVar14Array_2X1
.ends DP8TVar14Array_2X2

.subckt DP8TVar14Array_4X2 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TVar14Array_2X2
Xinst1x0 vss vdd wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TVar14Array_2X2
.ends DP8TVar14Array_4X2

.subckt DP8TVar14Array_4X4 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TVar14Array_4X2
Xinst0x1 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar14Array_4X2
.ends DP8TVar14Array_4X4

.subckt DP8TVar14Array_8X4 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar14Array_4X4
Xinst1x0 vss vdd wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar14Array_4X4
.ends DP8TVar14Array_8X4

.subckt DP8TVar14Array_8X8 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar14Array_8X4
Xinst0x1 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar14Array_8X4
.ends DP8TVar14Array_8X8

.subckt DP8TVar14BulkConn vdd vss bl1 bl2 bl1_n bl2_n
.ends DP8TVar14BulkConn

.subckt DP8TVar14BulkConnRow_2 vss vdd bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1]
Xinst0 vdd vss bl1[0] bl2[0] bl1_n[0] bl2_n[0] DP8TVar14BulkConn
Xinst1 vdd vss bl1[1] bl2[1] bl1_n[1] bl2_n[1] DP8TVar14BulkConn
.ends DP8TVar14BulkConnRow_2

.subckt DP8TVar14BulkConnRow_4 vss vdd bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3]
Xinst0 vss vdd bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TVar14BulkConnRow_2
Xinst1 vss vdd bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar14BulkConnRow_2
.ends DP8TVar14BulkConnRow_4

.subckt DP8TVar14BulkConnRow_8 vss vdd bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0 vss vdd bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar14BulkConnRow_4
Xinst1 vss vdd bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar14BulkConnRow_4
.ends DP8TVar14BulkConnRow_8

.subckt DP8TVar14Array_16X8BC vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] wl1[8] wl2[8] wl1[9] wl2[9] wl1[10] wl2[10] wl1[11] wl2[11] wl1[12] wl2[12] wl1[13] wl2[13] wl1[14] wl2[14] wl1[15] wl2[15] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar14Array_8X8
Xinst1x0 vss vdd wl1[8] wl2[8] wl1[9] wl2[9] wl1[10] wl2[10] wl1[11] wl2[11] wl1[12] wl2[12] wl1[13] wl2[13] wl1[14] wl2[14] wl1[15] wl2[15] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar14Array_8X8
Xbottombcrow vss vdd bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar14BulkConnRow_8
Xtopbcrow vss vdd bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar14BulkConnRow_8
.ends DP8TVar14Array_16X8BC

.subckt DP8TVar14TestArray_16X8 vss vdd wl1 wl2 bl1 bl1_n bl2 bl2_n
Xarray vss vdd zero zero zero zero zero zero zero zero zero zero zero zero zero zero zero zero wl1 wl2 zero zero zero zero zero zero zero zero zero zero zero zero zero zero bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1 bl1_n bl2 bl2_n bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar14Array_16X8BC
Xzero vdd vss zero zero_x1
.ends DP8TVar14TestArray_16X8

.subckt DP8TVar14Array_4X8 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar14Array_4X4
Xinst0x1 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar14Array_4X4
.ends DP8TVar14Array_4X8

.subckt DP8TVar14Array_2X4 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TVar14Array_2X2
Xinst0x1 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar14Array_2X2
.ends DP8TVar14Array_2X4

.subckt DP8TVar14Array_2X8 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar14Array_2X4
Xinst0x1 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar14Array_2X4
.ends DP8TVar14Array_2X8

.subckt DP8TVar14Array_1X2 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1]
Xinst0x0 wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] vdd vss DP8TVar14Cell
Xinst0x1 wl1[0] wl2[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] vdd vss DP8TVar14Cell
.ends DP8TVar14Array_1X2

.subckt DP8TVar14Array_1X4 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3]
Xinst0x0 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TVar14Array_1X2
Xinst0x1 vss vdd wl1[0] wl2[0] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar14Array_1X2
.ends DP8TVar14Array_1X4

.subckt DP8TVar14Array_1X8 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar14Array_1X4
Xinst0x1 vss vdd wl1[0] wl2[0] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar14Array_1X4
.ends DP8TVar14Array_1X8

.subckt DP8TVar14Array_7X8 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar14Array_4X8
Xinst1x0 vss vdd wl1[4] wl2[4] wl1[5] wl2[5] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar14Array_2X8
Xinst2x0 vss vdd wl1[6] wl2[6] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar14Array_1X8
.ends DP8TVar14Array_7X8

.subckt DP8TVar14CellShWL1 wl1 wl2 bl1 bl1_n bl2 bl2_n vdd vss
Xpu1 vdd bit_n bit vdd sg13_lv_pmos l=1.3e-07 w=3e-07
Xpd1 bit bit_n vss vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpu2 vdd bit bit_n vdd sg13_lv_pmos l=1.3e-07 w=3e-07
Xpd2 bit_n bit vss vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg1 bit wl1 bl1 vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg1n bit_n wl1 bl1_n vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg2 bit wl1 bl2 vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg2n bit_n wl1 bl2_n vss sg13_lv_nmos l=1.3e-07 w=3e-07
.ends DP8TVar14CellShWL1

.subckt DP8TVar14ArrayShWL1_1X2 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1]
Xinst0x0 wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] vdd vss DP8TVar14CellShWL1
Xinst0x1 wl1[0] wl2[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] vdd vss DP8TVar14CellShWL1
.ends DP8TVar14ArrayShWL1_1X2

.subckt DP8TVar14ArrayShWL1_1X4 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3]
Xinst0x0 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TVar14ArrayShWL1_1X2
Xinst0x1 vss vdd wl1[0] wl2[0] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar14ArrayShWL1_1X2
.ends DP8TVar14ArrayShWL1_1X4

.subckt DP8TVar14ArrayShWL1_1X8 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar14ArrayShWL1_1X4
Xinst0x1 vss vdd wl1[0] wl2[0] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar14ArrayShWL1_1X4
.ends DP8TVar14ArrayShWL1_1X8

.subckt DP8TVar14CellConnectOut wl1 wl2 bl1 bl1_n bl2 bl2_n vdd vss bit bit_n
Xpu1 vdd bit_n bit vdd sg13_lv_pmos l=1.3e-07 w=3e-07
Xpd1 bit bit_n vss vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpu2 vdd bit bit_n vdd sg13_lv_pmos l=1.3e-07 w=3e-07
Xpd2 bit_n bit vss vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg1 bit wl1 bl1 vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg1n bit_n wl1 bl1_n vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg2 bit wl2 bl2 vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg2n bit_n wl2 bl2_n vss sg13_lv_nmos l=1.3e-07 w=3e-07
.ends DP8TVar14CellConnectOut

.subckt DP8TVar14CellShWL2 wl1 wl2 bl1 bl1_n bl2 bl2_n vdd vss
Xpu1 vdd bit_n bit vdd sg13_lv_pmos l=1.3e-07 w=3e-07
Xpd1 bit bit_n vss vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpu2 vdd bit bit_n vdd sg13_lv_pmos l=1.3e-07 w=3e-07
Xpd2 bit_n bit vss vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg1 bit wl2 bl1 vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg1n bit_n wl2 bl1_n vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg2 bit wl2 bl2 vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg2n bit_n wl2 bl2_n vss sg13_lv_nmos l=1.3e-07 w=3e-07
.ends DP8TVar14CellShWL2

.subckt DP8TVar14ArrayShWL2_1X2 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1]
Xinst0x0 wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] vdd vss DP8TVar14CellShWL2
Xinst0x1 wl1[0] wl2[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] vdd vss DP8TVar14CellShWL2
.ends DP8TVar14ArrayShWL2_1X2

.subckt DP8TVar14ArrayShWL2_1X4 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3]
Xinst0x0 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TVar14ArrayShWL2_1X2
Xinst0x1 vss vdd wl1[0] wl2[0] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar14ArrayShWL2_1X2
.ends DP8TVar14ArrayShWL2_1X4

.subckt DP8TVar14ArrayShWL2_1X8 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar14ArrayShWL2_1X4
Xinst0x1 vss vdd wl1[0] wl2[0] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar14ArrayShWL2_1X4
.ends DP8TVar14ArrayShWL2_1X8

.subckt DP8TVar14Array_6X8 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar14Array_4X8
Xinst1x0 vss vdd wl1[4] wl2[4] wl1[5] wl2[5] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar14Array_2X8
.ends DP8TVar14Array_6X8

.subckt DP8TVar14TestArray_16X8C vss vdd wl1 wl2 bl1 bl1_n bl2 bl2_n bit bit_n
Xbcconn_bot vss vdd bcconn_bot_bl1[0] bcconn_bot_bl1_n[0] bcconn_bot_bl2[0] bcconn_bot_bl2_n[0] bcconn_bot_bl1[1] bcconn_bot_bl1_n[1] bcconn_bot_bl2[1] bcconn_bot_bl2_n[1] bcconn_bot_bl1[2] bcconn_bot_bl1_n[2] bcconn_bot_bl2[2] bcconn_bot_bl2_n[2] bcconn_bot_bl1[3] bcconn_bot_bl1_n[3] bcconn_bot_bl2[3] bcconn_bot_bl2_n[3] bl1 bl1_n bl2 bl2_n bcconn_bot_bl1[5] bcconn_bot_bl1_n[5] bcconn_bot_bl2[5] bcconn_bot_bl2_n[5] bcconn_bot_bl1[6] bcconn_bot_bl1_n[6] bcconn_bot_bl2[6] bcconn_bot_bl2_n[6] bcconn_bot_bl1[7] bcconn_bot_bl1_n[7] bcconn_bot_bl2[7] bcconn_bot_bl2_n[7] DP8TVar14BulkConnRow_8
Xbcconn_top vss vdd bcconn_top_bl1[0] bcconn_top_bl1_n[0] bcconn_top_bl2[0] bcconn_top_bl2_n[0] bcconn_top_bl1[1] bcconn_top_bl1_n[1] bcconn_top_bl2[1] bcconn_top_bl2_n[1] bcconn_top_bl1[2] bcconn_top_bl1_n[2] bcconn_top_bl2[2] bcconn_top_bl2_n[2] bcconn_top_bl1[3] bcconn_top_bl1_n[3] bcconn_top_bl2[3] bcconn_top_bl2_n[3] bl1 bl1_n bl2 bl2_n bcconn_top_bl1[5] bcconn_top_bl1_n[5] bcconn_top_bl2[5] bcconn_top_bl2_n[5] bcconn_top_bl1[6] bcconn_top_bl1_n[6] bcconn_top_bl2[6] bcconn_top_bl2_n[6] bcconn_top_bl1[7] bcconn_top_bl1_n[7] bcconn_top_bl2[7] bcconn_top_bl2_n[7] DP8TVar14BulkConnRow_8
Xarray_bot vss vdd zero zero zero zero zero zero zero zero zero zero zero zero zero zero array_bot_bl1[0] array_bot_bl1_n[0] array_bot_bl2[0] array_bot_bl2_n[0] array_bot_bl1[1] array_bot_bl1_n[1] array_bot_bl2[1] array_bot_bl2_n[1] array_bot_bl1[2] array_bot_bl1_n[2] array_bot_bl2[2] array_bot_bl2_n[2] array_bot_bl1[3] array_bot_bl1_n[3] array_bot_bl2[3] array_bot_bl2_n[3] bl1 bl1_n bl2 bl2_n array_bot_bl1[5] array_bot_bl1_n[5] array_bot_bl2[5] array_bot_bl2_n[5] array_bot_bl1[6] array_bot_bl1_n[6] array_bot_bl2[6] array_bot_bl2_n[6] array_bot_bl1[7] array_bot_bl1_n[7] array_bot_bl2[7] array_bot_bl2_n[7] DP8TVar14Array_7X8
Xshwl1_row vss vdd zero bit shwl1_row_bl1[0] shwl1_row_bl1_n[0] shwl1_row_bl2[0] shwl1_row_bl2_n[0] shwl1_row_bl1[1] shwl1_row_bl1_n[1] shwl1_row_bl2[1] shwl1_row_bl2_n[1] shwl1_row_bl1[2] shwl1_row_bl1_n[2] shwl1_row_bl2[2] shwl1_row_bl2_n[2] shwl1_row_bl1[3] shwl1_row_bl1_n[3] shwl1_row_bl2[3] shwl1_row_bl2_n[3] bl1 bl1_n bl2 bl2_n shwl1_row_bl1[5] shwl1_row_bl1_n[5] shwl1_row_bl2[5] shwl1_row_bl2_n[5] shwl1_row_bl1[6] shwl1_row_bl1_n[6] shwl1_row_bl2[6] shwl1_row_bl2_n[6] shwl1_row_bl1[7] shwl1_row_bl1_n[7] shwl1_row_bl2[7] shwl1_row_bl2_n[7] DP8TVar14ArrayShWL1_1X8
Xcell_cols_left vss vdd wl1 wl2 cell_cols_left_bl1[0] cell_cols_left_bl1_n[0] cell_cols_left_bl2[0] cell_cols_left_bl2_n[0] cell_cols_left_bl1[1] cell_cols_left_bl1_n[1] cell_cols_left_bl2[1] cell_cols_left_bl2_n[1] cell_cols_left_bl1[2] cell_cols_left_bl1_n[2] cell_cols_left_bl2[2] cell_cols_left_bl2_n[2] cell_cols_left_bl1[3] cell_cols_left_bl1_n[3] cell_cols_left_bl2[3] cell_cols_left_bl2_n[3] DP8TVar14Array_1X4
Xconncell wl1 wl2 bl1 bl1_n bl2 bl2_n vdd vss bit bit_n DP8TVar14CellConnectOut
Xfillcell wl1 wl2 fillcell_bl1 fillcell_bl1_n fillcell_bl2 fillcell_bl2_n vdd vss DP8TVar14Cell
Xcell_cols_right vss vdd wl1 wl2 cell_cols_right_bl1[0] cell_cols_right_bl1_n[0] cell_cols_right_bl2[0] cell_cols_right_bl2_n[0] cell_cols_right_bl1[1] cell_cols_right_bl1_n[1] cell_cols_right_bl2[1] cell_cols_right_bl2_n[1] DP8TVar14Array_1X2
Xshwl2_row vss vdd bit_n zero shwl2_row_bl1[0] shwl2_row_bl1_n[0] shwl2_row_bl2[0] shwl2_row_bl2_n[0] shwl2_row_bl1[1] shwl2_row_bl1_n[1] shwl2_row_bl2[1] shwl2_row_bl2_n[1] shwl2_row_bl1[2] shwl2_row_bl1_n[2] shwl2_row_bl2[2] shwl2_row_bl2_n[2] shwl2_row_bl1[3] shwl2_row_bl1_n[3] shwl2_row_bl2[3] shwl2_row_bl2_n[3] bl1 bl1_n bl2 bl2_n shwl2_row_bl1[5] shwl2_row_bl1_n[5] shwl2_row_bl2[5] shwl2_row_bl2_n[5] shwl2_row_bl1[6] shwl2_row_bl1_n[6] shwl2_row_bl2[6] shwl2_row_bl2_n[6] shwl2_row_bl1[7] shwl2_row_bl1_n[7] shwl2_row_bl2[7] shwl2_row_bl2_n[7] DP8TVar14ArrayShWL2_1X8
Xarray_top vss vdd zero zero zero zero zero zero zero zero zero zero zero zero array_top_bl1[0] array_top_bl1_n[0] array_top_bl2[0] array_top_bl2_n[0] array_top_bl1[1] array_top_bl1_n[1] array_top_bl2[1] array_top_bl2_n[1] array_top_bl1[2] array_top_bl1_n[2] array_top_bl2[2] array_top_bl2_n[2] array_top_bl1[3] array_top_bl1_n[3] array_top_bl2[3] array_top_bl2_n[3] bl1 bl1_n bl2 bl2_n array_top_bl1[5] array_top_bl1_n[5] array_top_bl2[5] array_top_bl2_n[5] array_top_bl1[6] array_top_bl1_n[6] array_top_bl2[6] array_top_bl2_n[6] array_top_bl1[7] array_top_bl1_n[7] array_top_bl2[7] array_top_bl2_n[7] DP8TVar14Array_6X8
Xzero vdd vss zero zero_x1
.ends DP8TVar14TestArray_16X8C

.subckt DP8TVar14 vss noco_vdd noco_wl1 noco_wl2 noco_bl1 noco_bl1_n noco_bl2 noco_bl2_n co_vdd co_bit co_bit_n co_wl1 co_wl2 co_bl1 co_bl1_n co_bl2_n co_bl2
Xframe noco_vdd noco_wl1 noco_wl2 noco_bl2 co_vdd co_bit co_bit_n co_wl1 co_wl2 NoConn_PAD0x9 vss noco_bl1 noco_bl1_n noco_bl2_n vss co_bl1 co_bl1_n co_bl2_n co_bl2 NoConn_PAD1x9 PadFrame_DP14
Xtestarray_noco vss noco_vdd noco_wl1 noco_wl2 noco_bl1 noco_bl1_n noco_bl2 noco_bl2_n DP8TVar14TestArray_16X8
Xtestarray_co vss co_vdd co_wl1 co_wl2 co_bl1 co_bl1_n co_bl2 co_bl2_n co_bit co_bit_n DP8TVar14TestArray_16X8C
.ends DP8TVar14

.subckt PadFrame_DP15 PAD0x0 PAD0x1 PAD0x2 PAD0x3 PAD0x4 PAD0x5 PAD0x6 PAD0x7 PAD0x8 PAD0x9 PAD1x0 PAD1x1 PAD1x2 PAD1x3 PAD1x4 PAD1x5 PAD1x6 PAD1x7 PAD1x8 PAD1x9
XPAD0x0 PAD0x0 BondPad
XPAD0x1 PAD0x1 BondPad
XPAD0x2 PAD0x2 BondPad
XPAD0x3 PAD0x3 BondPad
XPAD0x4 PAD0x4 BondPad
XPAD0x5 PAD0x5 BondPad
XPAD0x6 PAD0x6 BondPad
XPAD0x7 PAD0x7 BondPad
XPAD0x8 PAD0x8 BondPad
XPAD0x9 PAD0x9 BondPad
XPAD1x0 PAD1x0 BondPad
XPAD1x1 PAD1x1 BondPad
XPAD1x2 PAD1x2 BondPad
XPAD1x3 PAD1x3 BondPad
XPAD1x4 PAD1x4 BondPad
XPAD1x5 PAD1x5 BondPad
XPAD1x6 PAD1x6 BondPad
XPAD1x7 PAD1x7 BondPad
XPAD1x8 PAD1x8 BondPad
XPAD1x9 PAD1x9 BondPad
.ends PadFrame_DP15

.subckt DP8TVar15Cell wl1 wl2 bl1 bl1_n bl2 bl2_n vdd vss
Xpu1 vdd bit_n bit vdd sg13_lv_pmos l=1.3e-07 w=2e-07
Xpd1 bit bit_n vss vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpu2 vdd bit bit_n vdd sg13_lv_pmos l=1.3e-07 w=2e-07
Xpd2 bit_n bit vss vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg1 bit wl1 bl1 vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg1n bit_n wl1 bl1_n vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg2 bit wl2 bl2 vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg2n bit_n wl2 bl2_n vss sg13_lv_nmos l=1.3e-07 w=3e-07
.ends DP8TVar15Cell

.subckt DP8TVar15Array_2X1 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0]
Xinst0x0 wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] vdd vss DP8TVar15Cell
Xinst1x0 wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0] vdd vss DP8TVar15Cell
.ends DP8TVar15Array_2X1

.subckt DP8TVar15Array_2X2 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0] DP8TVar15Array_2X1
Xinst0x1 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TVar15Array_2X1
.ends DP8TVar15Array_2X2

.subckt DP8TVar15Array_4X2 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TVar15Array_2X2
Xinst1x0 vss vdd wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TVar15Array_2X2
.ends DP8TVar15Array_4X2

.subckt DP8TVar15Array_4X4 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TVar15Array_4X2
Xinst0x1 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar15Array_4X2
.ends DP8TVar15Array_4X4

.subckt DP8TVar15Array_8X4 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar15Array_4X4
Xinst1x0 vss vdd wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar15Array_4X4
.ends DP8TVar15Array_8X4

.subckt DP8TVar15Array_8X8 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar15Array_8X4
Xinst0x1 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar15Array_8X4
.ends DP8TVar15Array_8X8

.subckt DP8TVar15BulkConn vdd vss bl1 bl2 bl1_n bl2_n
.ends DP8TVar15BulkConn

.subckt DP8TVar15BulkConnRow_2 vss vdd bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1]
Xinst0 vdd vss bl1[0] bl2[0] bl1_n[0] bl2_n[0] DP8TVar15BulkConn
Xinst1 vdd vss bl1[1] bl2[1] bl1_n[1] bl2_n[1] DP8TVar15BulkConn
.ends DP8TVar15BulkConnRow_2

.subckt DP8TVar15BulkConnRow_4 vss vdd bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3]
Xinst0 vss vdd bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TVar15BulkConnRow_2
Xinst1 vss vdd bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar15BulkConnRow_2
.ends DP8TVar15BulkConnRow_4

.subckt DP8TVar15BulkConnRow_8 vss vdd bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0 vss vdd bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar15BulkConnRow_4
Xinst1 vss vdd bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar15BulkConnRow_4
.ends DP8TVar15BulkConnRow_8

.subckt DP8TVar15Array_16X8BC vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] wl1[8] wl2[8] wl1[9] wl2[9] wl1[10] wl2[10] wl1[11] wl2[11] wl1[12] wl2[12] wl1[13] wl2[13] wl1[14] wl2[14] wl1[15] wl2[15] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar15Array_8X8
Xinst1x0 vss vdd wl1[8] wl2[8] wl1[9] wl2[9] wl1[10] wl2[10] wl1[11] wl2[11] wl1[12] wl2[12] wl1[13] wl2[13] wl1[14] wl2[14] wl1[15] wl2[15] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar15Array_8X8
Xbottombcrow vss vdd bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar15BulkConnRow_8
Xtopbcrow vss vdd bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar15BulkConnRow_8
.ends DP8TVar15Array_16X8BC

.subckt DP8TVar15TestArray_16X8 vss vdd wl1 wl2 bl1 bl1_n bl2 bl2_n
Xarray vss vdd zero zero zero zero zero zero zero zero zero zero zero zero zero zero zero zero wl1 wl2 zero zero zero zero zero zero zero zero zero zero zero zero zero zero bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1 bl1_n bl2 bl2_n bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar15Array_16X8BC
Xzero vdd vss zero zero_x1
.ends DP8TVar15TestArray_16X8

.subckt DP8TVar15Array_4X8 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar15Array_4X4
Xinst0x1 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar15Array_4X4
.ends DP8TVar15Array_4X8

.subckt DP8TVar15Array_2X4 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TVar15Array_2X2
Xinst0x1 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar15Array_2X2
.ends DP8TVar15Array_2X4

.subckt DP8TVar15Array_2X8 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar15Array_2X4
Xinst0x1 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar15Array_2X4
.ends DP8TVar15Array_2X8

.subckt DP8TVar15Array_1X2 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1]
Xinst0x0 wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] vdd vss DP8TVar15Cell
Xinst0x1 wl1[0] wl2[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] vdd vss DP8TVar15Cell
.ends DP8TVar15Array_1X2

.subckt DP8TVar15Array_1X4 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3]
Xinst0x0 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TVar15Array_1X2
Xinst0x1 vss vdd wl1[0] wl2[0] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar15Array_1X2
.ends DP8TVar15Array_1X4

.subckt DP8TVar15Array_1X8 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar15Array_1X4
Xinst0x1 vss vdd wl1[0] wl2[0] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar15Array_1X4
.ends DP8TVar15Array_1X8

.subckt DP8TVar15Array_7X8 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar15Array_4X8
Xinst1x0 vss vdd wl1[4] wl2[4] wl1[5] wl2[5] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar15Array_2X8
Xinst2x0 vss vdd wl1[6] wl2[6] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar15Array_1X8
.ends DP8TVar15Array_7X8

.subckt DP8TVar15CellShWL1 wl1 wl2 bl1 bl1_n bl2 bl2_n vdd vss
Xpu1 vdd bit_n bit vdd sg13_lv_pmos l=1.3e-07 w=2e-07
Xpd1 bit bit_n vss vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpu2 vdd bit bit_n vdd sg13_lv_pmos l=1.3e-07 w=2e-07
Xpd2 bit_n bit vss vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg1 bit wl1 bl1 vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg1n bit_n wl1 bl1_n vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg2 bit wl1 bl2 vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg2n bit_n wl1 bl2_n vss sg13_lv_nmos l=1.3e-07 w=3e-07
.ends DP8TVar15CellShWL1

.subckt DP8TVar15ArrayShWL1_1X2 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1]
Xinst0x0 wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] vdd vss DP8TVar15CellShWL1
Xinst0x1 wl1[0] wl2[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] vdd vss DP8TVar15CellShWL1
.ends DP8TVar15ArrayShWL1_1X2

.subckt DP8TVar15ArrayShWL1_1X4 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3]
Xinst0x0 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TVar15ArrayShWL1_1X2
Xinst0x1 vss vdd wl1[0] wl2[0] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar15ArrayShWL1_1X2
.ends DP8TVar15ArrayShWL1_1X4

.subckt DP8TVar15ArrayShWL1_1X8 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar15ArrayShWL1_1X4
Xinst0x1 vss vdd wl1[0] wl2[0] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar15ArrayShWL1_1X4
.ends DP8TVar15ArrayShWL1_1X8

.subckt DP8TVar15CellConnectOut wl1 wl2 bl1 bl1_n bl2 bl2_n vdd vss bit bit_n
Xpu1 vdd bit_n bit vdd sg13_lv_pmos l=1.3e-07 w=2e-07
Xpd1 bit bit_n vss vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpu2 vdd bit bit_n vdd sg13_lv_pmos l=1.3e-07 w=2e-07
Xpd2 bit_n bit vss vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg1 bit wl1 bl1 vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg1n bit_n wl1 bl1_n vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg2 bit wl2 bl2 vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg2n bit_n wl2 bl2_n vss sg13_lv_nmos l=1.3e-07 w=3e-07
.ends DP8TVar15CellConnectOut

.subckt DP8TVar15CellShWL2 wl1 wl2 bl1 bl1_n bl2 bl2_n vdd vss
Xpu1 vdd bit_n bit vdd sg13_lv_pmos l=1.3e-07 w=2e-07
Xpd1 bit bit_n vss vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpu2 vdd bit bit_n vdd sg13_lv_pmos l=1.3e-07 w=2e-07
Xpd2 bit_n bit vss vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg1 bit wl2 bl1 vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg1n bit_n wl2 bl1_n vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg2 bit wl2 bl2 vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg2n bit_n wl2 bl2_n vss sg13_lv_nmos l=1.3e-07 w=3e-07
.ends DP8TVar15CellShWL2

.subckt DP8TVar15ArrayShWL2_1X2 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1]
Xinst0x0 wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] vdd vss DP8TVar15CellShWL2
Xinst0x1 wl1[0] wl2[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] vdd vss DP8TVar15CellShWL2
.ends DP8TVar15ArrayShWL2_1X2

.subckt DP8TVar15ArrayShWL2_1X4 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3]
Xinst0x0 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TVar15ArrayShWL2_1X2
Xinst0x1 vss vdd wl1[0] wl2[0] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar15ArrayShWL2_1X2
.ends DP8TVar15ArrayShWL2_1X4

.subckt DP8TVar15ArrayShWL2_1X8 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar15ArrayShWL2_1X4
Xinst0x1 vss vdd wl1[0] wl2[0] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar15ArrayShWL2_1X4
.ends DP8TVar15ArrayShWL2_1X8

.subckt DP8TVar15Array_6X8 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar15Array_4X8
Xinst1x0 vss vdd wl1[4] wl2[4] wl1[5] wl2[5] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar15Array_2X8
.ends DP8TVar15Array_6X8

.subckt DP8TVar15TestArray_16X8C vss vdd wl1 wl2 bl1 bl1_n bl2 bl2_n bit bit_n
Xbcconn_bot vss vdd bcconn_bot_bl1[0] bcconn_bot_bl1_n[0] bcconn_bot_bl2[0] bcconn_bot_bl2_n[0] bcconn_bot_bl1[1] bcconn_bot_bl1_n[1] bcconn_bot_bl2[1] bcconn_bot_bl2_n[1] bcconn_bot_bl1[2] bcconn_bot_bl1_n[2] bcconn_bot_bl2[2] bcconn_bot_bl2_n[2] bcconn_bot_bl1[3] bcconn_bot_bl1_n[3] bcconn_bot_bl2[3] bcconn_bot_bl2_n[3] bl1 bl1_n bl2 bl2_n bcconn_bot_bl1[5] bcconn_bot_bl1_n[5] bcconn_bot_bl2[5] bcconn_bot_bl2_n[5] bcconn_bot_bl1[6] bcconn_bot_bl1_n[6] bcconn_bot_bl2[6] bcconn_bot_bl2_n[6] bcconn_bot_bl1[7] bcconn_bot_bl1_n[7] bcconn_bot_bl2[7] bcconn_bot_bl2_n[7] DP8TVar15BulkConnRow_8
Xbcconn_top vss vdd bcconn_top_bl1[0] bcconn_top_bl1_n[0] bcconn_top_bl2[0] bcconn_top_bl2_n[0] bcconn_top_bl1[1] bcconn_top_bl1_n[1] bcconn_top_bl2[1] bcconn_top_bl2_n[1] bcconn_top_bl1[2] bcconn_top_bl1_n[2] bcconn_top_bl2[2] bcconn_top_bl2_n[2] bcconn_top_bl1[3] bcconn_top_bl1_n[3] bcconn_top_bl2[3] bcconn_top_bl2_n[3] bl1 bl1_n bl2 bl2_n bcconn_top_bl1[5] bcconn_top_bl1_n[5] bcconn_top_bl2[5] bcconn_top_bl2_n[5] bcconn_top_bl1[6] bcconn_top_bl1_n[6] bcconn_top_bl2[6] bcconn_top_bl2_n[6] bcconn_top_bl1[7] bcconn_top_bl1_n[7] bcconn_top_bl2[7] bcconn_top_bl2_n[7] DP8TVar15BulkConnRow_8
Xarray_bot vss vdd zero zero zero zero zero zero zero zero zero zero zero zero zero zero array_bot_bl1[0] array_bot_bl1_n[0] array_bot_bl2[0] array_bot_bl2_n[0] array_bot_bl1[1] array_bot_bl1_n[1] array_bot_bl2[1] array_bot_bl2_n[1] array_bot_bl1[2] array_bot_bl1_n[2] array_bot_bl2[2] array_bot_bl2_n[2] array_bot_bl1[3] array_bot_bl1_n[3] array_bot_bl2[3] array_bot_bl2_n[3] bl1 bl1_n bl2 bl2_n array_bot_bl1[5] array_bot_bl1_n[5] array_bot_bl2[5] array_bot_bl2_n[5] array_bot_bl1[6] array_bot_bl1_n[6] array_bot_bl2[6] array_bot_bl2_n[6] array_bot_bl1[7] array_bot_bl1_n[7] array_bot_bl2[7] array_bot_bl2_n[7] DP8TVar15Array_7X8
Xshwl1_row vss vdd zero bit shwl1_row_bl1[0] shwl1_row_bl1_n[0] shwl1_row_bl2[0] shwl1_row_bl2_n[0] shwl1_row_bl1[1] shwl1_row_bl1_n[1] shwl1_row_bl2[1] shwl1_row_bl2_n[1] shwl1_row_bl1[2] shwl1_row_bl1_n[2] shwl1_row_bl2[2] shwl1_row_bl2_n[2] shwl1_row_bl1[3] shwl1_row_bl1_n[3] shwl1_row_bl2[3] shwl1_row_bl2_n[3] bl1 bl1_n bl2 bl2_n shwl1_row_bl1[5] shwl1_row_bl1_n[5] shwl1_row_bl2[5] shwl1_row_bl2_n[5] shwl1_row_bl1[6] shwl1_row_bl1_n[6] shwl1_row_bl2[6] shwl1_row_bl2_n[6] shwl1_row_bl1[7] shwl1_row_bl1_n[7] shwl1_row_bl2[7] shwl1_row_bl2_n[7] DP8TVar15ArrayShWL1_1X8
Xcell_cols_left vss vdd wl1 wl2 cell_cols_left_bl1[0] cell_cols_left_bl1_n[0] cell_cols_left_bl2[0] cell_cols_left_bl2_n[0] cell_cols_left_bl1[1] cell_cols_left_bl1_n[1] cell_cols_left_bl2[1] cell_cols_left_bl2_n[1] cell_cols_left_bl1[2] cell_cols_left_bl1_n[2] cell_cols_left_bl2[2] cell_cols_left_bl2_n[2] cell_cols_left_bl1[3] cell_cols_left_bl1_n[3] cell_cols_left_bl2[3] cell_cols_left_bl2_n[3] DP8TVar15Array_1X4
Xconncell wl1 wl2 bl1 bl1_n bl2 bl2_n vdd vss bit bit_n DP8TVar15CellConnectOut
Xfillcell wl1 wl2 fillcell_bl1 fillcell_bl1_n fillcell_bl2 fillcell_bl2_n vdd vss DP8TVar15Cell
Xcell_cols_right vss vdd wl1 wl2 cell_cols_right_bl1[0] cell_cols_right_bl1_n[0] cell_cols_right_bl2[0] cell_cols_right_bl2_n[0] cell_cols_right_bl1[1] cell_cols_right_bl1_n[1] cell_cols_right_bl2[1] cell_cols_right_bl2_n[1] DP8TVar15Array_1X2
Xshwl2_row vss vdd bit_n zero shwl2_row_bl1[0] shwl2_row_bl1_n[0] shwl2_row_bl2[0] shwl2_row_bl2_n[0] shwl2_row_bl1[1] shwl2_row_bl1_n[1] shwl2_row_bl2[1] shwl2_row_bl2_n[1] shwl2_row_bl1[2] shwl2_row_bl1_n[2] shwl2_row_bl2[2] shwl2_row_bl2_n[2] shwl2_row_bl1[3] shwl2_row_bl1_n[3] shwl2_row_bl2[3] shwl2_row_bl2_n[3] bl1 bl1_n bl2 bl2_n shwl2_row_bl1[5] shwl2_row_bl1_n[5] shwl2_row_bl2[5] shwl2_row_bl2_n[5] shwl2_row_bl1[6] shwl2_row_bl1_n[6] shwl2_row_bl2[6] shwl2_row_bl2_n[6] shwl2_row_bl1[7] shwl2_row_bl1_n[7] shwl2_row_bl2[7] shwl2_row_bl2_n[7] DP8TVar15ArrayShWL2_1X8
Xarray_top vss vdd zero zero zero zero zero zero zero zero zero zero zero zero array_top_bl1[0] array_top_bl1_n[0] array_top_bl2[0] array_top_bl2_n[0] array_top_bl1[1] array_top_bl1_n[1] array_top_bl2[1] array_top_bl2_n[1] array_top_bl1[2] array_top_bl1_n[2] array_top_bl2[2] array_top_bl2_n[2] array_top_bl1[3] array_top_bl1_n[3] array_top_bl2[3] array_top_bl2_n[3] bl1 bl1_n bl2 bl2_n array_top_bl1[5] array_top_bl1_n[5] array_top_bl2[5] array_top_bl2_n[5] array_top_bl1[6] array_top_bl1_n[6] array_top_bl2[6] array_top_bl2_n[6] array_top_bl1[7] array_top_bl1_n[7] array_top_bl2[7] array_top_bl2_n[7] DP8TVar15Array_6X8
Xzero vdd vss zero zero_x1
.ends DP8TVar15TestArray_16X8C

.subckt DP8TVar15 vss noco_vdd noco_wl1 noco_wl2 noco_bl1 noco_bl1_n noco_bl2 noco_bl2_n co_vdd co_bit co_bit_n co_wl1 co_wl2 co_bl1 co_bl1_n co_bl2_n co_bl2
Xframe noco_vdd noco_wl1 noco_wl2 noco_bl2 co_vdd co_bit co_bit_n co_wl1 co_wl2 NoConn_PAD0x9 vss noco_bl1 noco_bl1_n noco_bl2_n vss co_bl1 co_bl1_n co_bl2_n co_bl2 NoConn_PAD1x9 PadFrame_DP15
Xtestarray_noco vss noco_vdd noco_wl1 noco_wl2 noco_bl1 noco_bl1_n noco_bl2 noco_bl2_n DP8TVar15TestArray_16X8
Xtestarray_co vss co_vdd co_wl1 co_wl2 co_bl1 co_bl1_n co_bl2 co_bl2_n co_bit co_bit_n DP8TVar15TestArray_16X8C
.ends DP8TVar15

.subckt PadFrame_DP16 PAD0x0 PAD0x1 PAD0x2 PAD0x3 PAD0x4 PAD0x5 PAD0x6 PAD0x7 PAD0x8 PAD0x9 PAD1x0 PAD1x1 PAD1x2 PAD1x3 PAD1x4 PAD1x5 PAD1x6 PAD1x7 PAD1x8 PAD1x9
XPAD0x0 PAD0x0 BondPad
XPAD0x1 PAD0x1 BondPad
XPAD0x2 PAD0x2 BondPad
XPAD0x3 PAD0x3 BondPad
XPAD0x4 PAD0x4 BondPad
XPAD0x5 PAD0x5 BondPad
XPAD0x6 PAD0x6 BondPad
XPAD0x7 PAD0x7 BondPad
XPAD0x8 PAD0x8 BondPad
XPAD0x9 PAD0x9 BondPad
XPAD1x0 PAD1x0 BondPad
XPAD1x1 PAD1x1 BondPad
XPAD1x2 PAD1x2 BondPad
XPAD1x3 PAD1x3 BondPad
XPAD1x4 PAD1x4 BondPad
XPAD1x5 PAD1x5 BondPad
XPAD1x6 PAD1x6 BondPad
XPAD1x7 PAD1x7 BondPad
XPAD1x8 PAD1x8 BondPad
XPAD1x9 PAD1x9 BondPad
.ends PadFrame_DP16

.subckt DP8TVar16Cell wl1 wl2 bl1 bl1_n bl2 bl2_n vdd vss
Xpu1 vdd bit_n bit vdd sg13_lv_pmos l=1.3e-07 w=1.5e-07
Xpd1 bit bit_n vss vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpu2 vdd bit bit_n vdd sg13_lv_pmos l=1.3e-07 w=1.5e-07
Xpd2 bit_n bit vss vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg1 bit wl1 bl1 vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg1n bit_n wl1 bl1_n vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg2 bit wl2 bl2 vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg2n bit_n wl2 bl2_n vss sg13_lv_nmos l=1.3e-07 w=3e-07
.ends DP8TVar16Cell

.subckt DP8TVar16Array_2X1 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0]
Xinst0x0 wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] vdd vss DP8TVar16Cell
Xinst1x0 wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0] vdd vss DP8TVar16Cell
.ends DP8TVar16Array_2X1

.subckt DP8TVar16Array_2X2 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0] DP8TVar16Array_2X1
Xinst0x1 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TVar16Array_2X1
.ends DP8TVar16Array_2X2

.subckt DP8TVar16Array_4X2 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TVar16Array_2X2
Xinst1x0 vss vdd wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TVar16Array_2X2
.ends DP8TVar16Array_4X2

.subckt DP8TVar16Array_4X4 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TVar16Array_4X2
Xinst0x1 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar16Array_4X2
.ends DP8TVar16Array_4X4

.subckt DP8TVar16Array_8X4 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar16Array_4X4
Xinst1x0 vss vdd wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar16Array_4X4
.ends DP8TVar16Array_8X4

.subckt DP8TVar16Array_8X8 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar16Array_8X4
Xinst0x1 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar16Array_8X4
.ends DP8TVar16Array_8X8

.subckt DP8TVar16BulkConn vdd vss bl1 bl2 bl1_n bl2_n
.ends DP8TVar16BulkConn

.subckt DP8TVar16BulkConnRow_2 vss vdd bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1]
Xinst0 vdd vss bl1[0] bl2[0] bl1_n[0] bl2_n[0] DP8TVar16BulkConn
Xinst1 vdd vss bl1[1] bl2[1] bl1_n[1] bl2_n[1] DP8TVar16BulkConn
.ends DP8TVar16BulkConnRow_2

.subckt DP8TVar16BulkConnRow_4 vss vdd bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3]
Xinst0 vss vdd bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TVar16BulkConnRow_2
Xinst1 vss vdd bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar16BulkConnRow_2
.ends DP8TVar16BulkConnRow_4

.subckt DP8TVar16BulkConnRow_8 vss vdd bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0 vss vdd bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar16BulkConnRow_4
Xinst1 vss vdd bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar16BulkConnRow_4
.ends DP8TVar16BulkConnRow_8

.subckt DP8TVar16Array_16X8BC vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] wl1[8] wl2[8] wl1[9] wl2[9] wl1[10] wl2[10] wl1[11] wl2[11] wl1[12] wl2[12] wl1[13] wl2[13] wl1[14] wl2[14] wl1[15] wl2[15] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar16Array_8X8
Xinst1x0 vss vdd wl1[8] wl2[8] wl1[9] wl2[9] wl1[10] wl2[10] wl1[11] wl2[11] wl1[12] wl2[12] wl1[13] wl2[13] wl1[14] wl2[14] wl1[15] wl2[15] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar16Array_8X8
Xbottombcrow vss vdd bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar16BulkConnRow_8
Xtopbcrow vss vdd bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar16BulkConnRow_8
.ends DP8TVar16Array_16X8BC

.subckt DP8TVar16TestArray_16X8 vss vdd wl1 wl2 bl1 bl1_n bl2 bl2_n
Xarray vss vdd zero zero zero zero zero zero zero zero zero zero zero zero zero zero zero zero wl1 wl2 zero zero zero zero zero zero zero zero zero zero zero zero zero zero bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1 bl1_n bl2 bl2_n bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar16Array_16X8BC
Xzero vdd vss zero zero_x1
.ends DP8TVar16TestArray_16X8

.subckt DP8TVar16Array_4X8 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar16Array_4X4
Xinst0x1 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar16Array_4X4
.ends DP8TVar16Array_4X8

.subckt DP8TVar16Array_2X4 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TVar16Array_2X2
Xinst0x1 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar16Array_2X2
.ends DP8TVar16Array_2X4

.subckt DP8TVar16Array_2X8 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar16Array_2X4
Xinst0x1 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar16Array_2X4
.ends DP8TVar16Array_2X8

.subckt DP8TVar16Array_1X2 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1]
Xinst0x0 wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] vdd vss DP8TVar16Cell
Xinst0x1 wl1[0] wl2[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] vdd vss DP8TVar16Cell
.ends DP8TVar16Array_1X2

.subckt DP8TVar16Array_1X4 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3]
Xinst0x0 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TVar16Array_1X2
Xinst0x1 vss vdd wl1[0] wl2[0] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar16Array_1X2
.ends DP8TVar16Array_1X4

.subckt DP8TVar16Array_1X8 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar16Array_1X4
Xinst0x1 vss vdd wl1[0] wl2[0] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar16Array_1X4
.ends DP8TVar16Array_1X8

.subckt DP8TVar16Array_7X8 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar16Array_4X8
Xinst1x0 vss vdd wl1[4] wl2[4] wl1[5] wl2[5] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar16Array_2X8
Xinst2x0 vss vdd wl1[6] wl2[6] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar16Array_1X8
.ends DP8TVar16Array_7X8

.subckt DP8TVar16CellShWL1 wl1 wl2 bl1 bl1_n bl2 bl2_n vdd vss
Xpu1 vdd bit_n bit vdd sg13_lv_pmos l=1.3e-07 w=1.5e-07
Xpd1 bit bit_n vss vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpu2 vdd bit bit_n vdd sg13_lv_pmos l=1.3e-07 w=1.5e-07
Xpd2 bit_n bit vss vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg1 bit wl1 bl1 vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg1n bit_n wl1 bl1_n vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg2 bit wl1 bl2 vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg2n bit_n wl1 bl2_n vss sg13_lv_nmos l=1.3e-07 w=3e-07
.ends DP8TVar16CellShWL1

.subckt DP8TVar16ArrayShWL1_1X2 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1]
Xinst0x0 wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] vdd vss DP8TVar16CellShWL1
Xinst0x1 wl1[0] wl2[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] vdd vss DP8TVar16CellShWL1
.ends DP8TVar16ArrayShWL1_1X2

.subckt DP8TVar16ArrayShWL1_1X4 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3]
Xinst0x0 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TVar16ArrayShWL1_1X2
Xinst0x1 vss vdd wl1[0] wl2[0] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar16ArrayShWL1_1X2
.ends DP8TVar16ArrayShWL1_1X4

.subckt DP8TVar16ArrayShWL1_1X8 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar16ArrayShWL1_1X4
Xinst0x1 vss vdd wl1[0] wl2[0] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar16ArrayShWL1_1X4
.ends DP8TVar16ArrayShWL1_1X8

.subckt DP8TVar16CellConnectOut wl1 wl2 bl1 bl1_n bl2 bl2_n vdd vss bit bit_n
Xpu1 vdd bit_n bit vdd sg13_lv_pmos l=1.3e-07 w=1.5e-07
Xpd1 bit bit_n vss vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpu2 vdd bit bit_n vdd sg13_lv_pmos l=1.3e-07 w=1.5e-07
Xpd2 bit_n bit vss vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg1 bit wl1 bl1 vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg1n bit_n wl1 bl1_n vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg2 bit wl2 bl2 vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg2n bit_n wl2 bl2_n vss sg13_lv_nmos l=1.3e-07 w=3e-07
.ends DP8TVar16CellConnectOut

.subckt DP8TVar16CellShWL2 wl1 wl2 bl1 bl1_n bl2 bl2_n vdd vss
Xpu1 vdd bit_n bit vdd sg13_lv_pmos l=1.3e-07 w=1.5e-07
Xpd1 bit bit_n vss vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpu2 vdd bit bit_n vdd sg13_lv_pmos l=1.3e-07 w=1.5e-07
Xpd2 bit_n bit vss vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg1 bit wl2 bl1 vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg1n bit_n wl2 bl1_n vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg2 bit wl2 bl2 vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg2n bit_n wl2 bl2_n vss sg13_lv_nmos l=1.3e-07 w=3e-07
.ends DP8TVar16CellShWL2

.subckt DP8TVar16ArrayShWL2_1X2 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1]
Xinst0x0 wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] vdd vss DP8TVar16CellShWL2
Xinst0x1 wl1[0] wl2[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] vdd vss DP8TVar16CellShWL2
.ends DP8TVar16ArrayShWL2_1X2

.subckt DP8TVar16ArrayShWL2_1X4 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3]
Xinst0x0 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TVar16ArrayShWL2_1X2
Xinst0x1 vss vdd wl1[0] wl2[0] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar16ArrayShWL2_1X2
.ends DP8TVar16ArrayShWL2_1X4

.subckt DP8TVar16ArrayShWL2_1X8 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar16ArrayShWL2_1X4
Xinst0x1 vss vdd wl1[0] wl2[0] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar16ArrayShWL2_1X4
.ends DP8TVar16ArrayShWL2_1X8

.subckt DP8TVar16Array_6X8 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar16Array_4X8
Xinst1x0 vss vdd wl1[4] wl2[4] wl1[5] wl2[5] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar16Array_2X8
.ends DP8TVar16Array_6X8

.subckt DP8TVar16TestArray_16X8C vss vdd wl1 wl2 bl1 bl1_n bl2 bl2_n bit bit_n
Xbcconn_bot vss vdd bcconn_bot_bl1[0] bcconn_bot_bl1_n[0] bcconn_bot_bl2[0] bcconn_bot_bl2_n[0] bcconn_bot_bl1[1] bcconn_bot_bl1_n[1] bcconn_bot_bl2[1] bcconn_bot_bl2_n[1] bcconn_bot_bl1[2] bcconn_bot_bl1_n[2] bcconn_bot_bl2[2] bcconn_bot_bl2_n[2] bcconn_bot_bl1[3] bcconn_bot_bl1_n[3] bcconn_bot_bl2[3] bcconn_bot_bl2_n[3] bl1 bl1_n bl2 bl2_n bcconn_bot_bl1[5] bcconn_bot_bl1_n[5] bcconn_bot_bl2[5] bcconn_bot_bl2_n[5] bcconn_bot_bl1[6] bcconn_bot_bl1_n[6] bcconn_bot_bl2[6] bcconn_bot_bl2_n[6] bcconn_bot_bl1[7] bcconn_bot_bl1_n[7] bcconn_bot_bl2[7] bcconn_bot_bl2_n[7] DP8TVar16BulkConnRow_8
Xbcconn_top vss vdd bcconn_top_bl1[0] bcconn_top_bl1_n[0] bcconn_top_bl2[0] bcconn_top_bl2_n[0] bcconn_top_bl1[1] bcconn_top_bl1_n[1] bcconn_top_bl2[1] bcconn_top_bl2_n[1] bcconn_top_bl1[2] bcconn_top_bl1_n[2] bcconn_top_bl2[2] bcconn_top_bl2_n[2] bcconn_top_bl1[3] bcconn_top_bl1_n[3] bcconn_top_bl2[3] bcconn_top_bl2_n[3] bl1 bl1_n bl2 bl2_n bcconn_top_bl1[5] bcconn_top_bl1_n[5] bcconn_top_bl2[5] bcconn_top_bl2_n[5] bcconn_top_bl1[6] bcconn_top_bl1_n[6] bcconn_top_bl2[6] bcconn_top_bl2_n[6] bcconn_top_bl1[7] bcconn_top_bl1_n[7] bcconn_top_bl2[7] bcconn_top_bl2_n[7] DP8TVar16BulkConnRow_8
Xarray_bot vss vdd zero zero zero zero zero zero zero zero zero zero zero zero zero zero array_bot_bl1[0] array_bot_bl1_n[0] array_bot_bl2[0] array_bot_bl2_n[0] array_bot_bl1[1] array_bot_bl1_n[1] array_bot_bl2[1] array_bot_bl2_n[1] array_bot_bl1[2] array_bot_bl1_n[2] array_bot_bl2[2] array_bot_bl2_n[2] array_bot_bl1[3] array_bot_bl1_n[3] array_bot_bl2[3] array_bot_bl2_n[3] bl1 bl1_n bl2 bl2_n array_bot_bl1[5] array_bot_bl1_n[5] array_bot_bl2[5] array_bot_bl2_n[5] array_bot_bl1[6] array_bot_bl1_n[6] array_bot_bl2[6] array_bot_bl2_n[6] array_bot_bl1[7] array_bot_bl1_n[7] array_bot_bl2[7] array_bot_bl2_n[7] DP8TVar16Array_7X8
Xshwl1_row vss vdd zero bit shwl1_row_bl1[0] shwl1_row_bl1_n[0] shwl1_row_bl2[0] shwl1_row_bl2_n[0] shwl1_row_bl1[1] shwl1_row_bl1_n[1] shwl1_row_bl2[1] shwl1_row_bl2_n[1] shwl1_row_bl1[2] shwl1_row_bl1_n[2] shwl1_row_bl2[2] shwl1_row_bl2_n[2] shwl1_row_bl1[3] shwl1_row_bl1_n[3] shwl1_row_bl2[3] shwl1_row_bl2_n[3] bl1 bl1_n bl2 bl2_n shwl1_row_bl1[5] shwl1_row_bl1_n[5] shwl1_row_bl2[5] shwl1_row_bl2_n[5] shwl1_row_bl1[6] shwl1_row_bl1_n[6] shwl1_row_bl2[6] shwl1_row_bl2_n[6] shwl1_row_bl1[7] shwl1_row_bl1_n[7] shwl1_row_bl2[7] shwl1_row_bl2_n[7] DP8TVar16ArrayShWL1_1X8
Xcell_cols_left vss vdd wl1 wl2 cell_cols_left_bl1[0] cell_cols_left_bl1_n[0] cell_cols_left_bl2[0] cell_cols_left_bl2_n[0] cell_cols_left_bl1[1] cell_cols_left_bl1_n[1] cell_cols_left_bl2[1] cell_cols_left_bl2_n[1] cell_cols_left_bl1[2] cell_cols_left_bl1_n[2] cell_cols_left_bl2[2] cell_cols_left_bl2_n[2] cell_cols_left_bl1[3] cell_cols_left_bl1_n[3] cell_cols_left_bl2[3] cell_cols_left_bl2_n[3] DP8TVar16Array_1X4
Xconncell wl1 wl2 bl1 bl1_n bl2 bl2_n vdd vss bit bit_n DP8TVar16CellConnectOut
Xfillcell wl1 wl2 fillcell_bl1 fillcell_bl1_n fillcell_bl2 fillcell_bl2_n vdd vss DP8TVar16Cell
Xcell_cols_right vss vdd wl1 wl2 cell_cols_right_bl1[0] cell_cols_right_bl1_n[0] cell_cols_right_bl2[0] cell_cols_right_bl2_n[0] cell_cols_right_bl1[1] cell_cols_right_bl1_n[1] cell_cols_right_bl2[1] cell_cols_right_bl2_n[1] DP8TVar16Array_1X2
Xshwl2_row vss vdd bit_n zero shwl2_row_bl1[0] shwl2_row_bl1_n[0] shwl2_row_bl2[0] shwl2_row_bl2_n[0] shwl2_row_bl1[1] shwl2_row_bl1_n[1] shwl2_row_bl2[1] shwl2_row_bl2_n[1] shwl2_row_bl1[2] shwl2_row_bl1_n[2] shwl2_row_bl2[2] shwl2_row_bl2_n[2] shwl2_row_bl1[3] shwl2_row_bl1_n[3] shwl2_row_bl2[3] shwl2_row_bl2_n[3] bl1 bl1_n bl2 bl2_n shwl2_row_bl1[5] shwl2_row_bl1_n[5] shwl2_row_bl2[5] shwl2_row_bl2_n[5] shwl2_row_bl1[6] shwl2_row_bl1_n[6] shwl2_row_bl2[6] shwl2_row_bl2_n[6] shwl2_row_bl1[7] shwl2_row_bl1_n[7] shwl2_row_bl2[7] shwl2_row_bl2_n[7] DP8TVar16ArrayShWL2_1X8
Xarray_top vss vdd zero zero zero zero zero zero zero zero zero zero zero zero array_top_bl1[0] array_top_bl1_n[0] array_top_bl2[0] array_top_bl2_n[0] array_top_bl1[1] array_top_bl1_n[1] array_top_bl2[1] array_top_bl2_n[1] array_top_bl1[2] array_top_bl1_n[2] array_top_bl2[2] array_top_bl2_n[2] array_top_bl1[3] array_top_bl1_n[3] array_top_bl2[3] array_top_bl2_n[3] bl1 bl1_n bl2 bl2_n array_top_bl1[5] array_top_bl1_n[5] array_top_bl2[5] array_top_bl2_n[5] array_top_bl1[6] array_top_bl1_n[6] array_top_bl2[6] array_top_bl2_n[6] array_top_bl1[7] array_top_bl1_n[7] array_top_bl2[7] array_top_bl2_n[7] DP8TVar16Array_6X8
Xzero vdd vss zero zero_x1
.ends DP8TVar16TestArray_16X8C

.subckt DP8TVar16 vss noco_vdd noco_wl1 noco_wl2 noco_bl1 noco_bl1_n noco_bl2 noco_bl2_n co_vdd co_bit co_bit_n co_wl1 co_wl2 co_bl1 co_bl1_n co_bl2_n co_bl2
Xframe noco_vdd noco_wl1 noco_wl2 noco_bl2 co_vdd co_bit co_bit_n co_wl1 co_wl2 NoConn_PAD0x9 vss noco_bl1 noco_bl1_n noco_bl2_n vss co_bl1 co_bl1_n co_bl2_n co_bl2 NoConn_PAD1x9 PadFrame_DP16
Xtestarray_noco vss noco_vdd noco_wl1 noco_wl2 noco_bl1 noco_bl1_n noco_bl2 noco_bl2_n DP8TVar16TestArray_16X8
Xtestarray_co vss co_vdd co_wl1 co_wl2 co_bl1 co_bl1_n co_bl2 co_bl2_n co_bit co_bit_n DP8TVar16TestArray_16X8C
.ends DP8TVar16

.subckt PadFrame_DP17 PAD0x0 PAD0x1 PAD0x2 PAD0x3 PAD0x4 PAD0x5 PAD0x6 PAD0x7 PAD0x8 PAD0x9 PAD1x0 PAD1x1 PAD1x2 PAD1x3 PAD1x4 PAD1x5 PAD1x6 PAD1x7 PAD1x8 PAD1x9
XPAD0x0 PAD0x0 BondPad
XPAD0x1 PAD0x1 BondPad
XPAD0x2 PAD0x2 BondPad
XPAD0x3 PAD0x3 BondPad
XPAD0x4 PAD0x4 BondPad
XPAD0x5 PAD0x5 BondPad
XPAD0x6 PAD0x6 BondPad
XPAD0x7 PAD0x7 BondPad
XPAD0x8 PAD0x8 BondPad
XPAD0x9 PAD0x9 BondPad
XPAD1x0 PAD1x0 BondPad
XPAD1x1 PAD1x1 BondPad
XPAD1x2 PAD1x2 BondPad
XPAD1x3 PAD1x3 BondPad
XPAD1x4 PAD1x4 BondPad
XPAD1x5 PAD1x5 BondPad
XPAD1x6 PAD1x6 BondPad
XPAD1x7 PAD1x7 BondPad
XPAD1x8 PAD1x8 BondPad
XPAD1x9 PAD1x9 BondPad
.ends PadFrame_DP17

.subckt DP8TVar17Cell wl1 wl2 bl1 bl1_n bl2 bl2_n vdd vss
Xpu1 vdd bit_n bit vdd sg13_lv_pmos l=1.3e-07 w=2e-07
Xpd1 bit bit_n vss vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpu2 vdd bit bit_n vdd sg13_lv_pmos l=1.3e-07 w=2e-07
Xpd2 bit_n bit vss vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg1 bit wl1 bl1 vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg1n bit_n wl1 bl1_n vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg2 bit wl2 bl2 vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg2n bit_n wl2 bl2_n vss sg13_lv_nmos l=1.3e-07 w=2e-07
.ends DP8TVar17Cell

.subckt DP8TVar17Array_2X1 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0]
Xinst0x0 wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] vdd vss DP8TVar17Cell
Xinst1x0 wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0] vdd vss DP8TVar17Cell
.ends DP8TVar17Array_2X1

.subckt DP8TVar17Array_2X2 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0] DP8TVar17Array_2X1
Xinst0x1 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TVar17Array_2X1
.ends DP8TVar17Array_2X2

.subckt DP8TVar17Array_4X2 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TVar17Array_2X2
Xinst1x0 vss vdd wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TVar17Array_2X2
.ends DP8TVar17Array_4X2

.subckt DP8TVar17Array_4X4 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TVar17Array_4X2
Xinst0x1 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar17Array_4X2
.ends DP8TVar17Array_4X4

.subckt DP8TVar17Array_8X4 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar17Array_4X4
Xinst1x0 vss vdd wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar17Array_4X4
.ends DP8TVar17Array_8X4

.subckt DP8TVar17Array_8X8 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar17Array_8X4
Xinst0x1 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar17Array_8X4
.ends DP8TVar17Array_8X8

.subckt DP8TVar17BulkConn vdd vss bl1 bl2 bl1_n bl2_n
.ends DP8TVar17BulkConn

.subckt DP8TVar17BulkConnRow_2 vss vdd bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1]
Xinst0 vdd vss bl1[0] bl2[0] bl1_n[0] bl2_n[0] DP8TVar17BulkConn
Xinst1 vdd vss bl1[1] bl2[1] bl1_n[1] bl2_n[1] DP8TVar17BulkConn
.ends DP8TVar17BulkConnRow_2

.subckt DP8TVar17BulkConnRow_4 vss vdd bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3]
Xinst0 vss vdd bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TVar17BulkConnRow_2
Xinst1 vss vdd bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar17BulkConnRow_2
.ends DP8TVar17BulkConnRow_4

.subckt DP8TVar17BulkConnRow_8 vss vdd bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0 vss vdd bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar17BulkConnRow_4
Xinst1 vss vdd bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar17BulkConnRow_4
.ends DP8TVar17BulkConnRow_8

.subckt DP8TVar17Array_16X8BC vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] wl1[8] wl2[8] wl1[9] wl2[9] wl1[10] wl2[10] wl1[11] wl2[11] wl1[12] wl2[12] wl1[13] wl2[13] wl1[14] wl2[14] wl1[15] wl2[15] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar17Array_8X8
Xinst1x0 vss vdd wl1[8] wl2[8] wl1[9] wl2[9] wl1[10] wl2[10] wl1[11] wl2[11] wl1[12] wl2[12] wl1[13] wl2[13] wl1[14] wl2[14] wl1[15] wl2[15] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar17Array_8X8
Xbottombcrow vss vdd bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar17BulkConnRow_8
Xtopbcrow vss vdd bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar17BulkConnRow_8
.ends DP8TVar17Array_16X8BC

.subckt DP8TVar17TestArray_16X8 vss vdd wl1 wl2 bl1 bl1_n bl2 bl2_n
Xarray vss vdd zero zero zero zero zero zero zero zero zero zero zero zero zero zero zero zero wl1 wl2 zero zero zero zero zero zero zero zero zero zero zero zero zero zero bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1 bl1_n bl2 bl2_n bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar17Array_16X8BC
Xzero vdd vss zero zero_x1
.ends DP8TVar17TestArray_16X8

.subckt DP8TVar17Array_4X8 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar17Array_4X4
Xinst0x1 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar17Array_4X4
.ends DP8TVar17Array_4X8

.subckt DP8TVar17Array_2X4 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TVar17Array_2X2
Xinst0x1 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar17Array_2X2
.ends DP8TVar17Array_2X4

.subckt DP8TVar17Array_2X8 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar17Array_2X4
Xinst0x1 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar17Array_2X4
.ends DP8TVar17Array_2X8

.subckt DP8TVar17Array_1X2 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1]
Xinst0x0 wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] vdd vss DP8TVar17Cell
Xinst0x1 wl1[0] wl2[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] vdd vss DP8TVar17Cell
.ends DP8TVar17Array_1X2

.subckt DP8TVar17Array_1X4 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3]
Xinst0x0 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TVar17Array_1X2
Xinst0x1 vss vdd wl1[0] wl2[0] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar17Array_1X2
.ends DP8TVar17Array_1X4

.subckt DP8TVar17Array_1X8 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar17Array_1X4
Xinst0x1 vss vdd wl1[0] wl2[0] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar17Array_1X4
.ends DP8TVar17Array_1X8

.subckt DP8TVar17Array_7X8 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar17Array_4X8
Xinst1x0 vss vdd wl1[4] wl2[4] wl1[5] wl2[5] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar17Array_2X8
Xinst2x0 vss vdd wl1[6] wl2[6] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar17Array_1X8
.ends DP8TVar17Array_7X8

.subckt DP8TVar17CellShWL1 wl1 wl2 bl1 bl1_n bl2 bl2_n vdd vss
Xpu1 vdd bit_n bit vdd sg13_lv_pmos l=1.3e-07 w=2e-07
Xpd1 bit bit_n vss vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpu2 vdd bit bit_n vdd sg13_lv_pmos l=1.3e-07 w=2e-07
Xpd2 bit_n bit vss vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg1 bit wl1 bl1 vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg1n bit_n wl1 bl1_n vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg2 bit wl1 bl2 vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg2n bit_n wl1 bl2_n vss sg13_lv_nmos l=1.3e-07 w=2e-07
.ends DP8TVar17CellShWL1

.subckt DP8TVar17ArrayShWL1_1X2 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1]
Xinst0x0 wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] vdd vss DP8TVar17CellShWL1
Xinst0x1 wl1[0] wl2[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] vdd vss DP8TVar17CellShWL1
.ends DP8TVar17ArrayShWL1_1X2

.subckt DP8TVar17ArrayShWL1_1X4 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3]
Xinst0x0 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TVar17ArrayShWL1_1X2
Xinst0x1 vss vdd wl1[0] wl2[0] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar17ArrayShWL1_1X2
.ends DP8TVar17ArrayShWL1_1X4

.subckt DP8TVar17ArrayShWL1_1X8 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar17ArrayShWL1_1X4
Xinst0x1 vss vdd wl1[0] wl2[0] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar17ArrayShWL1_1X4
.ends DP8TVar17ArrayShWL1_1X8

.subckt DP8TVar17CellConnectOut wl1 wl2 bl1 bl1_n bl2 bl2_n vdd vss bit bit_n
Xpu1 vdd bit_n bit vdd sg13_lv_pmos l=1.3e-07 w=2e-07
Xpd1 bit bit_n vss vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpu2 vdd bit bit_n vdd sg13_lv_pmos l=1.3e-07 w=2e-07
Xpd2 bit_n bit vss vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg1 bit wl1 bl1 vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg1n bit_n wl1 bl1_n vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg2 bit wl2 bl2 vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg2n bit_n wl2 bl2_n vss sg13_lv_nmos l=1.3e-07 w=2e-07
.ends DP8TVar17CellConnectOut

.subckt DP8TVar17CellShWL2 wl1 wl2 bl1 bl1_n bl2 bl2_n vdd vss
Xpu1 vdd bit_n bit vdd sg13_lv_pmos l=1.3e-07 w=2e-07
Xpd1 bit bit_n vss vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpu2 vdd bit bit_n vdd sg13_lv_pmos l=1.3e-07 w=2e-07
Xpd2 bit_n bit vss vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg1 bit wl2 bl1 vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg1n bit_n wl2 bl1_n vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg2 bit wl2 bl2 vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg2n bit_n wl2 bl2_n vss sg13_lv_nmos l=1.3e-07 w=2e-07
.ends DP8TVar17CellShWL2

.subckt DP8TVar17ArrayShWL2_1X2 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1]
Xinst0x0 wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] vdd vss DP8TVar17CellShWL2
Xinst0x1 wl1[0] wl2[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] vdd vss DP8TVar17CellShWL2
.ends DP8TVar17ArrayShWL2_1X2

.subckt DP8TVar17ArrayShWL2_1X4 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3]
Xinst0x0 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TVar17ArrayShWL2_1X2
Xinst0x1 vss vdd wl1[0] wl2[0] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar17ArrayShWL2_1X2
.ends DP8TVar17ArrayShWL2_1X4

.subckt DP8TVar17ArrayShWL2_1X8 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar17ArrayShWL2_1X4
Xinst0x1 vss vdd wl1[0] wl2[0] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar17ArrayShWL2_1X4
.ends DP8TVar17ArrayShWL2_1X8

.subckt DP8TVar17Array_6X8 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar17Array_4X8
Xinst1x0 vss vdd wl1[4] wl2[4] wl1[5] wl2[5] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar17Array_2X8
.ends DP8TVar17Array_6X8

.subckt DP8TVar17TestArray_16X8C vss vdd wl1 wl2 bl1 bl1_n bl2 bl2_n bit bit_n
Xbcconn_bot vss vdd bcconn_bot_bl1[0] bcconn_bot_bl1_n[0] bcconn_bot_bl2[0] bcconn_bot_bl2_n[0] bcconn_bot_bl1[1] bcconn_bot_bl1_n[1] bcconn_bot_bl2[1] bcconn_bot_bl2_n[1] bcconn_bot_bl1[2] bcconn_bot_bl1_n[2] bcconn_bot_bl2[2] bcconn_bot_bl2_n[2] bcconn_bot_bl1[3] bcconn_bot_bl1_n[3] bcconn_bot_bl2[3] bcconn_bot_bl2_n[3] bl1 bl1_n bl2 bl2_n bcconn_bot_bl1[5] bcconn_bot_bl1_n[5] bcconn_bot_bl2[5] bcconn_bot_bl2_n[5] bcconn_bot_bl1[6] bcconn_bot_bl1_n[6] bcconn_bot_bl2[6] bcconn_bot_bl2_n[6] bcconn_bot_bl1[7] bcconn_bot_bl1_n[7] bcconn_bot_bl2[7] bcconn_bot_bl2_n[7] DP8TVar17BulkConnRow_8
Xbcconn_top vss vdd bcconn_top_bl1[0] bcconn_top_bl1_n[0] bcconn_top_bl2[0] bcconn_top_bl2_n[0] bcconn_top_bl1[1] bcconn_top_bl1_n[1] bcconn_top_bl2[1] bcconn_top_bl2_n[1] bcconn_top_bl1[2] bcconn_top_bl1_n[2] bcconn_top_bl2[2] bcconn_top_bl2_n[2] bcconn_top_bl1[3] bcconn_top_bl1_n[3] bcconn_top_bl2[3] bcconn_top_bl2_n[3] bl1 bl1_n bl2 bl2_n bcconn_top_bl1[5] bcconn_top_bl1_n[5] bcconn_top_bl2[5] bcconn_top_bl2_n[5] bcconn_top_bl1[6] bcconn_top_bl1_n[6] bcconn_top_bl2[6] bcconn_top_bl2_n[6] bcconn_top_bl1[7] bcconn_top_bl1_n[7] bcconn_top_bl2[7] bcconn_top_bl2_n[7] DP8TVar17BulkConnRow_8
Xarray_bot vss vdd zero zero zero zero zero zero zero zero zero zero zero zero zero zero array_bot_bl1[0] array_bot_bl1_n[0] array_bot_bl2[0] array_bot_bl2_n[0] array_bot_bl1[1] array_bot_bl1_n[1] array_bot_bl2[1] array_bot_bl2_n[1] array_bot_bl1[2] array_bot_bl1_n[2] array_bot_bl2[2] array_bot_bl2_n[2] array_bot_bl1[3] array_bot_bl1_n[3] array_bot_bl2[3] array_bot_bl2_n[3] bl1 bl1_n bl2 bl2_n array_bot_bl1[5] array_bot_bl1_n[5] array_bot_bl2[5] array_bot_bl2_n[5] array_bot_bl1[6] array_bot_bl1_n[6] array_bot_bl2[6] array_bot_bl2_n[6] array_bot_bl1[7] array_bot_bl1_n[7] array_bot_bl2[7] array_bot_bl2_n[7] DP8TVar17Array_7X8
Xshwl1_row vss vdd zero bit shwl1_row_bl1[0] shwl1_row_bl1_n[0] shwl1_row_bl2[0] shwl1_row_bl2_n[0] shwl1_row_bl1[1] shwl1_row_bl1_n[1] shwl1_row_bl2[1] shwl1_row_bl2_n[1] shwl1_row_bl1[2] shwl1_row_bl1_n[2] shwl1_row_bl2[2] shwl1_row_bl2_n[2] shwl1_row_bl1[3] shwl1_row_bl1_n[3] shwl1_row_bl2[3] shwl1_row_bl2_n[3] bl1 bl1_n bl2 bl2_n shwl1_row_bl1[5] shwl1_row_bl1_n[5] shwl1_row_bl2[5] shwl1_row_bl2_n[5] shwl1_row_bl1[6] shwl1_row_bl1_n[6] shwl1_row_bl2[6] shwl1_row_bl2_n[6] shwl1_row_bl1[7] shwl1_row_bl1_n[7] shwl1_row_bl2[7] shwl1_row_bl2_n[7] DP8TVar17ArrayShWL1_1X8
Xcell_cols_left vss vdd wl1 wl2 cell_cols_left_bl1[0] cell_cols_left_bl1_n[0] cell_cols_left_bl2[0] cell_cols_left_bl2_n[0] cell_cols_left_bl1[1] cell_cols_left_bl1_n[1] cell_cols_left_bl2[1] cell_cols_left_bl2_n[1] cell_cols_left_bl1[2] cell_cols_left_bl1_n[2] cell_cols_left_bl2[2] cell_cols_left_bl2_n[2] cell_cols_left_bl1[3] cell_cols_left_bl1_n[3] cell_cols_left_bl2[3] cell_cols_left_bl2_n[3] DP8TVar17Array_1X4
Xconncell wl1 wl2 bl1 bl1_n bl2 bl2_n vdd vss bit bit_n DP8TVar17CellConnectOut
Xfillcell wl1 wl2 fillcell_bl1 fillcell_bl1_n fillcell_bl2 fillcell_bl2_n vdd vss DP8TVar17Cell
Xcell_cols_right vss vdd wl1 wl2 cell_cols_right_bl1[0] cell_cols_right_bl1_n[0] cell_cols_right_bl2[0] cell_cols_right_bl2_n[0] cell_cols_right_bl1[1] cell_cols_right_bl1_n[1] cell_cols_right_bl2[1] cell_cols_right_bl2_n[1] DP8TVar17Array_1X2
Xshwl2_row vss vdd bit_n zero shwl2_row_bl1[0] shwl2_row_bl1_n[0] shwl2_row_bl2[0] shwl2_row_bl2_n[0] shwl2_row_bl1[1] shwl2_row_bl1_n[1] shwl2_row_bl2[1] shwl2_row_bl2_n[1] shwl2_row_bl1[2] shwl2_row_bl1_n[2] shwl2_row_bl2[2] shwl2_row_bl2_n[2] shwl2_row_bl1[3] shwl2_row_bl1_n[3] shwl2_row_bl2[3] shwl2_row_bl2_n[3] bl1 bl1_n bl2 bl2_n shwl2_row_bl1[5] shwl2_row_bl1_n[5] shwl2_row_bl2[5] shwl2_row_bl2_n[5] shwl2_row_bl1[6] shwl2_row_bl1_n[6] shwl2_row_bl2[6] shwl2_row_bl2_n[6] shwl2_row_bl1[7] shwl2_row_bl1_n[7] shwl2_row_bl2[7] shwl2_row_bl2_n[7] DP8TVar17ArrayShWL2_1X8
Xarray_top vss vdd zero zero zero zero zero zero zero zero zero zero zero zero array_top_bl1[0] array_top_bl1_n[0] array_top_bl2[0] array_top_bl2_n[0] array_top_bl1[1] array_top_bl1_n[1] array_top_bl2[1] array_top_bl2_n[1] array_top_bl1[2] array_top_bl1_n[2] array_top_bl2[2] array_top_bl2_n[2] array_top_bl1[3] array_top_bl1_n[3] array_top_bl2[3] array_top_bl2_n[3] bl1 bl1_n bl2 bl2_n array_top_bl1[5] array_top_bl1_n[5] array_top_bl2[5] array_top_bl2_n[5] array_top_bl1[6] array_top_bl1_n[6] array_top_bl2[6] array_top_bl2_n[6] array_top_bl1[7] array_top_bl1_n[7] array_top_bl2[7] array_top_bl2_n[7] DP8TVar17Array_6X8
Xzero vdd vss zero zero_x1
.ends DP8TVar17TestArray_16X8C

.subckt DP8TVar17 vss noco_vdd noco_wl1 noco_wl2 noco_bl1 noco_bl1_n noco_bl2 noco_bl2_n co_vdd co_bit co_bit_n co_wl1 co_wl2 co_bl1 co_bl1_n co_bl2_n co_bl2
Xframe noco_vdd noco_wl1 noco_wl2 noco_bl2 co_vdd co_bit co_bit_n co_wl1 co_wl2 NoConn_PAD0x9 vss noco_bl1 noco_bl1_n noco_bl2_n vss co_bl1 co_bl1_n co_bl2_n co_bl2 NoConn_PAD1x9 PadFrame_DP17
Xtestarray_noco vss noco_vdd noco_wl1 noco_wl2 noco_bl1 noco_bl1_n noco_bl2 noco_bl2_n DP8TVar17TestArray_16X8
Xtestarray_co vss co_vdd co_wl1 co_wl2 co_bl1 co_bl1_n co_bl2 co_bl2_n co_bit co_bit_n DP8TVar17TestArray_16X8C
.ends DP8TVar17

.subckt PadFrame_DP18 PAD0x0 PAD0x1 PAD0x2 PAD0x3 PAD0x4 PAD0x5 PAD0x6 PAD0x7 PAD0x8 PAD0x9 PAD1x0 PAD1x1 PAD1x2 PAD1x3 PAD1x4 PAD1x5 PAD1x6 PAD1x7 PAD1x8 PAD1x9
XPAD0x0 PAD0x0 BondPad
XPAD0x1 PAD0x1 BondPad
XPAD0x2 PAD0x2 BondPad
XPAD0x3 PAD0x3 BondPad
XPAD0x4 PAD0x4 BondPad
XPAD0x5 PAD0x5 BondPad
XPAD0x6 PAD0x6 BondPad
XPAD0x7 PAD0x7 BondPad
XPAD0x8 PAD0x8 BondPad
XPAD0x9 PAD0x9 BondPad
XPAD1x0 PAD1x0 BondPad
XPAD1x1 PAD1x1 BondPad
XPAD1x2 PAD1x2 BondPad
XPAD1x3 PAD1x3 BondPad
XPAD1x4 PAD1x4 BondPad
XPAD1x5 PAD1x5 BondPad
XPAD1x6 PAD1x6 BondPad
XPAD1x7 PAD1x7 BondPad
XPAD1x8 PAD1x8 BondPad
XPAD1x9 PAD1x9 BondPad
.ends PadFrame_DP18

.subckt DP8TVar18Cell wl1 wl2 bl1 bl1_n bl2 bl2_n vdd vss
Xpu1 vdd bit_n bit vdd sg13_lv_pmos l=1.3e-07 w=1.5e-07
Xpd1 bit bit_n vss vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpu2 vdd bit bit_n vdd sg13_lv_pmos l=1.3e-07 w=1.5e-07
Xpd2 bit_n bit vss vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg1 bit wl1 bl1 vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg1n bit_n wl1 bl1_n vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg2 bit wl2 bl2 vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg2n bit_n wl2 bl2_n vss sg13_lv_nmos l=1.3e-07 w=2e-07
.ends DP8TVar18Cell

.subckt DP8TVar18Array_2X1 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0]
Xinst0x0 wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] vdd vss DP8TVar18Cell
Xinst1x0 wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0] vdd vss DP8TVar18Cell
.ends DP8TVar18Array_2X1

.subckt DP8TVar18Array_2X2 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0] DP8TVar18Array_2X1
Xinst0x1 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TVar18Array_2X1
.ends DP8TVar18Array_2X2

.subckt DP8TVar18Array_4X2 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TVar18Array_2X2
Xinst1x0 vss vdd wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TVar18Array_2X2
.ends DP8TVar18Array_4X2

.subckt DP8TVar18Array_4X4 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TVar18Array_4X2
Xinst0x1 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar18Array_4X2
.ends DP8TVar18Array_4X4

.subckt DP8TVar18Array_8X4 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar18Array_4X4
Xinst1x0 vss vdd wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar18Array_4X4
.ends DP8TVar18Array_8X4

.subckt DP8TVar18Array_8X8 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar18Array_8X4
Xinst0x1 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar18Array_8X4
.ends DP8TVar18Array_8X8

.subckt DP8TVar18BulkConn vdd vss bl1 bl2 bl1_n bl2_n
.ends DP8TVar18BulkConn

.subckt DP8TVar18BulkConnRow_2 vss vdd bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1]
Xinst0 vdd vss bl1[0] bl2[0] bl1_n[0] bl2_n[0] DP8TVar18BulkConn
Xinst1 vdd vss bl1[1] bl2[1] bl1_n[1] bl2_n[1] DP8TVar18BulkConn
.ends DP8TVar18BulkConnRow_2

.subckt DP8TVar18BulkConnRow_4 vss vdd bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3]
Xinst0 vss vdd bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TVar18BulkConnRow_2
Xinst1 vss vdd bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar18BulkConnRow_2
.ends DP8TVar18BulkConnRow_4

.subckt DP8TVar18BulkConnRow_8 vss vdd bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0 vss vdd bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar18BulkConnRow_4
Xinst1 vss vdd bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar18BulkConnRow_4
.ends DP8TVar18BulkConnRow_8

.subckt DP8TVar18Array_16X8BC vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] wl1[8] wl2[8] wl1[9] wl2[9] wl1[10] wl2[10] wl1[11] wl2[11] wl1[12] wl2[12] wl1[13] wl2[13] wl1[14] wl2[14] wl1[15] wl2[15] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar18Array_8X8
Xinst1x0 vss vdd wl1[8] wl2[8] wl1[9] wl2[9] wl1[10] wl2[10] wl1[11] wl2[11] wl1[12] wl2[12] wl1[13] wl2[13] wl1[14] wl2[14] wl1[15] wl2[15] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar18Array_8X8
Xbottombcrow vss vdd bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar18BulkConnRow_8
Xtopbcrow vss vdd bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar18BulkConnRow_8
.ends DP8TVar18Array_16X8BC

.subckt DP8TVar18TestArray_16X8 vss vdd wl1 wl2 bl1 bl1_n bl2 bl2_n
Xarray vss vdd zero zero zero zero zero zero zero zero zero zero zero zero zero zero zero zero wl1 wl2 zero zero zero zero zero zero zero zero zero zero zero zero zero zero bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1 bl1_n bl2 bl2_n bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar18Array_16X8BC
Xzero vdd vss zero zero_x1
.ends DP8TVar18TestArray_16X8

.subckt DP8TVar18Array_4X8 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar18Array_4X4
Xinst0x1 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar18Array_4X4
.ends DP8TVar18Array_4X8

.subckt DP8TVar18Array_2X4 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TVar18Array_2X2
Xinst0x1 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar18Array_2X2
.ends DP8TVar18Array_2X4

.subckt DP8TVar18Array_2X8 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar18Array_2X4
Xinst0x1 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar18Array_2X4
.ends DP8TVar18Array_2X8

.subckt DP8TVar18Array_1X2 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1]
Xinst0x0 wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] vdd vss DP8TVar18Cell
Xinst0x1 wl1[0] wl2[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] vdd vss DP8TVar18Cell
.ends DP8TVar18Array_1X2

.subckt DP8TVar18Array_1X4 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3]
Xinst0x0 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TVar18Array_1X2
Xinst0x1 vss vdd wl1[0] wl2[0] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar18Array_1X2
.ends DP8TVar18Array_1X4

.subckt DP8TVar18Array_1X8 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar18Array_1X4
Xinst0x1 vss vdd wl1[0] wl2[0] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar18Array_1X4
.ends DP8TVar18Array_1X8

.subckt DP8TVar18Array_7X8 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar18Array_4X8
Xinst1x0 vss vdd wl1[4] wl2[4] wl1[5] wl2[5] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar18Array_2X8
Xinst2x0 vss vdd wl1[6] wl2[6] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar18Array_1X8
.ends DP8TVar18Array_7X8

.subckt DP8TVar18CellShWL1 wl1 wl2 bl1 bl1_n bl2 bl2_n vdd vss
Xpu1 vdd bit_n bit vdd sg13_lv_pmos l=1.3e-07 w=1.5e-07
Xpd1 bit bit_n vss vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpu2 vdd bit bit_n vdd sg13_lv_pmos l=1.3e-07 w=1.5e-07
Xpd2 bit_n bit vss vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg1 bit wl1 bl1 vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg1n bit_n wl1 bl1_n vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg2 bit wl1 bl2 vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg2n bit_n wl1 bl2_n vss sg13_lv_nmos l=1.3e-07 w=2e-07
.ends DP8TVar18CellShWL1

.subckt DP8TVar18ArrayShWL1_1X2 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1]
Xinst0x0 wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] vdd vss DP8TVar18CellShWL1
Xinst0x1 wl1[0] wl2[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] vdd vss DP8TVar18CellShWL1
.ends DP8TVar18ArrayShWL1_1X2

.subckt DP8TVar18ArrayShWL1_1X4 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3]
Xinst0x0 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TVar18ArrayShWL1_1X2
Xinst0x1 vss vdd wl1[0] wl2[0] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar18ArrayShWL1_1X2
.ends DP8TVar18ArrayShWL1_1X4

.subckt DP8TVar18ArrayShWL1_1X8 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar18ArrayShWL1_1X4
Xinst0x1 vss vdd wl1[0] wl2[0] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar18ArrayShWL1_1X4
.ends DP8TVar18ArrayShWL1_1X8

.subckt DP8TVar18CellConnectOut wl1 wl2 bl1 bl1_n bl2 bl2_n vdd vss bit bit_n
Xpu1 vdd bit_n bit vdd sg13_lv_pmos l=1.3e-07 w=1.5e-07
Xpd1 bit bit_n vss vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpu2 vdd bit bit_n vdd sg13_lv_pmos l=1.3e-07 w=1.5e-07
Xpd2 bit_n bit vss vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg1 bit wl1 bl1 vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg1n bit_n wl1 bl1_n vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg2 bit wl2 bl2 vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg2n bit_n wl2 bl2_n vss sg13_lv_nmos l=1.3e-07 w=2e-07
.ends DP8TVar18CellConnectOut

.subckt DP8TVar18CellShWL2 wl1 wl2 bl1 bl1_n bl2 bl2_n vdd vss
Xpu1 vdd bit_n bit vdd sg13_lv_pmos l=1.3e-07 w=1.5e-07
Xpd1 bit bit_n vss vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpu2 vdd bit bit_n vdd sg13_lv_pmos l=1.3e-07 w=1.5e-07
Xpd2 bit_n bit vss vss sg13_lv_nmos l=1.3e-07 w=3e-07
Xpg1 bit wl2 bl1 vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg1n bit_n wl2 bl1_n vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg2 bit wl2 bl2 vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg2n bit_n wl2 bl2_n vss sg13_lv_nmos l=1.3e-07 w=2e-07
.ends DP8TVar18CellShWL2

.subckt DP8TVar18ArrayShWL2_1X2 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1]
Xinst0x0 wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] vdd vss DP8TVar18CellShWL2
Xinst0x1 wl1[0] wl2[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] vdd vss DP8TVar18CellShWL2
.ends DP8TVar18ArrayShWL2_1X2

.subckt DP8TVar18ArrayShWL2_1X4 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3]
Xinst0x0 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TVar18ArrayShWL2_1X2
Xinst0x1 vss vdd wl1[0] wl2[0] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar18ArrayShWL2_1X2
.ends DP8TVar18ArrayShWL2_1X4

.subckt DP8TVar18ArrayShWL2_1X8 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar18ArrayShWL2_1X4
Xinst0x1 vss vdd wl1[0] wl2[0] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar18ArrayShWL2_1X4
.ends DP8TVar18ArrayShWL2_1X8

.subckt DP8TVar18Array_6X8 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar18Array_4X8
Xinst1x0 vss vdd wl1[4] wl2[4] wl1[5] wl2[5] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar18Array_2X8
.ends DP8TVar18Array_6X8

.subckt DP8TVar18TestArray_16X8C vss vdd wl1 wl2 bl1 bl1_n bl2 bl2_n bit bit_n
Xbcconn_bot vss vdd bcconn_bot_bl1[0] bcconn_bot_bl1_n[0] bcconn_bot_bl2[0] bcconn_bot_bl2_n[0] bcconn_bot_bl1[1] bcconn_bot_bl1_n[1] bcconn_bot_bl2[1] bcconn_bot_bl2_n[1] bcconn_bot_bl1[2] bcconn_bot_bl1_n[2] bcconn_bot_bl2[2] bcconn_bot_bl2_n[2] bcconn_bot_bl1[3] bcconn_bot_bl1_n[3] bcconn_bot_bl2[3] bcconn_bot_bl2_n[3] bl1 bl1_n bl2 bl2_n bcconn_bot_bl1[5] bcconn_bot_bl1_n[5] bcconn_bot_bl2[5] bcconn_bot_bl2_n[5] bcconn_bot_bl1[6] bcconn_bot_bl1_n[6] bcconn_bot_bl2[6] bcconn_bot_bl2_n[6] bcconn_bot_bl1[7] bcconn_bot_bl1_n[7] bcconn_bot_bl2[7] bcconn_bot_bl2_n[7] DP8TVar18BulkConnRow_8
Xbcconn_top vss vdd bcconn_top_bl1[0] bcconn_top_bl1_n[0] bcconn_top_bl2[0] bcconn_top_bl2_n[0] bcconn_top_bl1[1] bcconn_top_bl1_n[1] bcconn_top_bl2[1] bcconn_top_bl2_n[1] bcconn_top_bl1[2] bcconn_top_bl1_n[2] bcconn_top_bl2[2] bcconn_top_bl2_n[2] bcconn_top_bl1[3] bcconn_top_bl1_n[3] bcconn_top_bl2[3] bcconn_top_bl2_n[3] bl1 bl1_n bl2 bl2_n bcconn_top_bl1[5] bcconn_top_bl1_n[5] bcconn_top_bl2[5] bcconn_top_bl2_n[5] bcconn_top_bl1[6] bcconn_top_bl1_n[6] bcconn_top_bl2[6] bcconn_top_bl2_n[6] bcconn_top_bl1[7] bcconn_top_bl1_n[7] bcconn_top_bl2[7] bcconn_top_bl2_n[7] DP8TVar18BulkConnRow_8
Xarray_bot vss vdd zero zero zero zero zero zero zero zero zero zero zero zero zero zero array_bot_bl1[0] array_bot_bl1_n[0] array_bot_bl2[0] array_bot_bl2_n[0] array_bot_bl1[1] array_bot_bl1_n[1] array_bot_bl2[1] array_bot_bl2_n[1] array_bot_bl1[2] array_bot_bl1_n[2] array_bot_bl2[2] array_bot_bl2_n[2] array_bot_bl1[3] array_bot_bl1_n[3] array_bot_bl2[3] array_bot_bl2_n[3] bl1 bl1_n bl2 bl2_n array_bot_bl1[5] array_bot_bl1_n[5] array_bot_bl2[5] array_bot_bl2_n[5] array_bot_bl1[6] array_bot_bl1_n[6] array_bot_bl2[6] array_bot_bl2_n[6] array_bot_bl1[7] array_bot_bl1_n[7] array_bot_bl2[7] array_bot_bl2_n[7] DP8TVar18Array_7X8
Xshwl1_row vss vdd zero bit shwl1_row_bl1[0] shwl1_row_bl1_n[0] shwl1_row_bl2[0] shwl1_row_bl2_n[0] shwl1_row_bl1[1] shwl1_row_bl1_n[1] shwl1_row_bl2[1] shwl1_row_bl2_n[1] shwl1_row_bl1[2] shwl1_row_bl1_n[2] shwl1_row_bl2[2] shwl1_row_bl2_n[2] shwl1_row_bl1[3] shwl1_row_bl1_n[3] shwl1_row_bl2[3] shwl1_row_bl2_n[3] bl1 bl1_n bl2 bl2_n shwl1_row_bl1[5] shwl1_row_bl1_n[5] shwl1_row_bl2[5] shwl1_row_bl2_n[5] shwl1_row_bl1[6] shwl1_row_bl1_n[6] shwl1_row_bl2[6] shwl1_row_bl2_n[6] shwl1_row_bl1[7] shwl1_row_bl1_n[7] shwl1_row_bl2[7] shwl1_row_bl2_n[7] DP8TVar18ArrayShWL1_1X8
Xcell_cols_left vss vdd wl1 wl2 cell_cols_left_bl1[0] cell_cols_left_bl1_n[0] cell_cols_left_bl2[0] cell_cols_left_bl2_n[0] cell_cols_left_bl1[1] cell_cols_left_bl1_n[1] cell_cols_left_bl2[1] cell_cols_left_bl2_n[1] cell_cols_left_bl1[2] cell_cols_left_bl1_n[2] cell_cols_left_bl2[2] cell_cols_left_bl2_n[2] cell_cols_left_bl1[3] cell_cols_left_bl1_n[3] cell_cols_left_bl2[3] cell_cols_left_bl2_n[3] DP8TVar18Array_1X4
Xconncell wl1 wl2 bl1 bl1_n bl2 bl2_n vdd vss bit bit_n DP8TVar18CellConnectOut
Xfillcell wl1 wl2 fillcell_bl1 fillcell_bl1_n fillcell_bl2 fillcell_bl2_n vdd vss DP8TVar18Cell
Xcell_cols_right vss vdd wl1 wl2 cell_cols_right_bl1[0] cell_cols_right_bl1_n[0] cell_cols_right_bl2[0] cell_cols_right_bl2_n[0] cell_cols_right_bl1[1] cell_cols_right_bl1_n[1] cell_cols_right_bl2[1] cell_cols_right_bl2_n[1] DP8TVar18Array_1X2
Xshwl2_row vss vdd bit_n zero shwl2_row_bl1[0] shwl2_row_bl1_n[0] shwl2_row_bl2[0] shwl2_row_bl2_n[0] shwl2_row_bl1[1] shwl2_row_bl1_n[1] shwl2_row_bl2[1] shwl2_row_bl2_n[1] shwl2_row_bl1[2] shwl2_row_bl1_n[2] shwl2_row_bl2[2] shwl2_row_bl2_n[2] shwl2_row_bl1[3] shwl2_row_bl1_n[3] shwl2_row_bl2[3] shwl2_row_bl2_n[3] bl1 bl1_n bl2 bl2_n shwl2_row_bl1[5] shwl2_row_bl1_n[5] shwl2_row_bl2[5] shwl2_row_bl2_n[5] shwl2_row_bl1[6] shwl2_row_bl1_n[6] shwl2_row_bl2[6] shwl2_row_bl2_n[6] shwl2_row_bl1[7] shwl2_row_bl1_n[7] shwl2_row_bl2[7] shwl2_row_bl2_n[7] DP8TVar18ArrayShWL2_1X8
Xarray_top vss vdd zero zero zero zero zero zero zero zero zero zero zero zero array_top_bl1[0] array_top_bl1_n[0] array_top_bl2[0] array_top_bl2_n[0] array_top_bl1[1] array_top_bl1_n[1] array_top_bl2[1] array_top_bl2_n[1] array_top_bl1[2] array_top_bl1_n[2] array_top_bl2[2] array_top_bl2_n[2] array_top_bl1[3] array_top_bl1_n[3] array_top_bl2[3] array_top_bl2_n[3] bl1 bl1_n bl2 bl2_n array_top_bl1[5] array_top_bl1_n[5] array_top_bl2[5] array_top_bl2_n[5] array_top_bl1[6] array_top_bl1_n[6] array_top_bl2[6] array_top_bl2_n[6] array_top_bl1[7] array_top_bl1_n[7] array_top_bl2[7] array_top_bl2_n[7] DP8TVar18Array_6X8
Xzero vdd vss zero zero_x1
.ends DP8TVar18TestArray_16X8C

.subckt DP8TVar18 vss noco_vdd noco_wl1 noco_wl2 noco_bl1 noco_bl1_n noco_bl2 noco_bl2_n co_vdd co_bit co_bit_n co_wl1 co_wl2 co_bl1 co_bl1_n co_bl2_n co_bl2
Xframe noco_vdd noco_wl1 noco_wl2 noco_bl2 co_vdd co_bit co_bit_n co_wl1 co_wl2 NoConn_PAD0x9 vss noco_bl1 noco_bl1_n noco_bl2_n vss co_bl1 co_bl1_n co_bl2_n co_bl2 NoConn_PAD1x9 PadFrame_DP18
Xtestarray_noco vss noco_vdd noco_wl1 noco_wl2 noco_bl1 noco_bl1_n noco_bl2 noco_bl2_n DP8TVar18TestArray_16X8
Xtestarray_co vss co_vdd co_wl1 co_wl2 co_bl1 co_bl1_n co_bl2 co_bl2_n co_bit co_bit_n DP8TVar18TestArray_16X8C
.ends DP8TVar18

.subckt PadFrame_DP19 PAD0x0 PAD0x1 PAD0x2 PAD0x3 PAD0x4 PAD0x5 PAD0x6 PAD0x7 PAD0x8 PAD0x9 PAD1x0 PAD1x1 PAD1x2 PAD1x3 PAD1x4 PAD1x5 PAD1x6 PAD1x7 PAD1x8 PAD1x9
XPAD0x0 PAD0x0 BondPad
XPAD0x1 PAD0x1 BondPad
XPAD0x2 PAD0x2 BondPad
XPAD0x3 PAD0x3 BondPad
XPAD0x4 PAD0x4 BondPad
XPAD0x5 PAD0x5 BondPad
XPAD0x6 PAD0x6 BondPad
XPAD0x7 PAD0x7 BondPad
XPAD0x8 PAD0x8 BondPad
XPAD0x9 PAD0x9 BondPad
XPAD1x0 PAD1x0 BondPad
XPAD1x1 PAD1x1 BondPad
XPAD1x2 PAD1x2 BondPad
XPAD1x3 PAD1x3 BondPad
XPAD1x4 PAD1x4 BondPad
XPAD1x5 PAD1x5 BondPad
XPAD1x6 PAD1x6 BondPad
XPAD1x7 PAD1x7 BondPad
XPAD1x8 PAD1x8 BondPad
XPAD1x9 PAD1x9 BondPad
.ends PadFrame_DP19

.subckt DP8TVar19Cell wl1 wl2 bl1 bl1_n bl2 bl2_n vdd vss
Xpu1 vdd bit_n bit vdd sg13_lv_pmos l=1.3e-07 w=2e-07
Xpd1 bit bit_n vss vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpu2 vdd bit bit_n vdd sg13_lv_pmos l=1.3e-07 w=2e-07
Xpd2 bit_n bit vss vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg1 bit wl1 bl1 vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg1n bit_n wl1 bl1_n vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg2 bit wl2 bl2 vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg2n bit_n wl2 bl2_n vss sg13_lv_nmos l=1.3e-07 w=2e-07
.ends DP8TVar19Cell

.subckt DP8TVar19Array_2X1 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0]
Xinst0x0 wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] vdd vss DP8TVar19Cell
Xinst1x0 wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0] vdd vss DP8TVar19Cell
.ends DP8TVar19Array_2X1

.subckt DP8TVar19Array_2X2 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0] DP8TVar19Array_2X1
Xinst0x1 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TVar19Array_2X1
.ends DP8TVar19Array_2X2

.subckt DP8TVar19Array_4X2 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TVar19Array_2X2
Xinst1x0 vss vdd wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TVar19Array_2X2
.ends DP8TVar19Array_4X2

.subckt DP8TVar19Array_4X4 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TVar19Array_4X2
Xinst0x1 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar19Array_4X2
.ends DP8TVar19Array_4X4

.subckt DP8TVar19Array_8X4 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar19Array_4X4
Xinst1x0 vss vdd wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar19Array_4X4
.ends DP8TVar19Array_8X4

.subckt DP8TVar19Array_8X8 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar19Array_8X4
Xinst0x1 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar19Array_8X4
.ends DP8TVar19Array_8X8

.subckt DP8TVar19BulkConn vdd vss bl1 bl2 bl1_n bl2_n
.ends DP8TVar19BulkConn

.subckt DP8TVar19BulkConnRow_2 vss vdd bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1]
Xinst0 vdd vss bl1[0] bl2[0] bl1_n[0] bl2_n[0] DP8TVar19BulkConn
Xinst1 vdd vss bl1[1] bl2[1] bl1_n[1] bl2_n[1] DP8TVar19BulkConn
.ends DP8TVar19BulkConnRow_2

.subckt DP8TVar19BulkConnRow_4 vss vdd bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3]
Xinst0 vss vdd bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TVar19BulkConnRow_2
Xinst1 vss vdd bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar19BulkConnRow_2
.ends DP8TVar19BulkConnRow_4

.subckt DP8TVar19BulkConnRow_8 vss vdd bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0 vss vdd bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar19BulkConnRow_4
Xinst1 vss vdd bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar19BulkConnRow_4
.ends DP8TVar19BulkConnRow_8

.subckt DP8TVar19Array_16X8BC vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] wl1[8] wl2[8] wl1[9] wl2[9] wl1[10] wl2[10] wl1[11] wl2[11] wl1[12] wl2[12] wl1[13] wl2[13] wl1[14] wl2[14] wl1[15] wl2[15] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar19Array_8X8
Xinst1x0 vss vdd wl1[8] wl2[8] wl1[9] wl2[9] wl1[10] wl2[10] wl1[11] wl2[11] wl1[12] wl2[12] wl1[13] wl2[13] wl1[14] wl2[14] wl1[15] wl2[15] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar19Array_8X8
Xbottombcrow vss vdd bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar19BulkConnRow_8
Xtopbcrow vss vdd bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar19BulkConnRow_8
.ends DP8TVar19Array_16X8BC

.subckt DP8TVar19TestArray_16X8 vss vdd wl1 wl2 bl1 bl1_n bl2 bl2_n
Xarray vss vdd zero zero zero zero zero zero zero zero zero zero zero zero zero zero zero zero wl1 wl2 zero zero zero zero zero zero zero zero zero zero zero zero zero zero bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1 bl1_n bl2 bl2_n bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar19Array_16X8BC
Xzero vdd vss zero zero_x1
.ends DP8TVar19TestArray_16X8

.subckt DP8TVar19Array_4X8 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar19Array_4X4
Xinst0x1 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar19Array_4X4
.ends DP8TVar19Array_4X8

.subckt DP8TVar19Array_2X4 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TVar19Array_2X2
Xinst0x1 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar19Array_2X2
.ends DP8TVar19Array_2X4

.subckt DP8TVar19Array_2X8 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar19Array_2X4
Xinst0x1 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar19Array_2X4
.ends DP8TVar19Array_2X8

.subckt DP8TVar19Array_1X2 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1]
Xinst0x0 wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] vdd vss DP8TVar19Cell
Xinst0x1 wl1[0] wl2[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] vdd vss DP8TVar19Cell
.ends DP8TVar19Array_1X2

.subckt DP8TVar19Array_1X4 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3]
Xinst0x0 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TVar19Array_1X2
Xinst0x1 vss vdd wl1[0] wl2[0] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar19Array_1X2
.ends DP8TVar19Array_1X4

.subckt DP8TVar19Array_1X8 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar19Array_1X4
Xinst0x1 vss vdd wl1[0] wl2[0] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar19Array_1X4
.ends DP8TVar19Array_1X8

.subckt DP8TVar19Array_7X8 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar19Array_4X8
Xinst1x0 vss vdd wl1[4] wl2[4] wl1[5] wl2[5] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar19Array_2X8
Xinst2x0 vss vdd wl1[6] wl2[6] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar19Array_1X8
.ends DP8TVar19Array_7X8

.subckt DP8TVar19CellShWL1 wl1 wl2 bl1 bl1_n bl2 bl2_n vdd vss
Xpu1 vdd bit_n bit vdd sg13_lv_pmos l=1.3e-07 w=2e-07
Xpd1 bit bit_n vss vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpu2 vdd bit bit_n vdd sg13_lv_pmos l=1.3e-07 w=2e-07
Xpd2 bit_n bit vss vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg1 bit wl1 bl1 vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg1n bit_n wl1 bl1_n vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg2 bit wl1 bl2 vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg2n bit_n wl1 bl2_n vss sg13_lv_nmos l=1.3e-07 w=2e-07
.ends DP8TVar19CellShWL1

.subckt DP8TVar19ArrayShWL1_1X2 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1]
Xinst0x0 wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] vdd vss DP8TVar19CellShWL1
Xinst0x1 wl1[0] wl2[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] vdd vss DP8TVar19CellShWL1
.ends DP8TVar19ArrayShWL1_1X2

.subckt DP8TVar19ArrayShWL1_1X4 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3]
Xinst0x0 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TVar19ArrayShWL1_1X2
Xinst0x1 vss vdd wl1[0] wl2[0] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar19ArrayShWL1_1X2
.ends DP8TVar19ArrayShWL1_1X4

.subckt DP8TVar19ArrayShWL1_1X8 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar19ArrayShWL1_1X4
Xinst0x1 vss vdd wl1[0] wl2[0] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar19ArrayShWL1_1X4
.ends DP8TVar19ArrayShWL1_1X8

.subckt DP8TVar19CellConnectOut wl1 wl2 bl1 bl1_n bl2 bl2_n vdd vss bit bit_n
Xpu1 vdd bit_n bit vdd sg13_lv_pmos l=1.3e-07 w=2e-07
Xpd1 bit bit_n vss vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpu2 vdd bit bit_n vdd sg13_lv_pmos l=1.3e-07 w=2e-07
Xpd2 bit_n bit vss vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg1 bit wl1 bl1 vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg1n bit_n wl1 bl1_n vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg2 bit wl2 bl2 vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg2n bit_n wl2 bl2_n vss sg13_lv_nmos l=1.3e-07 w=2e-07
.ends DP8TVar19CellConnectOut

.subckt DP8TVar19CellShWL2 wl1 wl2 bl1 bl1_n bl2 bl2_n vdd vss
Xpu1 vdd bit_n bit vdd sg13_lv_pmos l=1.3e-07 w=2e-07
Xpd1 bit bit_n vss vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpu2 vdd bit bit_n vdd sg13_lv_pmos l=1.3e-07 w=2e-07
Xpd2 bit_n bit vss vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg1 bit wl2 bl1 vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg1n bit_n wl2 bl1_n vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg2 bit wl2 bl2 vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg2n bit_n wl2 bl2_n vss sg13_lv_nmos l=1.3e-07 w=2e-07
.ends DP8TVar19CellShWL2

.subckt DP8TVar19ArrayShWL2_1X2 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1]
Xinst0x0 wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] vdd vss DP8TVar19CellShWL2
Xinst0x1 wl1[0] wl2[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] vdd vss DP8TVar19CellShWL2
.ends DP8TVar19ArrayShWL2_1X2

.subckt DP8TVar19ArrayShWL2_1X4 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3]
Xinst0x0 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TVar19ArrayShWL2_1X2
Xinst0x1 vss vdd wl1[0] wl2[0] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar19ArrayShWL2_1X2
.ends DP8TVar19ArrayShWL2_1X4

.subckt DP8TVar19ArrayShWL2_1X8 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar19ArrayShWL2_1X4
Xinst0x1 vss vdd wl1[0] wl2[0] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar19ArrayShWL2_1X4
.ends DP8TVar19ArrayShWL2_1X8

.subckt DP8TVar19Array_6X8 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar19Array_4X8
Xinst1x0 vss vdd wl1[4] wl2[4] wl1[5] wl2[5] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar19Array_2X8
.ends DP8TVar19Array_6X8

.subckt DP8TVar19TestArray_16X8C vss vdd wl1 wl2 bl1 bl1_n bl2 bl2_n bit bit_n
Xbcconn_bot vss vdd bcconn_bot_bl1[0] bcconn_bot_bl1_n[0] bcconn_bot_bl2[0] bcconn_bot_bl2_n[0] bcconn_bot_bl1[1] bcconn_bot_bl1_n[1] bcconn_bot_bl2[1] bcconn_bot_bl2_n[1] bcconn_bot_bl1[2] bcconn_bot_bl1_n[2] bcconn_bot_bl2[2] bcconn_bot_bl2_n[2] bcconn_bot_bl1[3] bcconn_bot_bl1_n[3] bcconn_bot_bl2[3] bcconn_bot_bl2_n[3] bl1 bl1_n bl2 bl2_n bcconn_bot_bl1[5] bcconn_bot_bl1_n[5] bcconn_bot_bl2[5] bcconn_bot_bl2_n[5] bcconn_bot_bl1[6] bcconn_bot_bl1_n[6] bcconn_bot_bl2[6] bcconn_bot_bl2_n[6] bcconn_bot_bl1[7] bcconn_bot_bl1_n[7] bcconn_bot_bl2[7] bcconn_bot_bl2_n[7] DP8TVar19BulkConnRow_8
Xbcconn_top vss vdd bcconn_top_bl1[0] bcconn_top_bl1_n[0] bcconn_top_bl2[0] bcconn_top_bl2_n[0] bcconn_top_bl1[1] bcconn_top_bl1_n[1] bcconn_top_bl2[1] bcconn_top_bl2_n[1] bcconn_top_bl1[2] bcconn_top_bl1_n[2] bcconn_top_bl2[2] bcconn_top_bl2_n[2] bcconn_top_bl1[3] bcconn_top_bl1_n[3] bcconn_top_bl2[3] bcconn_top_bl2_n[3] bl1 bl1_n bl2 bl2_n bcconn_top_bl1[5] bcconn_top_bl1_n[5] bcconn_top_bl2[5] bcconn_top_bl2_n[5] bcconn_top_bl1[6] bcconn_top_bl1_n[6] bcconn_top_bl2[6] bcconn_top_bl2_n[6] bcconn_top_bl1[7] bcconn_top_bl1_n[7] bcconn_top_bl2[7] bcconn_top_bl2_n[7] DP8TVar19BulkConnRow_8
Xarray_bot vss vdd zero zero zero zero zero zero zero zero zero zero zero zero zero zero array_bot_bl1[0] array_bot_bl1_n[0] array_bot_bl2[0] array_bot_bl2_n[0] array_bot_bl1[1] array_bot_bl1_n[1] array_bot_bl2[1] array_bot_bl2_n[1] array_bot_bl1[2] array_bot_bl1_n[2] array_bot_bl2[2] array_bot_bl2_n[2] array_bot_bl1[3] array_bot_bl1_n[3] array_bot_bl2[3] array_bot_bl2_n[3] bl1 bl1_n bl2 bl2_n array_bot_bl1[5] array_bot_bl1_n[5] array_bot_bl2[5] array_bot_bl2_n[5] array_bot_bl1[6] array_bot_bl1_n[6] array_bot_bl2[6] array_bot_bl2_n[6] array_bot_bl1[7] array_bot_bl1_n[7] array_bot_bl2[7] array_bot_bl2_n[7] DP8TVar19Array_7X8
Xshwl1_row vss vdd zero bit shwl1_row_bl1[0] shwl1_row_bl1_n[0] shwl1_row_bl2[0] shwl1_row_bl2_n[0] shwl1_row_bl1[1] shwl1_row_bl1_n[1] shwl1_row_bl2[1] shwl1_row_bl2_n[1] shwl1_row_bl1[2] shwl1_row_bl1_n[2] shwl1_row_bl2[2] shwl1_row_bl2_n[2] shwl1_row_bl1[3] shwl1_row_bl1_n[3] shwl1_row_bl2[3] shwl1_row_bl2_n[3] bl1 bl1_n bl2 bl2_n shwl1_row_bl1[5] shwl1_row_bl1_n[5] shwl1_row_bl2[5] shwl1_row_bl2_n[5] shwl1_row_bl1[6] shwl1_row_bl1_n[6] shwl1_row_bl2[6] shwl1_row_bl2_n[6] shwl1_row_bl1[7] shwl1_row_bl1_n[7] shwl1_row_bl2[7] shwl1_row_bl2_n[7] DP8TVar19ArrayShWL1_1X8
Xcell_cols_left vss vdd wl1 wl2 cell_cols_left_bl1[0] cell_cols_left_bl1_n[0] cell_cols_left_bl2[0] cell_cols_left_bl2_n[0] cell_cols_left_bl1[1] cell_cols_left_bl1_n[1] cell_cols_left_bl2[1] cell_cols_left_bl2_n[1] cell_cols_left_bl1[2] cell_cols_left_bl1_n[2] cell_cols_left_bl2[2] cell_cols_left_bl2_n[2] cell_cols_left_bl1[3] cell_cols_left_bl1_n[3] cell_cols_left_bl2[3] cell_cols_left_bl2_n[3] DP8TVar19Array_1X4
Xconncell wl1 wl2 bl1 bl1_n bl2 bl2_n vdd vss bit bit_n DP8TVar19CellConnectOut
Xfillcell wl1 wl2 fillcell_bl1 fillcell_bl1_n fillcell_bl2 fillcell_bl2_n vdd vss DP8TVar19Cell
Xcell_cols_right vss vdd wl1 wl2 cell_cols_right_bl1[0] cell_cols_right_bl1_n[0] cell_cols_right_bl2[0] cell_cols_right_bl2_n[0] cell_cols_right_bl1[1] cell_cols_right_bl1_n[1] cell_cols_right_bl2[1] cell_cols_right_bl2_n[1] DP8TVar19Array_1X2
Xshwl2_row vss vdd bit_n zero shwl2_row_bl1[0] shwl2_row_bl1_n[0] shwl2_row_bl2[0] shwl2_row_bl2_n[0] shwl2_row_bl1[1] shwl2_row_bl1_n[1] shwl2_row_bl2[1] shwl2_row_bl2_n[1] shwl2_row_bl1[2] shwl2_row_bl1_n[2] shwl2_row_bl2[2] shwl2_row_bl2_n[2] shwl2_row_bl1[3] shwl2_row_bl1_n[3] shwl2_row_bl2[3] shwl2_row_bl2_n[3] bl1 bl1_n bl2 bl2_n shwl2_row_bl1[5] shwl2_row_bl1_n[5] shwl2_row_bl2[5] shwl2_row_bl2_n[5] shwl2_row_bl1[6] shwl2_row_bl1_n[6] shwl2_row_bl2[6] shwl2_row_bl2_n[6] shwl2_row_bl1[7] shwl2_row_bl1_n[7] shwl2_row_bl2[7] shwl2_row_bl2_n[7] DP8TVar19ArrayShWL2_1X8
Xarray_top vss vdd zero zero zero zero zero zero zero zero zero zero zero zero array_top_bl1[0] array_top_bl1_n[0] array_top_bl2[0] array_top_bl2_n[0] array_top_bl1[1] array_top_bl1_n[1] array_top_bl2[1] array_top_bl2_n[1] array_top_bl1[2] array_top_bl1_n[2] array_top_bl2[2] array_top_bl2_n[2] array_top_bl1[3] array_top_bl1_n[3] array_top_bl2[3] array_top_bl2_n[3] bl1 bl1_n bl2 bl2_n array_top_bl1[5] array_top_bl1_n[5] array_top_bl2[5] array_top_bl2_n[5] array_top_bl1[6] array_top_bl1_n[6] array_top_bl2[6] array_top_bl2_n[6] array_top_bl1[7] array_top_bl1_n[7] array_top_bl2[7] array_top_bl2_n[7] DP8TVar19Array_6X8
Xzero vdd vss zero zero_x1
.ends DP8TVar19TestArray_16X8C

.subckt DP8TVar19 vss noco_vdd noco_wl1 noco_wl2 noco_bl1 noco_bl1_n noco_bl2 noco_bl2_n co_vdd co_bit co_bit_n co_wl1 co_wl2 co_bl1 co_bl1_n co_bl2_n co_bl2
Xframe noco_vdd noco_wl1 noco_wl2 noco_bl2 co_vdd co_bit co_bit_n co_wl1 co_wl2 NoConn_PAD0x9 vss noco_bl1 noco_bl1_n noco_bl2_n vss co_bl1 co_bl1_n co_bl2_n co_bl2 NoConn_PAD1x9 PadFrame_DP19
Xtestarray_noco vss noco_vdd noco_wl1 noco_wl2 noco_bl1 noco_bl1_n noco_bl2 noco_bl2_n DP8TVar19TestArray_16X8
Xtestarray_co vss co_vdd co_wl1 co_wl2 co_bl1 co_bl1_n co_bl2 co_bl2_n co_bit co_bit_n DP8TVar19TestArray_16X8C
.ends DP8TVar19

.subckt PadFrame_DP20 PAD0x0 PAD0x1 PAD0x2 PAD0x3 PAD0x4 PAD0x5 PAD0x6 PAD0x7 PAD0x8 PAD0x9 PAD1x0 PAD1x1 PAD1x2 PAD1x3 PAD1x4 PAD1x5 PAD1x6 PAD1x7 PAD1x8 PAD1x9
XPAD0x0 PAD0x0 BondPad
XPAD0x1 PAD0x1 BondPad
XPAD0x2 PAD0x2 BondPad
XPAD0x3 PAD0x3 BondPad
XPAD0x4 PAD0x4 BondPad
XPAD0x5 PAD0x5 BondPad
XPAD0x6 PAD0x6 BondPad
XPAD0x7 PAD0x7 BondPad
XPAD0x8 PAD0x8 BondPad
XPAD0x9 PAD0x9 BondPad
XPAD1x0 PAD1x0 BondPad
XPAD1x1 PAD1x1 BondPad
XPAD1x2 PAD1x2 BondPad
XPAD1x3 PAD1x3 BondPad
XPAD1x4 PAD1x4 BondPad
XPAD1x5 PAD1x5 BondPad
XPAD1x6 PAD1x6 BondPad
XPAD1x7 PAD1x7 BondPad
XPAD1x8 PAD1x8 BondPad
XPAD1x9 PAD1x9 BondPad
.ends PadFrame_DP20

.subckt DP8TVar20Cell wl1 wl2 bl1 bl1_n bl2 bl2_n vdd vss
Xpu1 vdd bit_n bit vdd sg13_lv_pmos l=1.3e-07 w=1.5e-07
Xpd1 bit bit_n vss vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpu2 vdd bit bit_n vdd sg13_lv_pmos l=1.3e-07 w=1.5e-07
Xpd2 bit_n bit vss vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg1 bit wl1 bl1 vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg1n bit_n wl1 bl1_n vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg2 bit wl2 bl2 vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg2n bit_n wl2 bl2_n vss sg13_lv_nmos l=1.3e-07 w=2e-07
.ends DP8TVar20Cell

.subckt DP8TVar20Array_2X1 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0]
Xinst0x0 wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] vdd vss DP8TVar20Cell
Xinst1x0 wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0] vdd vss DP8TVar20Cell
.ends DP8TVar20Array_2X1

.subckt DP8TVar20Array_2X2 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0] DP8TVar20Array_2X1
Xinst0x1 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TVar20Array_2X1
.ends DP8TVar20Array_2X2

.subckt DP8TVar20Array_4X2 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TVar20Array_2X2
Xinst1x0 vss vdd wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TVar20Array_2X2
.ends DP8TVar20Array_4X2

.subckt DP8TVar20Array_4X4 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TVar20Array_4X2
Xinst0x1 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar20Array_4X2
.ends DP8TVar20Array_4X4

.subckt DP8TVar20Array_8X4 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar20Array_4X4
Xinst1x0 vss vdd wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar20Array_4X4
.ends DP8TVar20Array_8X4

.subckt DP8TVar20Array_8X8 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar20Array_8X4
Xinst0x1 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar20Array_8X4
.ends DP8TVar20Array_8X8

.subckt DP8TVar20BulkConn vdd vss bl1 bl2 bl1_n bl2_n
.ends DP8TVar20BulkConn

.subckt DP8TVar20BulkConnRow_2 vss vdd bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1]
Xinst0 vdd vss bl1[0] bl2[0] bl1_n[0] bl2_n[0] DP8TVar20BulkConn
Xinst1 vdd vss bl1[1] bl2[1] bl1_n[1] bl2_n[1] DP8TVar20BulkConn
.ends DP8TVar20BulkConnRow_2

.subckt DP8TVar20BulkConnRow_4 vss vdd bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3]
Xinst0 vss vdd bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TVar20BulkConnRow_2
Xinst1 vss vdd bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar20BulkConnRow_2
.ends DP8TVar20BulkConnRow_4

.subckt DP8TVar20BulkConnRow_8 vss vdd bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0 vss vdd bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar20BulkConnRow_4
Xinst1 vss vdd bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar20BulkConnRow_4
.ends DP8TVar20BulkConnRow_8

.subckt DP8TVar20Array_16X8BC vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] wl1[8] wl2[8] wl1[9] wl2[9] wl1[10] wl2[10] wl1[11] wl2[11] wl1[12] wl2[12] wl1[13] wl2[13] wl1[14] wl2[14] wl1[15] wl2[15] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar20Array_8X8
Xinst1x0 vss vdd wl1[8] wl2[8] wl1[9] wl2[9] wl1[10] wl2[10] wl1[11] wl2[11] wl1[12] wl2[12] wl1[13] wl2[13] wl1[14] wl2[14] wl1[15] wl2[15] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar20Array_8X8
Xbottombcrow vss vdd bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar20BulkConnRow_8
Xtopbcrow vss vdd bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar20BulkConnRow_8
.ends DP8TVar20Array_16X8BC

.subckt DP8TVar20TestArray_16X8 vss vdd wl1 wl2 bl1 bl1_n bl2 bl2_n
Xarray vss vdd zero zero zero zero zero zero zero zero zero zero zero zero zero zero zero zero wl1 wl2 zero zero zero zero zero zero zero zero zero zero zero zero zero zero bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1 bl1_n bl2 bl2_n bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar20Array_16X8BC
Xzero vdd vss zero zero_x1
.ends DP8TVar20TestArray_16X8

.subckt DP8TVar20Array_4X8 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar20Array_4X4
Xinst0x1 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar20Array_4X4
.ends DP8TVar20Array_4X8

.subckt DP8TVar20Array_2X4 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TVar20Array_2X2
Xinst0x1 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar20Array_2X2
.ends DP8TVar20Array_2X4

.subckt DP8TVar20Array_2X8 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar20Array_2X4
Xinst0x1 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar20Array_2X4
.ends DP8TVar20Array_2X8

.subckt DP8TVar20Array_1X2 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1]
Xinst0x0 wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] vdd vss DP8TVar20Cell
Xinst0x1 wl1[0] wl2[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] vdd vss DP8TVar20Cell
.ends DP8TVar20Array_1X2

.subckt DP8TVar20Array_1X4 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3]
Xinst0x0 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TVar20Array_1X2
Xinst0x1 vss vdd wl1[0] wl2[0] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar20Array_1X2
.ends DP8TVar20Array_1X4

.subckt DP8TVar20Array_1X8 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar20Array_1X4
Xinst0x1 vss vdd wl1[0] wl2[0] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar20Array_1X4
.ends DP8TVar20Array_1X8

.subckt DP8TVar20Array_7X8 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar20Array_4X8
Xinst1x0 vss vdd wl1[4] wl2[4] wl1[5] wl2[5] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar20Array_2X8
Xinst2x0 vss vdd wl1[6] wl2[6] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar20Array_1X8
.ends DP8TVar20Array_7X8

.subckt DP8TVar20CellShWL1 wl1 wl2 bl1 bl1_n bl2 bl2_n vdd vss
Xpu1 vdd bit_n bit vdd sg13_lv_pmos l=1.3e-07 w=1.5e-07
Xpd1 bit bit_n vss vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpu2 vdd bit bit_n vdd sg13_lv_pmos l=1.3e-07 w=1.5e-07
Xpd2 bit_n bit vss vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg1 bit wl1 bl1 vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg1n bit_n wl1 bl1_n vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg2 bit wl1 bl2 vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg2n bit_n wl1 bl2_n vss sg13_lv_nmos l=1.3e-07 w=2e-07
.ends DP8TVar20CellShWL1

.subckt DP8TVar20ArrayShWL1_1X2 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1]
Xinst0x0 wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] vdd vss DP8TVar20CellShWL1
Xinst0x1 wl1[0] wl2[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] vdd vss DP8TVar20CellShWL1
.ends DP8TVar20ArrayShWL1_1X2

.subckt DP8TVar20ArrayShWL1_1X4 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3]
Xinst0x0 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TVar20ArrayShWL1_1X2
Xinst0x1 vss vdd wl1[0] wl2[0] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar20ArrayShWL1_1X2
.ends DP8TVar20ArrayShWL1_1X4

.subckt DP8TVar20ArrayShWL1_1X8 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar20ArrayShWL1_1X4
Xinst0x1 vss vdd wl1[0] wl2[0] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar20ArrayShWL1_1X4
.ends DP8TVar20ArrayShWL1_1X8

.subckt DP8TVar20CellConnectOut wl1 wl2 bl1 bl1_n bl2 bl2_n vdd vss bit bit_n
Xpu1 vdd bit_n bit vdd sg13_lv_pmos l=1.3e-07 w=1.5e-07
Xpd1 bit bit_n vss vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpu2 vdd bit bit_n vdd sg13_lv_pmos l=1.3e-07 w=1.5e-07
Xpd2 bit_n bit vss vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg1 bit wl1 bl1 vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg1n bit_n wl1 bl1_n vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg2 bit wl2 bl2 vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg2n bit_n wl2 bl2_n vss sg13_lv_nmos l=1.3e-07 w=2e-07
.ends DP8TVar20CellConnectOut

.subckt DP8TVar20CellShWL2 wl1 wl2 bl1 bl1_n bl2 bl2_n vdd vss
Xpu1 vdd bit_n bit vdd sg13_lv_pmos l=1.3e-07 w=1.5e-07
Xpd1 bit bit_n vss vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpu2 vdd bit bit_n vdd sg13_lv_pmos l=1.3e-07 w=1.5e-07
Xpd2 bit_n bit vss vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg1 bit wl2 bl1 vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg1n bit_n wl2 bl1_n vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg2 bit wl2 bl2 vss sg13_lv_nmos l=1.3e-07 w=2e-07
Xpg2n bit_n wl2 bl2_n vss sg13_lv_nmos l=1.3e-07 w=2e-07
.ends DP8TVar20CellShWL2

.subckt DP8TVar20ArrayShWL2_1X2 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1]
Xinst0x0 wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] vdd vss DP8TVar20CellShWL2
Xinst0x1 wl1[0] wl2[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] vdd vss DP8TVar20CellShWL2
.ends DP8TVar20ArrayShWL2_1X2

.subckt DP8TVar20ArrayShWL2_1X4 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3]
Xinst0x0 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TVar20ArrayShWL2_1X2
Xinst0x1 vss vdd wl1[0] wl2[0] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar20ArrayShWL2_1X2
.ends DP8TVar20ArrayShWL2_1X4

.subckt DP8TVar20ArrayShWL2_1X8 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss vdd wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TVar20ArrayShWL2_1X4
Xinst0x1 vss vdd wl1[0] wl2[0] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar20ArrayShWL2_1X4
.ends DP8TVar20ArrayShWL2_1X8

.subckt DP8TVar20Array_6X8 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar20Array_4X8
Xinst1x0 vss vdd wl1[4] wl2[4] wl1[5] wl2[5] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TVar20Array_2X8
.ends DP8TVar20Array_6X8

.subckt DP8TVar20TestArray_16X8C vss vdd wl1 wl2 bl1 bl1_n bl2 bl2_n bit bit_n
Xbcconn_bot vss vdd bcconn_bot_bl1[0] bcconn_bot_bl1_n[0] bcconn_bot_bl2[0] bcconn_bot_bl2_n[0] bcconn_bot_bl1[1] bcconn_bot_bl1_n[1] bcconn_bot_bl2[1] bcconn_bot_bl2_n[1] bcconn_bot_bl1[2] bcconn_bot_bl1_n[2] bcconn_bot_bl2[2] bcconn_bot_bl2_n[2] bcconn_bot_bl1[3] bcconn_bot_bl1_n[3] bcconn_bot_bl2[3] bcconn_bot_bl2_n[3] bl1 bl1_n bl2 bl2_n bcconn_bot_bl1[5] bcconn_bot_bl1_n[5] bcconn_bot_bl2[5] bcconn_bot_bl2_n[5] bcconn_bot_bl1[6] bcconn_bot_bl1_n[6] bcconn_bot_bl2[6] bcconn_bot_bl2_n[6] bcconn_bot_bl1[7] bcconn_bot_bl1_n[7] bcconn_bot_bl2[7] bcconn_bot_bl2_n[7] DP8TVar20BulkConnRow_8
Xbcconn_top vss vdd bcconn_top_bl1[0] bcconn_top_bl1_n[0] bcconn_top_bl2[0] bcconn_top_bl2_n[0] bcconn_top_bl1[1] bcconn_top_bl1_n[1] bcconn_top_bl2[1] bcconn_top_bl2_n[1] bcconn_top_bl1[2] bcconn_top_bl1_n[2] bcconn_top_bl2[2] bcconn_top_bl2_n[2] bcconn_top_bl1[3] bcconn_top_bl1_n[3] bcconn_top_bl2[3] bcconn_top_bl2_n[3] bl1 bl1_n bl2 bl2_n bcconn_top_bl1[5] bcconn_top_bl1_n[5] bcconn_top_bl2[5] bcconn_top_bl2_n[5] bcconn_top_bl1[6] bcconn_top_bl1_n[6] bcconn_top_bl2[6] bcconn_top_bl2_n[6] bcconn_top_bl1[7] bcconn_top_bl1_n[7] bcconn_top_bl2[7] bcconn_top_bl2_n[7] DP8TVar20BulkConnRow_8
Xarray_bot vss vdd zero zero zero zero zero zero zero zero zero zero zero zero zero zero array_bot_bl1[0] array_bot_bl1_n[0] array_bot_bl2[0] array_bot_bl2_n[0] array_bot_bl1[1] array_bot_bl1_n[1] array_bot_bl2[1] array_bot_bl2_n[1] array_bot_bl1[2] array_bot_bl1_n[2] array_bot_bl2[2] array_bot_bl2_n[2] array_bot_bl1[3] array_bot_bl1_n[3] array_bot_bl2[3] array_bot_bl2_n[3] bl1 bl1_n bl2 bl2_n array_bot_bl1[5] array_bot_bl1_n[5] array_bot_bl2[5] array_bot_bl2_n[5] array_bot_bl1[6] array_bot_bl1_n[6] array_bot_bl2[6] array_bot_bl2_n[6] array_bot_bl1[7] array_bot_bl1_n[7] array_bot_bl2[7] array_bot_bl2_n[7] DP8TVar20Array_7X8
Xshwl1_row vss vdd zero bit shwl1_row_bl1[0] shwl1_row_bl1_n[0] shwl1_row_bl2[0] shwl1_row_bl2_n[0] shwl1_row_bl1[1] shwl1_row_bl1_n[1] shwl1_row_bl2[1] shwl1_row_bl2_n[1] shwl1_row_bl1[2] shwl1_row_bl1_n[2] shwl1_row_bl2[2] shwl1_row_bl2_n[2] shwl1_row_bl1[3] shwl1_row_bl1_n[3] shwl1_row_bl2[3] shwl1_row_bl2_n[3] bl1 bl1_n bl2 bl2_n shwl1_row_bl1[5] shwl1_row_bl1_n[5] shwl1_row_bl2[5] shwl1_row_bl2_n[5] shwl1_row_bl1[6] shwl1_row_bl1_n[6] shwl1_row_bl2[6] shwl1_row_bl2_n[6] shwl1_row_bl1[7] shwl1_row_bl1_n[7] shwl1_row_bl2[7] shwl1_row_bl2_n[7] DP8TVar20ArrayShWL1_1X8
Xcell_cols_left vss vdd wl1 wl2 cell_cols_left_bl1[0] cell_cols_left_bl1_n[0] cell_cols_left_bl2[0] cell_cols_left_bl2_n[0] cell_cols_left_bl1[1] cell_cols_left_bl1_n[1] cell_cols_left_bl2[1] cell_cols_left_bl2_n[1] cell_cols_left_bl1[2] cell_cols_left_bl1_n[2] cell_cols_left_bl2[2] cell_cols_left_bl2_n[2] cell_cols_left_bl1[3] cell_cols_left_bl1_n[3] cell_cols_left_bl2[3] cell_cols_left_bl2_n[3] DP8TVar20Array_1X4
Xconncell wl1 wl2 bl1 bl1_n bl2 bl2_n vdd vss bit bit_n DP8TVar20CellConnectOut
Xfillcell wl1 wl2 fillcell_bl1 fillcell_bl1_n fillcell_bl2 fillcell_bl2_n vdd vss DP8TVar20Cell
Xcell_cols_right vss vdd wl1 wl2 cell_cols_right_bl1[0] cell_cols_right_bl1_n[0] cell_cols_right_bl2[0] cell_cols_right_bl2_n[0] cell_cols_right_bl1[1] cell_cols_right_bl1_n[1] cell_cols_right_bl2[1] cell_cols_right_bl2_n[1] DP8TVar20Array_1X2
Xshwl2_row vss vdd bit_n zero shwl2_row_bl1[0] shwl2_row_bl1_n[0] shwl2_row_bl2[0] shwl2_row_bl2_n[0] shwl2_row_bl1[1] shwl2_row_bl1_n[1] shwl2_row_bl2[1] shwl2_row_bl2_n[1] shwl2_row_bl1[2] shwl2_row_bl1_n[2] shwl2_row_bl2[2] shwl2_row_bl2_n[2] shwl2_row_bl1[3] shwl2_row_bl1_n[3] shwl2_row_bl2[3] shwl2_row_bl2_n[3] bl1 bl1_n bl2 bl2_n shwl2_row_bl1[5] shwl2_row_bl1_n[5] shwl2_row_bl2[5] shwl2_row_bl2_n[5] shwl2_row_bl1[6] shwl2_row_bl1_n[6] shwl2_row_bl2[6] shwl2_row_bl2_n[6] shwl2_row_bl1[7] shwl2_row_bl1_n[7] shwl2_row_bl2[7] shwl2_row_bl2_n[7] DP8TVar20ArrayShWL2_1X8
Xarray_top vss vdd zero zero zero zero zero zero zero zero zero zero zero zero array_top_bl1[0] array_top_bl1_n[0] array_top_bl2[0] array_top_bl2_n[0] array_top_bl1[1] array_top_bl1_n[1] array_top_bl2[1] array_top_bl2_n[1] array_top_bl1[2] array_top_bl1_n[2] array_top_bl2[2] array_top_bl2_n[2] array_top_bl1[3] array_top_bl1_n[3] array_top_bl2[3] array_top_bl2_n[3] bl1 bl1_n bl2 bl2_n array_top_bl1[5] array_top_bl1_n[5] array_top_bl2[5] array_top_bl2_n[5] array_top_bl1[6] array_top_bl1_n[6] array_top_bl2[6] array_top_bl2_n[6] array_top_bl1[7] array_top_bl1_n[7] array_top_bl2[7] array_top_bl2_n[7] DP8TVar20Array_6X8
Xzero vdd vss zero zero_x1
.ends DP8TVar20TestArray_16X8C

.subckt DP8TVar20 vss noco_vdd noco_wl1 noco_wl2 noco_bl1 noco_bl1_n noco_bl2 noco_bl2_n co_vdd co_bit co_bit_n co_wl1 co_wl2 co_bl1 co_bl1_n co_bl2_n co_bl2
Xframe noco_vdd noco_wl1 noco_wl2 noco_bl2 co_vdd co_bit co_bit_n co_wl1 co_wl2 NoConn_PAD0x9 vss noco_bl1 noco_bl1_n noco_bl2_n vss co_bl1 co_bl1_n co_bl2_n co_bl2 NoConn_PAD1x9 PadFrame_DP20
Xtestarray_noco vss noco_vdd noco_wl1 noco_wl2 noco_bl1 noco_bl1_n noco_bl2 noco_bl2_n DP8TVar20TestArray_16X8
Xtestarray_co vss co_vdd co_wl1 co_wl2 co_bl1 co_bl1_n co_bl2 co_bl2_n co_bit co_bit_n DP8TVar20TestArray_16X8C
.ends DP8TVar20

.subckt SingleCell_TestStructures vss sp6tvar0_noco_vdd sp6tvar0_noco_wl sp6tvar0_noco_bl sp6tvar0_noco_bl_n sp6tvar0_co_vdd sp6tvar0_co_bl sp6tvar0_co_bl_n sp6tvar0_co_bit sp6tvar0_co_bit_n sp6tvar0_co_wl sp6tvar1_noco_vdd sp6tvar1_noco_wl sp6tvar1_noco_bl sp6tvar1_noco_bl_n sp6tvar1_co_vdd sp6tvar1_co_bl sp6tvar1_co_bl_n sp6tvar1_co_bit sp6tvar1_co_bit_n sp6tvar1_co_wl sp6tvar2_noco_vdd sp6tvar2_noco_wl sp6tvar2_noco_bl sp6tvar2_noco_bl_n sp6tvar2_co_vdd sp6tvar2_co_bl sp6tvar2_co_bl_n sp6tvar2_co_bit sp6tvar2_co_bit_n sp6tvar2_co_wl sp6tvar3_noco_vdd sp6tvar3_noco_wl sp6tvar3_noco_bl sp6tvar3_noco_bl_n sp6tvar3_co_vdd sp6tvar3_co_bl sp6tvar3_co_bl_n sp6tvar3_co_bit sp6tvar3_co_bit_n sp6tvar3_co_wl sp6tvar4_noco_vdd sp6tvar4_noco_wl sp6tvar4_noco_bl sp6tvar4_noco_bl_n sp6tvar4_co_vdd sp6tvar4_co_bl sp6tvar4_co_bl_n sp6tvar4_co_bit sp6tvar4_co_bit_n sp6tvar4_co_wl sp6tvar5_noco_vdd sp6tvar5_noco_wl sp6tvar5_noco_bl sp6tvar5_noco_bl_n sp6tvar5_co_vdd sp6tvar5_co_bl sp6tvar5_co_bl_n sp6tvar5_co_bit sp6tvar5_co_bit_n sp6tvar5_co_wl sp6tvar6_noco_vdd sp6tvar6_noco_wl sp6tvar6_noco_bl sp6tvar6_noco_bl_n sp6tvar6_co_vdd sp6tvar6_co_bl sp6tvar6_co_bl_n sp6tvar6_co_bit sp6tvar6_co_bit_n sp6tvar6_co_wl sp6tvar7_noco_vdd sp6tvar7_noco_wl sp6tvar7_noco_bl sp6tvar7_noco_bl_n sp6tvar7_co_vdd sp6tvar7_co_bl sp6tvar7_co_bl_n sp6tvar7_co_bit sp6tvar7_co_bit_n sp6tvar7_co_wl sp6tvar8_noco_vdd sp6tvar8_noco_wl sp6tvar8_noco_bl sp6tvar8_noco_bl_n sp6tvar8_co_vdd sp6tvar8_co_bl sp6tvar8_co_bl_n sp6tvar8_co_bit sp6tvar8_co_bit_n sp6tvar8_co_wl sp6tvar9_noco_vdd sp6tvar9_noco_wl sp6tvar9_noco_bl sp6tvar9_noco_bl_n sp6tvar9_co_vdd sp6tvar9_co_bl sp6tvar9_co_bl_n sp6tvar9_co_bit sp6tvar9_co_bit_n sp6tvar9_co_wl sp6tvar10_noco_vdd sp6tvar10_noco_wl sp6tvar10_noco_bl sp6tvar10_noco_bl_n sp6tvar10_co_vdd sp6tvar10_co_bl sp6tvar10_co_bl_n sp6tvar10_co_bit sp6tvar10_co_bit_n sp6tvar10_co_wl sp6tvar11_noco_vdd sp6tvar11_noco_wl sp6tvar11_noco_bl sp6tvar11_noco_bl_n sp6tvar11_co_vdd sp6tvar11_co_bl sp6tvar11_co_bl_n sp6tvar11_co_bit sp6tvar11_co_bit_n sp6tvar11_co_wl sp6tvar12_noco_vdd sp6tvar12_noco_wl sp6tvar12_noco_bl sp6tvar12_noco_bl_n sp6tvar12_co_vdd sp6tvar12_co_bl sp6tvar12_co_bl_n sp6tvar12_co_bit sp6tvar12_co_bit_n sp6tvar12_co_wl sp6tvar13_noco_vdd sp6tvar13_noco_wl sp6tvar13_noco_bl sp6tvar13_noco_bl_n sp6tvar13_co_vdd sp6tvar13_co_bl sp6tvar13_co_bl_n sp6tvar13_co_bit sp6tvar13_co_bit_n sp6tvar13_co_wl sp6tvar14_noco_vdd sp6tvar14_noco_wl sp6tvar14_noco_bl sp6tvar14_noco_bl_n sp6tvar14_co_vdd sp6tvar14_co_bl sp6tvar14_co_bl_n sp6tvar14_co_bit sp6tvar14_co_bit_n sp6tvar14_co_wl sp6tvar15_noco_vdd sp6tvar15_noco_wl sp6tvar15_noco_bl sp6tvar15_noco_bl_n sp6tvar15_co_vdd sp6tvar15_co_bl sp6tvar15_co_bl_n sp6tvar15_co_bit sp6tvar15_co_bit_n sp6tvar15_co_wl sp6tvar16_noco_vdd sp6tvar16_noco_wl sp6tvar16_noco_bl sp6tvar16_noco_bl_n sp6tvar16_co_vdd sp6tvar16_co_bl sp6tvar16_co_bl_n sp6tvar16_co_bit sp6tvar16_co_bit_n sp6tvar16_co_wl sp6tvar17_noco_vdd sp6tvar17_noco_wl sp6tvar17_noco_bl sp6tvar17_noco_bl_n sp6tvar17_co_vdd sp6tvar17_co_bl sp6tvar17_co_bl_n sp6tvar17_co_bit sp6tvar17_co_bit_n sp6tvar17_co_wl sp6tvar18_noco_vdd sp6tvar18_noco_wl sp6tvar18_noco_bl sp6tvar18_noco_bl_n sp6tvar18_co_vdd sp6tvar18_co_bl sp6tvar18_co_bl_n sp6tvar18_co_bit sp6tvar18_co_bit_n sp6tvar18_co_wl sp6tvar19_noco_vdd sp6tvar19_noco_wl sp6tvar19_noco_bl sp6tvar19_noco_bl_n sp6tvar19_co_vdd sp6tvar19_co_bl sp6tvar19_co_bl_n sp6tvar19_co_bit sp6tvar19_co_bit_n sp6tvar19_co_wl sp6tvar20_noco_vdd sp6tvar20_noco_wl sp6tvar20_noco_bl sp6tvar20_noco_bl_n sp6tvar20_co_vdd sp6tvar20_co_bl sp6tvar20_co_bl_n sp6tvar20_co_bit sp6tvar20_co_bit_n sp6tvar20_co_wl sp6tvar21_noco_vdd sp6tvar21_noco_wl sp6tvar21_noco_bl sp6tvar21_noco_bl_n sp6tvar21_co_vdd sp6tvar21_co_bl sp6tvar21_co_bl_n sp6tvar21_co_bit sp6tvar21_co_bit_n sp6tvar21_co_wl sp6tvar22_noco_vdd sp6tvar22_noco_wl sp6tvar22_noco_bl sp6tvar22_noco_bl_n sp6tvar22_co_vdd sp6tvar22_co_bl sp6tvar22_co_bl_n sp6tvar22_co_bit sp6tvar22_co_bit_n sp6tvar22_co_wl dp8tvar0_noco_vdd dp8tvar0_noco_wl1 dp8tvar0_noco_wl2 dp8tvar0_noco_bl1 dp8tvar0_noco_bl1_n dp8tvar0_noco_bl2 dp8tvar0_noco_bl2_n dp8tvar0_co_vdd dp8tvar0_co_bit dp8tvar0_co_bit_n dp8tvar0_co_wl1 dp8tvar0_co_wl2 dp8tvar0_co_bl1 dp8tvar0_co_bl1_n dp8tvar0_co_bl2_n dp8tvar0_co_bl2 dp8tvar1_noco_vdd dp8tvar1_noco_wl1 dp8tvar1_noco_wl2 dp8tvar1_noco_bl1 dp8tvar1_noco_bl1_n dp8tvar1_noco_bl2 dp8tvar1_noco_bl2_n dp8tvar1_co_vdd dp8tvar1_co_bit dp8tvar1_co_bit_n dp8tvar1_co_wl1 dp8tvar1_co_wl2 dp8tvar1_co_bl1 dp8tvar1_co_bl1_n dp8tvar1_co_bl2_n dp8tvar1_co_bl2 dp8tvar2_noco_vdd dp8tvar2_noco_wl1 dp8tvar2_noco_wl2 dp8tvar2_noco_bl1 dp8tvar2_noco_bl1_n dp8tvar2_noco_bl2 dp8tvar2_noco_bl2_n dp8tvar2_co_vdd dp8tvar2_co_bit dp8tvar2_co_bit_n dp8tvar2_co_wl1 dp8tvar2_co_wl2 dp8tvar2_co_bl1 dp8tvar2_co_bl1_n dp8tvar2_co_bl2_n dp8tvar2_co_bl2 dp8tvar3_noco_vdd dp8tvar3_noco_wl1 dp8tvar3_noco_wl2 dp8tvar3_noco_bl1 dp8tvar3_noco_bl1_n dp8tvar3_noco_bl2 dp8tvar3_noco_bl2_n dp8tvar3_co_vdd dp8tvar3_co_bit dp8tvar3_co_bit_n dp8tvar3_co_wl1 dp8tvar3_co_wl2 dp8tvar3_co_bl1 dp8tvar3_co_bl1_n dp8tvar3_co_bl2_n dp8tvar3_co_bl2 dp8tvar4_noco_vdd dp8tvar4_noco_wl1 dp8tvar4_noco_wl2 dp8tvar4_noco_bl1 dp8tvar4_noco_bl1_n dp8tvar4_noco_bl2 dp8tvar4_noco_bl2_n dp8tvar4_co_vdd dp8tvar4_co_bit dp8tvar4_co_bit_n dp8tvar4_co_wl1 dp8tvar4_co_wl2 dp8tvar4_co_bl1 dp8tvar4_co_bl1_n dp8tvar4_co_bl2_n dp8tvar4_co_bl2 dp8tvar5_noco_vdd dp8tvar5_noco_wl1 dp8tvar5_noco_wl2 dp8tvar5_noco_bl1 dp8tvar5_noco_bl1_n dp8tvar5_noco_bl2 dp8tvar5_noco_bl2_n dp8tvar5_co_vdd dp8tvar5_co_bit dp8tvar5_co_bit_n dp8tvar5_co_wl1 dp8tvar5_co_wl2 dp8tvar5_co_bl1 dp8tvar5_co_bl1_n dp8tvar5_co_bl2_n dp8tvar5_co_bl2 dp8tvar6_noco_vdd dp8tvar6_noco_wl1 dp8tvar6_noco_wl2 dp8tvar6_noco_bl1 dp8tvar6_noco_bl1_n dp8tvar6_noco_bl2 dp8tvar6_noco_bl2_n dp8tvar6_co_vdd dp8tvar6_co_bit dp8tvar6_co_bit_n dp8tvar6_co_wl1 dp8tvar6_co_wl2 dp8tvar6_co_bl1 dp8tvar6_co_bl1_n dp8tvar6_co_bl2_n dp8tvar6_co_bl2 dp8tvar7_noco_vdd dp8tvar7_noco_wl1 dp8tvar7_noco_wl2 dp8tvar7_noco_bl1 dp8tvar7_noco_bl1_n dp8tvar7_noco_bl2 dp8tvar7_noco_bl2_n dp8tvar7_co_vdd dp8tvar7_co_bit dp8tvar7_co_bit_n dp8tvar7_co_wl1 dp8tvar7_co_wl2 dp8tvar7_co_bl1 dp8tvar7_co_bl1_n dp8tvar7_co_bl2_n dp8tvar7_co_bl2 dp8tvar8_noco_vdd dp8tvar8_noco_wl1 dp8tvar8_noco_wl2 dp8tvar8_noco_bl1 dp8tvar8_noco_bl1_n dp8tvar8_noco_bl2 dp8tvar8_noco_bl2_n dp8tvar8_co_vdd dp8tvar8_co_bit dp8tvar8_co_bit_n dp8tvar8_co_wl1 dp8tvar8_co_wl2 dp8tvar8_co_bl1 dp8tvar8_co_bl1_n dp8tvar8_co_bl2_n dp8tvar8_co_bl2 dp8tvar9_noco_vdd dp8tvar9_noco_wl1 dp8tvar9_noco_wl2 dp8tvar9_noco_bl1 dp8tvar9_noco_bl1_n dp8tvar9_noco_bl2 dp8tvar9_noco_bl2_n dp8tvar9_co_vdd dp8tvar9_co_bit dp8tvar9_co_bit_n dp8tvar9_co_wl1 dp8tvar9_co_wl2 dp8tvar9_co_bl1 dp8tvar9_co_bl1_n dp8tvar9_co_bl2_n dp8tvar9_co_bl2 dp8tvar10_noco_vdd dp8tvar10_noco_wl1 dp8tvar10_noco_wl2 dp8tvar10_noco_bl1 dp8tvar10_noco_bl1_n dp8tvar10_noco_bl2 dp8tvar10_noco_bl2_n dp8tvar10_co_vdd dp8tvar10_co_bit dp8tvar10_co_bit_n dp8tvar10_co_wl1 dp8tvar10_co_wl2 dp8tvar10_co_bl1 dp8tvar10_co_bl1_n dp8tvar10_co_bl2_n dp8tvar10_co_bl2 dp8tvar11_noco_vdd dp8tvar11_noco_wl1 dp8tvar11_noco_wl2 dp8tvar11_noco_bl1 dp8tvar11_noco_bl1_n dp8tvar11_noco_bl2 dp8tvar11_noco_bl2_n dp8tvar11_co_vdd dp8tvar11_co_bit dp8tvar11_co_bit_n dp8tvar11_co_wl1 dp8tvar11_co_wl2 dp8tvar11_co_bl1 dp8tvar11_co_bl1_n dp8tvar11_co_bl2_n dp8tvar11_co_bl2 dp8tvar12_noco_vdd dp8tvar12_noco_wl1 dp8tvar12_noco_wl2 dp8tvar12_noco_bl1 dp8tvar12_noco_bl1_n dp8tvar12_noco_bl2 dp8tvar12_noco_bl2_n dp8tvar12_co_vdd dp8tvar12_co_bit dp8tvar12_co_bit_n dp8tvar12_co_wl1 dp8tvar12_co_wl2 dp8tvar12_co_bl1 dp8tvar12_co_bl1_n dp8tvar12_co_bl2_n dp8tvar12_co_bl2 dp8tvar13_noco_vdd dp8tvar13_noco_wl1 dp8tvar13_noco_wl2 dp8tvar13_noco_bl1 dp8tvar13_noco_bl1_n dp8tvar13_noco_bl2 dp8tvar13_noco_bl2_n dp8tvar13_co_vdd dp8tvar13_co_bit dp8tvar13_co_bit_n dp8tvar13_co_wl1 dp8tvar13_co_wl2 dp8tvar13_co_bl1 dp8tvar13_co_bl1_n dp8tvar13_co_bl2_n dp8tvar13_co_bl2 dp8tvar14_noco_vdd dp8tvar14_noco_wl1 dp8tvar14_noco_wl2 dp8tvar14_noco_bl1 dp8tvar14_noco_bl1_n dp8tvar14_noco_bl2 dp8tvar14_noco_bl2_n dp8tvar14_co_vdd dp8tvar14_co_bit dp8tvar14_co_bit_n dp8tvar14_co_wl1 dp8tvar14_co_wl2 dp8tvar14_co_bl1 dp8tvar14_co_bl1_n dp8tvar14_co_bl2_n dp8tvar14_co_bl2 dp8tvar15_noco_vdd dp8tvar15_noco_wl1 dp8tvar15_noco_wl2 dp8tvar15_noco_bl1 dp8tvar15_noco_bl1_n dp8tvar15_noco_bl2 dp8tvar15_noco_bl2_n dp8tvar15_co_vdd dp8tvar15_co_bit dp8tvar15_co_bit_n dp8tvar15_co_wl1 dp8tvar15_co_wl2 dp8tvar15_co_bl1 dp8tvar15_co_bl1_n dp8tvar15_co_bl2_n dp8tvar15_co_bl2 dp8tvar16_noco_vdd dp8tvar16_noco_wl1 dp8tvar16_noco_wl2 dp8tvar16_noco_bl1 dp8tvar16_noco_bl1_n dp8tvar16_noco_bl2 dp8tvar16_noco_bl2_n dp8tvar16_co_vdd dp8tvar16_co_bit dp8tvar16_co_bit_n dp8tvar16_co_wl1 dp8tvar16_co_wl2 dp8tvar16_co_bl1 dp8tvar16_co_bl1_n dp8tvar16_co_bl2_n dp8tvar16_co_bl2 dp8tvar17_noco_vdd dp8tvar17_noco_wl1 dp8tvar17_noco_wl2 dp8tvar17_noco_bl1 dp8tvar17_noco_bl1_n dp8tvar17_noco_bl2 dp8tvar17_noco_bl2_n dp8tvar17_co_vdd dp8tvar17_co_bit dp8tvar17_co_bit_n dp8tvar17_co_wl1 dp8tvar17_co_wl2 dp8tvar17_co_bl1 dp8tvar17_co_bl1_n dp8tvar17_co_bl2_n dp8tvar17_co_bl2 dp8tvar18_noco_vdd dp8tvar18_noco_wl1 dp8tvar18_noco_wl2 dp8tvar18_noco_bl1 dp8tvar18_noco_bl1_n dp8tvar18_noco_bl2 dp8tvar18_noco_bl2_n dp8tvar18_co_vdd dp8tvar18_co_bit dp8tvar18_co_bit_n dp8tvar18_co_wl1 dp8tvar18_co_wl2 dp8tvar18_co_bl1 dp8tvar18_co_bl1_n dp8tvar18_co_bl2_n dp8tvar18_co_bl2 dp8tvar19_noco_vdd dp8tvar19_noco_wl1 dp8tvar19_noco_wl2 dp8tvar19_noco_bl1 dp8tvar19_noco_bl1_n dp8tvar19_noco_bl2 dp8tvar19_noco_bl2_n dp8tvar19_co_vdd dp8tvar19_co_bit dp8tvar19_co_bit_n dp8tvar19_co_wl1 dp8tvar19_co_wl2 dp8tvar19_co_bl1 dp8tvar19_co_bl1_n dp8tvar19_co_bl2_n dp8tvar19_co_bl2 dp8tvar20_noco_vdd dp8tvar20_noco_wl1 dp8tvar20_noco_wl2 dp8tvar20_noco_bl1 dp8tvar20_noco_bl1_n dp8tvar20_noco_bl2 dp8tvar20_noco_bl2_n dp8tvar20_co_vdd dp8tvar20_co_bit dp8tvar20_co_bit_n dp8tvar20_co_wl1 dp8tvar20_co_wl2 dp8tvar20_co_bl1 dp8tvar20_co_bl1_n dp8tvar20_co_bl2_n dp8tvar20_co_bl2
Xsp6tvar0 vss sp6tvar0_noco_vdd sp6tvar0_noco_wl sp6tvar0_noco_bl sp6tvar0_noco_bl_n sp6tvar0_co_vdd sp6tvar0_co_bl sp6tvar0_co_bl_n sp6tvar0_co_bit sp6tvar0_co_bit_n sp6tvar0_co_wl SP6TVar0
Xsp6tvar1 vss sp6tvar1_noco_vdd sp6tvar1_noco_wl sp6tvar1_noco_bl sp6tvar1_noco_bl_n sp6tvar1_co_vdd sp6tvar1_co_bl sp6tvar1_co_bl_n sp6tvar1_co_bit sp6tvar1_co_bit_n sp6tvar1_co_wl SP6TVar1
Xsp6tvar2 vss sp6tvar2_noco_vdd sp6tvar2_noco_wl sp6tvar2_noco_bl sp6tvar2_noco_bl_n sp6tvar2_co_vdd sp6tvar2_co_bl sp6tvar2_co_bl_n sp6tvar2_co_bit sp6tvar2_co_bit_n sp6tvar2_co_wl SP6TVar2
Xsp6tvar3 vss sp6tvar3_noco_vdd sp6tvar3_noco_wl sp6tvar3_noco_bl sp6tvar3_noco_bl_n sp6tvar3_co_vdd sp6tvar3_co_bl sp6tvar3_co_bl_n sp6tvar3_co_bit sp6tvar3_co_bit_n sp6tvar3_co_wl SP6TVar3
Xsp6tvar4 vss sp6tvar4_noco_vdd sp6tvar4_noco_wl sp6tvar4_noco_bl sp6tvar4_noco_bl_n sp6tvar4_co_vdd sp6tvar4_co_bl sp6tvar4_co_bl_n sp6tvar4_co_bit sp6tvar4_co_bit_n sp6tvar4_co_wl SP6TVar4
Xsp6tvar5 vss sp6tvar5_noco_vdd sp6tvar5_noco_wl sp6tvar5_noco_bl sp6tvar5_noco_bl_n sp6tvar5_co_vdd sp6tvar5_co_bl sp6tvar5_co_bl_n sp6tvar5_co_bit sp6tvar5_co_bit_n sp6tvar5_co_wl SP6TVar5
Xsp6tvar6 vss sp6tvar6_noco_vdd sp6tvar6_noco_wl sp6tvar6_noco_bl sp6tvar6_noco_bl_n sp6tvar6_co_vdd sp6tvar6_co_bl sp6tvar6_co_bl_n sp6tvar6_co_bit sp6tvar6_co_bit_n sp6tvar6_co_wl SP6TVar6
Xsp6tvar7 vss sp6tvar7_noco_vdd sp6tvar7_noco_wl sp6tvar7_noco_bl sp6tvar7_noco_bl_n sp6tvar7_co_vdd sp6tvar7_co_bl sp6tvar7_co_bl_n sp6tvar7_co_bit sp6tvar7_co_bit_n sp6tvar7_co_wl SP6TVar7
Xsp6tvar8 vss sp6tvar8_noco_vdd sp6tvar8_noco_wl sp6tvar8_noco_bl sp6tvar8_noco_bl_n sp6tvar8_co_vdd sp6tvar8_co_bl sp6tvar8_co_bl_n sp6tvar8_co_bit sp6tvar8_co_bit_n sp6tvar8_co_wl SP6TVar8
Xsp6tvar9 vss sp6tvar9_noco_vdd sp6tvar9_noco_wl sp6tvar9_noco_bl sp6tvar9_noco_bl_n sp6tvar9_co_vdd sp6tvar9_co_bl sp6tvar9_co_bl_n sp6tvar9_co_bit sp6tvar9_co_bit_n sp6tvar9_co_wl SP6TVar9
Xsp6tvar10 vss sp6tvar10_noco_vdd sp6tvar10_noco_wl sp6tvar10_noco_bl sp6tvar10_noco_bl_n sp6tvar10_co_vdd sp6tvar10_co_bl sp6tvar10_co_bl_n sp6tvar10_co_bit sp6tvar10_co_bit_n sp6tvar10_co_wl SP6TVar10
Xsp6tvar11 vss sp6tvar11_noco_vdd sp6tvar11_noco_wl sp6tvar11_noco_bl sp6tvar11_noco_bl_n sp6tvar11_co_vdd sp6tvar11_co_bl sp6tvar11_co_bl_n sp6tvar11_co_bit sp6tvar11_co_bit_n sp6tvar11_co_wl SP6TVar11
Xsp6tvar12 vss sp6tvar12_noco_vdd sp6tvar12_noco_wl sp6tvar12_noco_bl sp6tvar12_noco_bl_n sp6tvar12_co_vdd sp6tvar12_co_bl sp6tvar12_co_bl_n sp6tvar12_co_bit sp6tvar12_co_bit_n sp6tvar12_co_wl SP6TVar12
Xsp6tvar13 vss sp6tvar13_noco_vdd sp6tvar13_noco_wl sp6tvar13_noco_bl sp6tvar13_noco_bl_n sp6tvar13_co_vdd sp6tvar13_co_bl sp6tvar13_co_bl_n sp6tvar13_co_bit sp6tvar13_co_bit_n sp6tvar13_co_wl SP6TVar13
Xsp6tvar14 vss sp6tvar14_noco_vdd sp6tvar14_noco_wl sp6tvar14_noco_bl sp6tvar14_noco_bl_n sp6tvar14_co_vdd sp6tvar14_co_bl sp6tvar14_co_bl_n sp6tvar14_co_bit sp6tvar14_co_bit_n sp6tvar14_co_wl SP6TVar14
Xsp6tvar15 vss sp6tvar15_noco_vdd sp6tvar15_noco_wl sp6tvar15_noco_bl sp6tvar15_noco_bl_n sp6tvar15_co_vdd sp6tvar15_co_bl sp6tvar15_co_bl_n sp6tvar15_co_bit sp6tvar15_co_bit_n sp6tvar15_co_wl SP6TVar15
Xsp6tvar16 vss sp6tvar16_noco_vdd sp6tvar16_noco_wl sp6tvar16_noco_bl sp6tvar16_noco_bl_n sp6tvar16_co_vdd sp6tvar16_co_bl sp6tvar16_co_bl_n sp6tvar16_co_bit sp6tvar16_co_bit_n sp6tvar16_co_wl SP6TVar16
Xsp6tvar17 vss sp6tvar17_noco_vdd sp6tvar17_noco_wl sp6tvar17_noco_bl sp6tvar17_noco_bl_n sp6tvar17_co_vdd sp6tvar17_co_bl sp6tvar17_co_bl_n sp6tvar17_co_bit sp6tvar17_co_bit_n sp6tvar17_co_wl SP6TVar17
Xsp6tvar18 vss sp6tvar18_noco_vdd sp6tvar18_noco_wl sp6tvar18_noco_bl sp6tvar18_noco_bl_n sp6tvar18_co_vdd sp6tvar18_co_bl sp6tvar18_co_bl_n sp6tvar18_co_bit sp6tvar18_co_bit_n sp6tvar18_co_wl SP6TVar18
Xsp6tvar19 vss sp6tvar19_noco_vdd sp6tvar19_noco_wl sp6tvar19_noco_bl sp6tvar19_noco_bl_n sp6tvar19_co_vdd sp6tvar19_co_bl sp6tvar19_co_bl_n sp6tvar19_co_bit sp6tvar19_co_bit_n sp6tvar19_co_wl SP6TVar19
Xsp6tvar20 vss sp6tvar20_noco_vdd sp6tvar20_noco_wl sp6tvar20_noco_bl sp6tvar20_noco_bl_n sp6tvar20_co_vdd sp6tvar20_co_bl sp6tvar20_co_bl_n sp6tvar20_co_bit sp6tvar20_co_bit_n sp6tvar20_co_wl SP6TVar20
Xsp6tvar21 vss sp6tvar21_noco_vdd sp6tvar21_noco_wl sp6tvar21_noco_bl sp6tvar21_noco_bl_n sp6tvar21_co_vdd sp6tvar21_co_bl sp6tvar21_co_bl_n sp6tvar21_co_bit sp6tvar21_co_bit_n sp6tvar21_co_wl SP6TVar21
Xsp6tvar22 vss sp6tvar22_noco_vdd sp6tvar22_noco_wl sp6tvar22_noco_bl sp6tvar22_noco_bl_n sp6tvar22_co_vdd sp6tvar22_co_bl sp6tvar22_co_bl_n sp6tvar22_co_bit sp6tvar22_co_bit_n sp6tvar22_co_wl SP6TVar22
Xdp8tvar0 vss dp8tvar0_noco_vdd dp8tvar0_noco_wl1 dp8tvar0_noco_wl2 dp8tvar0_noco_bl1 dp8tvar0_noco_bl1_n dp8tvar0_noco_bl2 dp8tvar0_noco_bl2_n dp8tvar0_co_vdd dp8tvar0_co_bit dp8tvar0_co_bit_n dp8tvar0_co_wl1 dp8tvar0_co_wl2 dp8tvar0_co_bl1 dp8tvar0_co_bl1_n dp8tvar0_co_bl2_n dp8tvar0_co_bl2 DP8TVar0
Xdp8tvar1 vss dp8tvar1_noco_vdd dp8tvar1_noco_wl1 dp8tvar1_noco_wl2 dp8tvar1_noco_bl1 dp8tvar1_noco_bl1_n dp8tvar1_noco_bl2 dp8tvar1_noco_bl2_n dp8tvar1_co_vdd dp8tvar1_co_bit dp8tvar1_co_bit_n dp8tvar1_co_wl1 dp8tvar1_co_wl2 dp8tvar1_co_bl1 dp8tvar1_co_bl1_n dp8tvar1_co_bl2_n dp8tvar1_co_bl2 DP8TVar1
Xdp8tvar2 vss dp8tvar2_noco_vdd dp8tvar2_noco_wl1 dp8tvar2_noco_wl2 dp8tvar2_noco_bl1 dp8tvar2_noco_bl1_n dp8tvar2_noco_bl2 dp8tvar2_noco_bl2_n dp8tvar2_co_vdd dp8tvar2_co_bit dp8tvar2_co_bit_n dp8tvar2_co_wl1 dp8tvar2_co_wl2 dp8tvar2_co_bl1 dp8tvar2_co_bl1_n dp8tvar2_co_bl2_n dp8tvar2_co_bl2 DP8TVar2
Xdp8tvar3 vss dp8tvar3_noco_vdd dp8tvar3_noco_wl1 dp8tvar3_noco_wl2 dp8tvar3_noco_bl1 dp8tvar3_noco_bl1_n dp8tvar3_noco_bl2 dp8tvar3_noco_bl2_n dp8tvar3_co_vdd dp8tvar3_co_bit dp8tvar3_co_bit_n dp8tvar3_co_wl1 dp8tvar3_co_wl2 dp8tvar3_co_bl1 dp8tvar3_co_bl1_n dp8tvar3_co_bl2_n dp8tvar3_co_bl2 DP8TVar3
Xdp8tvar4 vss dp8tvar4_noco_vdd dp8tvar4_noco_wl1 dp8tvar4_noco_wl2 dp8tvar4_noco_bl1 dp8tvar4_noco_bl1_n dp8tvar4_noco_bl2 dp8tvar4_noco_bl2_n dp8tvar4_co_vdd dp8tvar4_co_bit dp8tvar4_co_bit_n dp8tvar4_co_wl1 dp8tvar4_co_wl2 dp8tvar4_co_bl1 dp8tvar4_co_bl1_n dp8tvar4_co_bl2_n dp8tvar4_co_bl2 DP8TVar4
Xdp8tvar5 vss dp8tvar5_noco_vdd dp8tvar5_noco_wl1 dp8tvar5_noco_wl2 dp8tvar5_noco_bl1 dp8tvar5_noco_bl1_n dp8tvar5_noco_bl2 dp8tvar5_noco_bl2_n dp8tvar5_co_vdd dp8tvar5_co_bit dp8tvar5_co_bit_n dp8tvar5_co_wl1 dp8tvar5_co_wl2 dp8tvar5_co_bl1 dp8tvar5_co_bl1_n dp8tvar5_co_bl2_n dp8tvar5_co_bl2 DP8TVar5
Xdp8tvar6 vss dp8tvar6_noco_vdd dp8tvar6_noco_wl1 dp8tvar6_noco_wl2 dp8tvar6_noco_bl1 dp8tvar6_noco_bl1_n dp8tvar6_noco_bl2 dp8tvar6_noco_bl2_n dp8tvar6_co_vdd dp8tvar6_co_bit dp8tvar6_co_bit_n dp8tvar6_co_wl1 dp8tvar6_co_wl2 dp8tvar6_co_bl1 dp8tvar6_co_bl1_n dp8tvar6_co_bl2_n dp8tvar6_co_bl2 DP8TVar6
Xdp8tvar7 vss dp8tvar7_noco_vdd dp8tvar7_noco_wl1 dp8tvar7_noco_wl2 dp8tvar7_noco_bl1 dp8tvar7_noco_bl1_n dp8tvar7_noco_bl2 dp8tvar7_noco_bl2_n dp8tvar7_co_vdd dp8tvar7_co_bit dp8tvar7_co_bit_n dp8tvar7_co_wl1 dp8tvar7_co_wl2 dp8tvar7_co_bl1 dp8tvar7_co_bl1_n dp8tvar7_co_bl2_n dp8tvar7_co_bl2 DP8TVar7
Xdp8tvar8 vss dp8tvar8_noco_vdd dp8tvar8_noco_wl1 dp8tvar8_noco_wl2 dp8tvar8_noco_bl1 dp8tvar8_noco_bl1_n dp8tvar8_noco_bl2 dp8tvar8_noco_bl2_n dp8tvar8_co_vdd dp8tvar8_co_bit dp8tvar8_co_bit_n dp8tvar8_co_wl1 dp8tvar8_co_wl2 dp8tvar8_co_bl1 dp8tvar8_co_bl1_n dp8tvar8_co_bl2_n dp8tvar8_co_bl2 DP8TVar8
Xdp8tvar9 vss dp8tvar9_noco_vdd dp8tvar9_noco_wl1 dp8tvar9_noco_wl2 dp8tvar9_noco_bl1 dp8tvar9_noco_bl1_n dp8tvar9_noco_bl2 dp8tvar9_noco_bl2_n dp8tvar9_co_vdd dp8tvar9_co_bit dp8tvar9_co_bit_n dp8tvar9_co_wl1 dp8tvar9_co_wl2 dp8tvar9_co_bl1 dp8tvar9_co_bl1_n dp8tvar9_co_bl2_n dp8tvar9_co_bl2 DP8TVar9
Xdp8tvar10 vss dp8tvar10_noco_vdd dp8tvar10_noco_wl1 dp8tvar10_noco_wl2 dp8tvar10_noco_bl1 dp8tvar10_noco_bl1_n dp8tvar10_noco_bl2 dp8tvar10_noco_bl2_n dp8tvar10_co_vdd dp8tvar10_co_bit dp8tvar10_co_bit_n dp8tvar10_co_wl1 dp8tvar10_co_wl2 dp8tvar10_co_bl1 dp8tvar10_co_bl1_n dp8tvar10_co_bl2_n dp8tvar10_co_bl2 DP8TVar10
Xdp8tvar11 vss dp8tvar11_noco_vdd dp8tvar11_noco_wl1 dp8tvar11_noco_wl2 dp8tvar11_noco_bl1 dp8tvar11_noco_bl1_n dp8tvar11_noco_bl2 dp8tvar11_noco_bl2_n dp8tvar11_co_vdd dp8tvar11_co_bit dp8tvar11_co_bit_n dp8tvar11_co_wl1 dp8tvar11_co_wl2 dp8tvar11_co_bl1 dp8tvar11_co_bl1_n dp8tvar11_co_bl2_n dp8tvar11_co_bl2 DP8TVar11
Xdp8tvar12 vss dp8tvar12_noco_vdd dp8tvar12_noco_wl1 dp8tvar12_noco_wl2 dp8tvar12_noco_bl1 dp8tvar12_noco_bl1_n dp8tvar12_noco_bl2 dp8tvar12_noco_bl2_n dp8tvar12_co_vdd dp8tvar12_co_bit dp8tvar12_co_bit_n dp8tvar12_co_wl1 dp8tvar12_co_wl2 dp8tvar12_co_bl1 dp8tvar12_co_bl1_n dp8tvar12_co_bl2_n dp8tvar12_co_bl2 DP8TVar12
Xdp8tvar13 vss dp8tvar13_noco_vdd dp8tvar13_noco_wl1 dp8tvar13_noco_wl2 dp8tvar13_noco_bl1 dp8tvar13_noco_bl1_n dp8tvar13_noco_bl2 dp8tvar13_noco_bl2_n dp8tvar13_co_vdd dp8tvar13_co_bit dp8tvar13_co_bit_n dp8tvar13_co_wl1 dp8tvar13_co_wl2 dp8tvar13_co_bl1 dp8tvar13_co_bl1_n dp8tvar13_co_bl2_n dp8tvar13_co_bl2 DP8TVar13
Xdp8tvar14 vss dp8tvar14_noco_vdd dp8tvar14_noco_wl1 dp8tvar14_noco_wl2 dp8tvar14_noco_bl1 dp8tvar14_noco_bl1_n dp8tvar14_noco_bl2 dp8tvar14_noco_bl2_n dp8tvar14_co_vdd dp8tvar14_co_bit dp8tvar14_co_bit_n dp8tvar14_co_wl1 dp8tvar14_co_wl2 dp8tvar14_co_bl1 dp8tvar14_co_bl1_n dp8tvar14_co_bl2_n dp8tvar14_co_bl2 DP8TVar14
Xdp8tvar15 vss dp8tvar15_noco_vdd dp8tvar15_noco_wl1 dp8tvar15_noco_wl2 dp8tvar15_noco_bl1 dp8tvar15_noco_bl1_n dp8tvar15_noco_bl2 dp8tvar15_noco_bl2_n dp8tvar15_co_vdd dp8tvar15_co_bit dp8tvar15_co_bit_n dp8tvar15_co_wl1 dp8tvar15_co_wl2 dp8tvar15_co_bl1 dp8tvar15_co_bl1_n dp8tvar15_co_bl2_n dp8tvar15_co_bl2 DP8TVar15
Xdp8tvar16 vss dp8tvar16_noco_vdd dp8tvar16_noco_wl1 dp8tvar16_noco_wl2 dp8tvar16_noco_bl1 dp8tvar16_noco_bl1_n dp8tvar16_noco_bl2 dp8tvar16_noco_bl2_n dp8tvar16_co_vdd dp8tvar16_co_bit dp8tvar16_co_bit_n dp8tvar16_co_wl1 dp8tvar16_co_wl2 dp8tvar16_co_bl1 dp8tvar16_co_bl1_n dp8tvar16_co_bl2_n dp8tvar16_co_bl2 DP8TVar16
Xdp8tvar17 vss dp8tvar17_noco_vdd dp8tvar17_noco_wl1 dp8tvar17_noco_wl2 dp8tvar17_noco_bl1 dp8tvar17_noco_bl1_n dp8tvar17_noco_bl2 dp8tvar17_noco_bl2_n dp8tvar17_co_vdd dp8tvar17_co_bit dp8tvar17_co_bit_n dp8tvar17_co_wl1 dp8tvar17_co_wl2 dp8tvar17_co_bl1 dp8tvar17_co_bl1_n dp8tvar17_co_bl2_n dp8tvar17_co_bl2 DP8TVar17
Xdp8tvar18 vss dp8tvar18_noco_vdd dp8tvar18_noco_wl1 dp8tvar18_noco_wl2 dp8tvar18_noco_bl1 dp8tvar18_noco_bl1_n dp8tvar18_noco_bl2 dp8tvar18_noco_bl2_n dp8tvar18_co_vdd dp8tvar18_co_bit dp8tvar18_co_bit_n dp8tvar18_co_wl1 dp8tvar18_co_wl2 dp8tvar18_co_bl1 dp8tvar18_co_bl1_n dp8tvar18_co_bl2_n dp8tvar18_co_bl2 DP8TVar18
Xdp8tvar19 vss dp8tvar19_noco_vdd dp8tvar19_noco_wl1 dp8tvar19_noco_wl2 dp8tvar19_noco_bl1 dp8tvar19_noco_bl1_n dp8tvar19_noco_bl2 dp8tvar19_noco_bl2_n dp8tvar19_co_vdd dp8tvar19_co_bit dp8tvar19_co_bit_n dp8tvar19_co_wl1 dp8tvar19_co_wl2 dp8tvar19_co_bl1 dp8tvar19_co_bl1_n dp8tvar19_co_bl2_n dp8tvar19_co_bl2 DP8TVar19
Xdp8tvar20 vss dp8tvar20_noco_vdd dp8tvar20_noco_wl1 dp8tvar20_noco_wl2 dp8tvar20_noco_bl1 dp8tvar20_noco_bl1_n dp8tvar20_noco_bl2 dp8tvar20_noco_bl2_n dp8tvar20_co_vdd dp8tvar20_co_bit dp8tvar20_co_bit_n dp8tvar20_co_wl1 dp8tvar20_co_wl2 dp8tvar20_co_bl1 dp8tvar20_co_bl1_n dp8tvar20_co_bl2_n dp8tvar20_co_bl2 DP8TVar20
.ends SingleCell_TestStructures

