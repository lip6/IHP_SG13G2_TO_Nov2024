** sch_path: /home/joerdson/ihp130_skel/xschem/chip/CryoChip.sch
.subckt CryoChip GPN SDP1 SDP2 SDP3 SDP4 SDP5 SDN5 SDN4 SDN3 SDN2 SDN1 SDN0 SDP6 SDP0 SDN6 BP BN BN SN1 DN1 GN1 BN SN2 DN2 GN2 BN SN3 DN3 GN3 BN SN4 DN4 GN4 BN SN5 DN5 GN5 BN SN6 DN6 GN6 BN SN7 DN7 GN7 BN SN8
+ DN8 GN8 BP1 SP1 DP1 GP1 BP2 SP2 DP2 GP2 BP3 SP3 DP3 GP3 BP4 SP4 DP4 GP4 BP5 SP5 DP5 GP5 BP6 SP6 DP6 GP6 BP7 SP7 DP7 GP7 BP8 SP8 DP8 GP8 VDD IN OUT BN
M1 SDN0 GPN SDN1 BN sg13_lv_nmos l=0.13u w=0.15u ng=1 m=1
M2 SDP1 GPN SDP0 BP sg13_lv_pmos l=0.13u w=0.15u ng=1 m=1
M3 SDN1 GPN SDN2 BN sg13_lv_nmos l=0.13u w=3.0u ng=1 m=1
M4 SDP2 GPN SDP1 BP sg13_lv_pmos l=0.13u w=3.0u ng=1 m=1
M5 SDN2 GPN SDN3 BN sg13_lv_nmos l=0.3u w=3.0u ng=1 m=1
M6 SDP3 GPN SDP2 BP sg13_lv_pmos l=0.3u w=3.0u ng=1 m=1
M7 SDN3 GPN SDN4 BN sg13_lv_nmos l=0.6u w=3.0u ng=1 m=1
M8 SDP4 GPN SDP3 BP sg13_lv_pmos l=0.6u w=3.0u ng=1 m=1
M9 SDN4 GPN SDN5 BN sg13_lv_nmos l=1.0u w=3.0u ng=1 m=1
M10 SDP5 GPN SDP4 BP sg13_lv_pmos l=1.0u w=3.0u ng=1 m=1
M11 SDN5 GPN SDN6 BN sg13_lv_nmos l=10u w=10u ng=1 m=1
M12 SDP6 GPN SDP5 BP sg13_lv_pmos l=10u w=10u ng=1 m=1
M13 DN1 GN1 SN1 BN sg13_lv_nmos w=0.15u l=0.13u ng=1 m=1
M14 DN2 GN2 SN2 BN sg13_lv_nmos w=3.0u l=0.13u ng=1 m=1
M15 DN3 GN3 SN3 BN sg13_lv_nmos w=3.0u l=0.3u ng=1 m=1
M16 DN4 GN4 SN4 BN sg13_lv_nmos w=3.0u l=0.6u ng=1 m=1
M17 DN5 GN5 SN5 BN sg13_lv_nmos w=3.0u l=1u ng=1 m=1
M18 DN6 GN6 SN6 BN sg13_lv_nmos w=10u l=10u ng=1 m=1
M19 DN7 GN7 SN7 BN sg13_lv_nmos w=1u l=1u ng=1 m=1
M20 DN8 GN8 SN8 BN sg13_lv_nmos w=0.5u l=1u ng=1 m=1
M21 DP1 GP1 SP1 BP1 sg13_lv_pmos w=0.15u l=0.13u ng=1 m=1
M22 DP2 GP2 SP2 BP2 sg13_lv_pmos w=3.0u l=0.13u ng=1 m=1
M23 DP3 GP3 SP3 BP3 sg13_lv_pmos w=3.0u l=0.3u ng=1 m=1
M24 DP4 GP4 SP4 BP4 sg13_lv_pmos w=3.0u l=0.6u ng=1 m=1
M25 DP5 GP5 SP5 BP5 sg13_lv_pmos w=3u l=1u ng=1 m=1
M26 DP6 GP6 SP6 BP6 sg13_lv_pmos w=10u l=10u ng=1 m=1
M27 DP7 GP7 SP7 BP7 sg13_lv_pmos w=1u l=1u ng=1 m=1
M28 DP8 GP8 SP8 BP8 sg13_lv_pmos w=0.5u l=1u ng=1 m=1
M29 BN IN OUT BN sg13_lv_nmos l=0.13u w=0.15u ng=1 m=1
M30 out IN VDD VDD sg13_lv_pmos l=0.13u w=0.6u ng=1 m=1
.ends
.end
