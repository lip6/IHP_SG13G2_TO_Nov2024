module chip_top (aux_enable_pad,
    clk_pad,
    lfsr_out_pad,
    rst_pad,
    shreg_in_pad,
    shreg_out_pad,
    wr_enable_pad,
    data_in_pad,
    data_out_pad,
    out_select_pad,
    reg_addr_pad);
 inout aux_enable_pad;
 inout clk_pad;
 inout lfsr_out_pad;
 inout rst_pad;
 inout shreg_in_pad;
 inout shreg_out_pad;
 inout wr_enable_pad;
 inout [7:0] data_in_pad;
 inout [7:0] data_out_pad;
 inout [1:0] out_select_pad;
 inout [2:0] reg_addr_pad;

 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire _04785_;
 wire _04786_;
 wire _04787_;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04809_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire _04907_;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire _04915_;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire _04927_;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire _04933_;
 wire _04934_;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire _04940_;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire _04952_;
 wire _04953_;
 wire _04954_;
 wire _04955_;
 wire _04956_;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire _04965_;
 wire _04966_;
 wire _04967_;
 wire _04968_;
 wire _04969_;
 wire _04970_;
 wire _04971_;
 wire _04972_;
 wire _04973_;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire _04977_;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire _04982_;
 wire _04983_;
 wire _04984_;
 wire _04985_;
 wire _04986_;
 wire _04987_;
 wire _04988_;
 wire _04989_;
 wire _04990_;
 wire _04991_;
 wire _04992_;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04997_;
 wire _04998_;
 wire _04999_;
 wire _05000_;
 wire _05001_;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire _05012_;
 wire _05013_;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire _05018_;
 wire _05019_;
 wire _05020_;
 wire _05021_;
 wire _05022_;
 wire _05023_;
 wire _05024_;
 wire _05025_;
 wire _05026_;
 wire _05027_;
 wire _05028_;
 wire _05029_;
 wire _05030_;
 wire _05031_;
 wire _05032_;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire _05036_;
 wire _05037_;
 wire _05038_;
 wire _05039_;
 wire _05040_;
 wire _05041_;
 wire _05042_;
 wire _05043_;
 wire _05044_;
 wire _05045_;
 wire _05046_;
 wire _05047_;
 wire _05048_;
 wire _05049_;
 wire _05050_;
 wire _05051_;
 wire _05052_;
 wire _05053_;
 wire _05054_;
 wire _05055_;
 wire _05056_;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire _05061_;
 wire _05062_;
 wire _05063_;
 wire _05064_;
 wire _05065_;
 wire _05066_;
 wire _05067_;
 wire _05068_;
 wire _05069_;
 wire _05070_;
 wire _05071_;
 wire _05072_;
 wire _05073_;
 wire _05074_;
 wire _05075_;
 wire _05076_;
 wire _05077_;
 wire _05078_;
 wire _05079_;
 wire _05080_;
 wire _05081_;
 wire _05082_;
 wire _05083_;
 wire _05084_;
 wire _05085_;
 wire _05086_;
 wire _05087_;
 wire _05088_;
 wire _05089_;
 wire _05090_;
 wire _05091_;
 wire _05092_;
 wire _05093_;
 wire _05094_;
 wire _05095_;
 wire _05096_;
 wire _05097_;
 wire _05098_;
 wire _05099_;
 wire _05100_;
 wire _05101_;
 wire _05102_;
 wire _05103_;
 wire _05104_;
 wire _05105_;
 wire _05106_;
 wire _05107_;
 wire _05108_;
 wire _05109_;
 wire _05110_;
 wire _05111_;
 wire _05112_;
 wire _05113_;
 wire _05114_;
 wire _05115_;
 wire _05116_;
 wire _05117_;
 wire _05118_;
 wire _05119_;
 wire _05120_;
 wire _05121_;
 wire _05122_;
 wire _05123_;
 wire _05124_;
 wire _05125_;
 wire _05126_;
 wire _05127_;
 wire _05128_;
 wire _05129_;
 wire _05130_;
 wire _05131_;
 wire _05132_;
 wire _05133_;
 wire _05134_;
 wire _05135_;
 wire _05136_;
 wire _05137_;
 wire _05138_;
 wire _05139_;
 wire _05140_;
 wire _05141_;
 wire _05142_;
 wire _05143_;
 wire _05144_;
 wire _05145_;
 wire _05146_;
 wire _05147_;
 wire _05148_;
 wire _05149_;
 wire _05150_;
 wire _05151_;
 wire _05152_;
 wire _05153_;
 wire _05154_;
 wire _05155_;
 wire _05156_;
 wire _05157_;
 wire _05158_;
 wire _05159_;
 wire _05160_;
 wire _05161_;
 wire _05162_;
 wire _05163_;
 wire _05164_;
 wire _05165_;
 wire _05166_;
 wire _05167_;
 wire _05168_;
 wire _05169_;
 wire _05170_;
 wire _05171_;
 wire _05172_;
 wire _05173_;
 wire _05174_;
 wire _05175_;
 wire _05176_;
 wire _05177_;
 wire _05178_;
 wire _05179_;
 wire _05180_;
 wire _05181_;
 wire _05182_;
 wire _05183_;
 wire _05184_;
 wire _05185_;
 wire _05186_;
 wire _05187_;
 wire _05188_;
 wire _05189_;
 wire _05190_;
 wire _05191_;
 wire _05192_;
 wire _05193_;
 wire _05194_;
 wire _05195_;
 wire _05196_;
 wire _05197_;
 wire _05198_;
 wire _05199_;
 wire _05200_;
 wire _05201_;
 wire _05202_;
 wire _05203_;
 wire _05204_;
 wire _05205_;
 wire _05206_;
 wire _05207_;
 wire _05208_;
 wire _05209_;
 wire _05210_;
 wire _05211_;
 wire _05212_;
 wire _05213_;
 wire _05214_;
 wire _05215_;
 wire _05216_;
 wire _05217_;
 wire _05218_;
 wire _05219_;
 wire _05220_;
 wire _05221_;
 wire _05222_;
 wire _05223_;
 wire _05224_;
 wire _05225_;
 wire _05226_;
 wire _05227_;
 wire _05228_;
 wire _05229_;
 wire _05230_;
 wire _05231_;
 wire _05232_;
 wire _05233_;
 wire _05234_;
 wire _05235_;
 wire _05236_;
 wire _05237_;
 wire _05238_;
 wire _05239_;
 wire _05240_;
 wire _05241_;
 wire _05242_;
 wire _05243_;
 wire _05244_;
 wire _05245_;
 wire _05246_;
 wire _05247_;
 wire _05248_;
 wire _05249_;
 wire _05250_;
 wire _05251_;
 wire _05252_;
 wire _05253_;
 wire _05254_;
 wire _05255_;
 wire _05256_;
 wire _05257_;
 wire _05258_;
 wire _05259_;
 wire _05260_;
 wire _05261_;
 wire _05262_;
 wire _05263_;
 wire _05264_;
 wire _05265_;
 wire _05266_;
 wire _05267_;
 wire _05268_;
 wire _05269_;
 wire _05270_;
 wire _05271_;
 wire _05272_;
 wire _05273_;
 wire _05274_;
 wire _05275_;
 wire _05276_;
 wire _05277_;
 wire _05278_;
 wire _05279_;
 wire _05280_;
 wire _05281_;
 wire _05282_;
 wire _05283_;
 wire _05284_;
 wire _05285_;
 wire _05286_;
 wire _05287_;
 wire _05288_;
 wire _05289_;
 wire _05290_;
 wire _05291_;
 wire _05292_;
 wire _05293_;
 wire _05294_;
 wire _05295_;
 wire _05296_;
 wire _05297_;
 wire _05298_;
 wire _05299_;
 wire _05300_;
 wire _05301_;
 wire _05302_;
 wire _05303_;
 wire _05304_;
 wire _05305_;
 wire _05306_;
 wire _05307_;
 wire _05308_;
 wire _05309_;
 wire _05310_;
 wire _05311_;
 wire _05312_;
 wire _05313_;
 wire _05314_;
 wire _05315_;
 wire _05316_;
 wire _05317_;
 wire _05318_;
 wire _05319_;
 wire _05320_;
 wire _05321_;
 wire _05322_;
 wire _05323_;
 wire _05324_;
 wire _05325_;
 wire _05326_;
 wire _05327_;
 wire _05328_;
 wire _05329_;
 wire _05330_;
 wire _05331_;
 wire _05332_;
 wire _05333_;
 wire _05334_;
 wire _05335_;
 wire _05336_;
 wire _05337_;
 wire _05338_;
 wire _05339_;
 wire _05340_;
 wire _05341_;
 wire _05342_;
 wire _05343_;
 wire _05344_;
 wire _05345_;
 wire _05346_;
 wire _05347_;
 wire _05348_;
 wire _05349_;
 wire _05350_;
 wire _05351_;
 wire _05352_;
 wire _05353_;
 wire _05354_;
 wire _05355_;
 wire _05356_;
 wire _05357_;
 wire _05358_;
 wire _05359_;
 wire _05360_;
 wire _05361_;
 wire _05362_;
 wire _05363_;
 wire _05364_;
 wire _05365_;
 wire _05366_;
 wire _05367_;
 wire _05368_;
 wire _05369_;
 wire _05370_;
 wire _05371_;
 wire _05372_;
 wire _05373_;
 wire _05374_;
 wire _05375_;
 wire _05376_;
 wire _05377_;
 wire _05378_;
 wire _05379_;
 wire _05380_;
 wire _05381_;
 wire _05382_;
 wire _05383_;
 wire _05384_;
 wire _05385_;
 wire _05386_;
 wire _05387_;
 wire _05388_;
 wire _05389_;
 wire _05390_;
 wire _05391_;
 wire _05392_;
 wire _05393_;
 wire _05394_;
 wire _05395_;
 wire _05396_;
 wire _05397_;
 wire _05398_;
 wire _05399_;
 wire _05400_;
 wire _05401_;
 wire _05402_;
 wire _05403_;
 wire _05404_;
 wire _05405_;
 wire _05406_;
 wire _05407_;
 wire _05408_;
 wire _05409_;
 wire _05410_;
 wire _05411_;
 wire _05412_;
 wire _05413_;
 wire _05414_;
 wire _05415_;
 wire _05416_;
 wire _05417_;
 wire _05418_;
 wire _05419_;
 wire _05420_;
 wire _05421_;
 wire _05422_;
 wire _05423_;
 wire _05424_;
 wire _05425_;
 wire _05426_;
 wire _05427_;
 wire _05428_;
 wire _05429_;
 wire _05430_;
 wire _05431_;
 wire _05432_;
 wire _05433_;
 wire _05434_;
 wire _05435_;
 wire _05436_;
 wire _05437_;
 wire _05438_;
 wire _05439_;
 wire _05440_;
 wire _05441_;
 wire _05442_;
 wire _05443_;
 wire _05444_;
 wire _05445_;
 wire _05446_;
 wire _05447_;
 wire _05448_;
 wire _05449_;
 wire _05450_;
 wire _05451_;
 wire _05452_;
 wire _05453_;
 wire _05454_;
 wire _05455_;
 wire _05456_;
 wire _05457_;
 wire _05458_;
 wire _05459_;
 wire _05460_;
 wire _05461_;
 wire _05462_;
 wire _05463_;
 wire _05464_;
 wire _05465_;
 wire _05466_;
 wire _05467_;
 wire _05468_;
 wire _05469_;
 wire _05470_;
 wire _05471_;
 wire _05472_;
 wire _05473_;
 wire _05474_;
 wire _05475_;
 wire _05476_;
 wire _05477_;
 wire _05478_;
 wire _05479_;
 wire _05480_;
 wire _05481_;
 wire _05482_;
 wire _05483_;
 wire _05484_;
 wire _05485_;
 wire _05486_;
 wire _05487_;
 wire _05488_;
 wire _05489_;
 wire _05490_;
 wire _05491_;
 wire _05492_;
 wire _05493_;
 wire _05494_;
 wire _05495_;
 wire _05496_;
 wire _05497_;
 wire _05498_;
 wire _05499_;
 wire _05500_;
 wire _05501_;
 wire _05502_;
 wire _05503_;
 wire _05504_;
 wire _05505_;
 wire _05506_;
 wire _05507_;
 wire _05508_;
 wire _05509_;
 wire _05510_;
 wire _05511_;
 wire _05512_;
 wire _05513_;
 wire _05514_;
 wire _05515_;
 wire _05516_;
 wire _05517_;
 wire _05518_;
 wire _05519_;
 wire _05520_;
 wire _05521_;
 wire _05522_;
 wire _05523_;
 wire _05524_;
 wire _05525_;
 wire _05526_;
 wire _05527_;
 wire _05528_;
 wire _05529_;
 wire _05530_;
 wire _05531_;
 wire _05532_;
 wire _05533_;
 wire _05534_;
 wire _05535_;
 wire _05536_;
 wire _05537_;
 wire _05538_;
 wire _05539_;
 wire _05540_;
 wire _05541_;
 wire _05542_;
 wire _05543_;
 wire _05544_;
 wire _05545_;
 wire _05546_;
 wire _05547_;
 wire _05548_;
 wire _05549_;
 wire _05550_;
 wire _05551_;
 wire _05552_;
 wire _05553_;
 wire _05554_;
 wire _05555_;
 wire _05556_;
 wire _05557_;
 wire _05558_;
 wire _05559_;
 wire _05560_;
 wire _05561_;
 wire _05562_;
 wire _05563_;
 wire _05564_;
 wire _05565_;
 wire _05566_;
 wire _05567_;
 wire _05568_;
 wire _05569_;
 wire _05570_;
 wire _05571_;
 wire _05572_;
 wire _05573_;
 wire _05574_;
 wire _05575_;
 wire _05576_;
 wire _05577_;
 wire _05578_;
 wire _05579_;
 wire _05580_;
 wire _05581_;
 wire _05582_;
 wire _05583_;
 wire _05584_;
 wire _05585_;
 wire _05586_;
 wire _05587_;
 wire _05588_;
 wire _05589_;
 wire _05590_;
 wire _05591_;
 wire _05592_;
 wire _05593_;
 wire _05594_;
 wire _05595_;
 wire _05596_;
 wire _05597_;
 wire _05598_;
 wire _05599_;
 wire _05600_;
 wire _05601_;
 wire _05602_;
 wire _05603_;
 wire _05604_;
 wire _05605_;
 wire _05606_;
 wire _05607_;
 wire _05608_;
 wire _05609_;
 wire _05610_;
 wire _05611_;
 wire _05612_;
 wire _05613_;
 wire _05614_;
 wire _05615_;
 wire _05616_;
 wire _05617_;
 wire _05618_;
 wire _05619_;
 wire _05620_;
 wire _05621_;
 wire _05622_;
 wire _05623_;
 wire _05624_;
 wire _05625_;
 wire _05626_;
 wire _05627_;
 wire _05628_;
 wire _05629_;
 wire _05630_;
 wire _05631_;
 wire _05632_;
 wire _05633_;
 wire _05634_;
 wire _05635_;
 wire _05636_;
 wire _05637_;
 wire _05638_;
 wire _05639_;
 wire _05640_;
 wire _05641_;
 wire _05642_;
 wire _05643_;
 wire _05644_;
 wire _05645_;
 wire _05646_;
 wire _05647_;
 wire _05648_;
 wire _05649_;
 wire _05650_;
 wire _05651_;
 wire _05652_;
 wire _05653_;
 wire _05654_;
 wire _05655_;
 wire _05656_;
 wire _05657_;
 wire _05658_;
 wire _05659_;
 wire _05660_;
 wire _05661_;
 wire _05662_;
 wire _05663_;
 wire _05664_;
 wire _05665_;
 wire _05666_;
 wire _05667_;
 wire _05668_;
 wire _05669_;
 wire _05670_;
 wire _05671_;
 wire _05672_;
 wire _05673_;
 wire _05674_;
 wire _05675_;
 wire _05676_;
 wire _05677_;
 wire _05678_;
 wire _05679_;
 wire _05680_;
 wire _05681_;
 wire _05682_;
 wire _05683_;
 wire _05684_;
 wire _05685_;
 wire _05686_;
 wire _05687_;
 wire _05688_;
 wire _05689_;
 wire _05690_;
 wire _05691_;
 wire _05692_;
 wire _05693_;
 wire _05694_;
 wire _05695_;
 wire _05696_;
 wire _05697_;
 wire _05698_;
 wire _05699_;
 wire _05700_;
 wire _05701_;
 wire _05702_;
 wire _05703_;
 wire _05704_;
 wire _05705_;
 wire _05706_;
 wire _05707_;
 wire _05708_;
 wire _05709_;
 wire _05710_;
 wire _05711_;
 wire _05712_;
 wire _05713_;
 wire _05714_;
 wire _05715_;
 wire _05716_;
 wire _05717_;
 wire _05718_;
 wire _05719_;
 wire _05720_;
 wire _05721_;
 wire _05722_;
 wire _05723_;
 wire _05724_;
 wire _05725_;
 wire _05726_;
 wire _05727_;
 wire _05728_;
 wire _05729_;
 wire _05730_;
 wire _05731_;
 wire _05732_;
 wire _05733_;
 wire _05734_;
 wire _05735_;
 wire _05736_;
 wire _05737_;
 wire _05738_;
 wire _05739_;
 wire _05740_;
 wire _05741_;
 wire _05742_;
 wire _05743_;
 wire _05744_;
 wire _05745_;
 wire _05746_;
 wire _05747_;
 wire _05748_;
 wire _05749_;
 wire _05750_;
 wire _05751_;
 wire _05752_;
 wire _05753_;
 wire _05754_;
 wire _05755_;
 wire _05756_;
 wire _05757_;
 wire _05758_;
 wire _05759_;
 wire _05760_;
 wire _05761_;
 wire _05762_;
 wire _05763_;
 wire _05764_;
 wire _05765_;
 wire _05766_;
 wire _05767_;
 wire _05768_;
 wire _05769_;
 wire _05770_;
 wire _05771_;
 wire _05772_;
 wire _05773_;
 wire _05774_;
 wire _05775_;
 wire _05776_;
 wire _05777_;
 wire _05778_;
 wire _05779_;
 wire _05780_;
 wire _05781_;
 wire _05782_;
 wire _05783_;
 wire _05784_;
 wire _05785_;
 wire _05786_;
 wire _05787_;
 wire _05788_;
 wire _05789_;
 wire _05790_;
 wire _05791_;
 wire _05792_;
 wire _05793_;
 wire _05794_;
 wire _05795_;
 wire _05796_;
 wire _05797_;
 wire _05798_;
 wire _05799_;
 wire _05800_;
 wire _05801_;
 wire _05802_;
 wire _05803_;
 wire _05804_;
 wire _05805_;
 wire _05806_;
 wire _05807_;
 wire _05808_;
 wire _05809_;
 wire _05810_;
 wire _05811_;
 wire _05812_;
 wire _05813_;
 wire _05814_;
 wire _05815_;
 wire _05816_;
 wire _05817_;
 wire _05818_;
 wire _05819_;
 wire _05820_;
 wire _05821_;
 wire _05822_;
 wire _05823_;
 wire _05824_;
 wire _05825_;
 wire _05826_;
 wire _05827_;
 wire _05828_;
 wire _05829_;
 wire _05830_;
 wire _05831_;
 wire _05832_;
 wire _05833_;
 wire _05834_;
 wire _05835_;
 wire _05836_;
 wire _05837_;
 wire _05838_;
 wire _05839_;
 wire _05840_;
 wire _05841_;
 wire _05842_;
 wire _05843_;
 wire _05844_;
 wire _05845_;
 wire _05846_;
 wire _05847_;
 wire _05848_;
 wire _05849_;
 wire _05850_;
 wire _05851_;
 wire _05852_;
 wire _05853_;
 wire _05854_;
 wire _05855_;
 wire _05856_;
 wire _05857_;
 wire _05858_;
 wire _05859_;
 wire _05860_;
 wire _05861_;
 wire _05862_;
 wire _05863_;
 wire _05864_;
 wire _05865_;
 wire _05866_;
 wire _05867_;
 wire _05868_;
 wire _05869_;
 wire _05870_;
 wire _05871_;
 wire _05872_;
 wire _05873_;
 wire _05874_;
 wire _05875_;
 wire _05876_;
 wire _05877_;
 wire _05878_;
 wire _05879_;
 wire _05880_;
 wire _05881_;
 wire _05882_;
 wire _05883_;
 wire _05884_;
 wire _05885_;
 wire _05886_;
 wire _05887_;
 wire _05888_;
 wire _05889_;
 wire _05890_;
 wire _05891_;
 wire _05892_;
 wire _05893_;
 wire _05894_;
 wire _05895_;
 wire _05896_;
 wire _05897_;
 wire _05898_;
 wire _05899_;
 wire _05900_;
 wire _05901_;
 wire _05902_;
 wire _05903_;
 wire _05904_;
 wire _05905_;
 wire _05906_;
 wire _05907_;
 wire _05908_;
 wire _05909_;
 wire _05910_;
 wire _05911_;
 wire _05912_;
 wire _05913_;
 wire _05914_;
 wire _05915_;
 wire _05916_;
 wire _05917_;
 wire _05918_;
 wire _05919_;
 wire _05920_;
 wire _05921_;
 wire _05922_;
 wire _05923_;
 wire _05924_;
 wire _05925_;
 wire _05926_;
 wire _05927_;
 wire _05928_;
 wire _05929_;
 wire _05930_;
 wire _05931_;
 wire _05932_;
 wire _05933_;
 wire _05934_;
 wire _05935_;
 wire _05936_;
 wire _05937_;
 wire _05938_;
 wire _05939_;
 wire _05940_;
 wire _05941_;
 wire _05942_;
 wire _05943_;
 wire _05944_;
 wire _05945_;
 wire _05946_;
 wire _05947_;
 wire _05948_;
 wire _05949_;
 wire _05950_;
 wire _05951_;
 wire _05952_;
 wire _05953_;
 wire _05954_;
 wire _05955_;
 wire _05956_;
 wire _05957_;
 wire _05958_;
 wire _05959_;
 wire _05960_;
 wire _05961_;
 wire _05962_;
 wire _05963_;
 wire _05964_;
 wire _05965_;
 wire _05966_;
 wire _05967_;
 wire _05968_;
 wire _05969_;
 wire _05970_;
 wire _05971_;
 wire _05972_;
 wire _05973_;
 wire _05974_;
 wire _05975_;
 wire _05976_;
 wire _05977_;
 wire _05978_;
 wire _05979_;
 wire _05980_;
 wire _05981_;
 wire _05982_;
 wire _05983_;
 wire _05984_;
 wire _05985_;
 wire _05986_;
 wire _05987_;
 wire _05988_;
 wire _05989_;
 wire _05990_;
 wire _05991_;
 wire _05992_;
 wire _05993_;
 wire _05994_;
 wire _05995_;
 wire _05996_;
 wire _05997_;
 wire _05998_;
 wire _05999_;
 wire _06000_;
 wire _06001_;
 wire _06002_;
 wire _06003_;
 wire _06004_;
 wire _06005_;
 wire _06006_;
 wire _06007_;
 wire _06008_;
 wire _06009_;
 wire _06010_;
 wire _06011_;
 wire _06012_;
 wire _06013_;
 wire _06014_;
 wire _06015_;
 wire _06016_;
 wire _06017_;
 wire _06018_;
 wire _06019_;
 wire _06020_;
 wire _06021_;
 wire _06022_;
 wire _06023_;
 wire _06024_;
 wire _06025_;
 wire _06026_;
 wire _06027_;
 wire _06028_;
 wire _06029_;
 wire _06030_;
 wire _06031_;
 wire _06032_;
 wire _06033_;
 wire _06034_;
 wire _06035_;
 wire _06036_;
 wire _06037_;
 wire _06038_;
 wire _06039_;
 wire _06040_;
 wire _06041_;
 wire _06042_;
 wire _06043_;
 wire _06044_;
 wire _06045_;
 wire _06046_;
 wire _06047_;
 wire _06048_;
 wire _06049_;
 wire _06050_;
 wire _06051_;
 wire _06052_;
 wire _06053_;
 wire _06054_;
 wire _06055_;
 wire _06056_;
 wire _06057_;
 wire _06058_;
 wire _06059_;
 wire _06060_;
 wire _06061_;
 wire _06062_;
 wire _06063_;
 wire _06064_;
 wire _06065_;
 wire _06066_;
 wire _06067_;
 wire _06068_;
 wire _06069_;
 wire _06070_;
 wire _06071_;
 wire _06072_;
 wire _06073_;
 wire _06074_;
 wire _06075_;
 wire _06076_;
 wire _06077_;
 wire _06078_;
 wire _06079_;
 wire _06080_;
 wire _06081_;
 wire _06082_;
 wire _06083_;
 wire _06084_;
 wire _06085_;
 wire _06086_;
 wire _06087_;
 wire _06088_;
 wire _06089_;
 wire _06090_;
 wire _06091_;
 wire _06092_;
 wire _06093_;
 wire _06094_;
 wire _06095_;
 wire _06096_;
 wire _06097_;
 wire _06098_;
 wire _06099_;
 wire _06100_;
 wire _06101_;
 wire _06102_;
 wire _06103_;
 wire _06104_;
 wire _06105_;
 wire _06106_;
 wire _06107_;
 wire _06108_;
 wire _06109_;
 wire _06110_;
 wire _06111_;
 wire _06112_;
 wire _06113_;
 wire _06114_;
 wire _06115_;
 wire _06116_;
 wire _06117_;
 wire _06118_;
 wire _06119_;
 wire _06120_;
 wire _06121_;
 wire _06122_;
 wire _06123_;
 wire _06124_;
 wire _06125_;
 wire _06126_;
 wire _06127_;
 wire _06128_;
 wire _06129_;
 wire _06130_;
 wire _06131_;
 wire _06132_;
 wire _06133_;
 wire _06134_;
 wire _06135_;
 wire _06136_;
 wire _06137_;
 wire _06138_;
 wire _06139_;
 wire _06140_;
 wire _06141_;
 wire _06142_;
 wire _06143_;
 wire _06144_;
 wire _06145_;
 wire _06146_;
 wire _06147_;
 wire _06148_;
 wire _06149_;
 wire _06150_;
 wire _06151_;
 wire _06152_;
 wire _06153_;
 wire _06154_;
 wire _06155_;
 wire _06156_;
 wire _06157_;
 wire _06158_;
 wire _06159_;
 wire _06160_;
 wire _06161_;
 wire _06162_;
 wire _06163_;
 wire _06164_;
 wire _06165_;
 wire _06166_;
 wire _06167_;
 wire _06168_;
 wire _06169_;
 wire _06170_;
 wire _06171_;
 wire _06172_;
 wire _06173_;
 wire _06174_;
 wire _06175_;
 wire _06176_;
 wire _06177_;
 wire _06178_;
 wire _06179_;
 wire _06180_;
 wire _06181_;
 wire _06182_;
 wire _06183_;
 wire _06184_;
 wire _06185_;
 wire _06186_;
 wire _06187_;
 wire _06188_;
 wire _06189_;
 wire _06190_;
 wire _06191_;
 wire _06192_;
 wire _06193_;
 wire _06194_;
 wire _06195_;
 wire _06196_;
 wire _06197_;
 wire _06198_;
 wire _06199_;
 wire _06200_;
 wire _06201_;
 wire _06202_;
 wire _06203_;
 wire _06204_;
 wire _06205_;
 wire _06206_;
 wire _06207_;
 wire _06208_;
 wire _06209_;
 wire _06210_;
 wire _06211_;
 wire _06212_;
 wire _06213_;
 wire _06214_;
 wire _06215_;
 wire _06216_;
 wire _06217_;
 wire _06218_;
 wire _06219_;
 wire _06220_;
 wire _06221_;
 wire _06222_;
 wire _06223_;
 wire _06224_;
 wire _06225_;
 wire _06226_;
 wire _06227_;
 wire _06228_;
 wire _06229_;
 wire _06230_;
 wire _06231_;
 wire _06232_;
 wire _06233_;
 wire _06234_;
 wire _06235_;
 wire _06236_;
 wire _06237_;
 wire _06238_;
 wire _06239_;
 wire _06240_;
 wire _06241_;
 wire _06242_;
 wire _06243_;
 wire _06244_;
 wire _06245_;
 wire _06246_;
 wire _06247_;
 wire _06248_;
 wire _06249_;
 wire _06250_;
 wire _06251_;
 wire _06252_;
 wire _06253_;
 wire _06254_;
 wire _06255_;
 wire _06256_;
 wire _06257_;
 wire _06258_;
 wire _06259_;
 wire _06260_;
 wire _06261_;
 wire _06262_;
 wire _06263_;
 wire _06264_;
 wire _06265_;
 wire _06266_;
 wire _06267_;
 wire _06268_;
 wire _06269_;
 wire _06270_;
 wire _06271_;
 wire _06272_;
 wire _06273_;
 wire _06274_;
 wire _06275_;
 wire _06276_;
 wire _06277_;
 wire _06278_;
 wire _06279_;
 wire _06280_;
 wire _06281_;
 wire _06282_;
 wire _06283_;
 wire _06284_;
 wire _06285_;
 wire _06286_;
 wire _06287_;
 wire _06288_;
 wire _06289_;
 wire _06290_;
 wire _06291_;
 wire _06292_;
 wire _06293_;
 wire _06294_;
 wire _06295_;
 wire _06296_;
 wire _06297_;
 wire _06298_;
 wire _06299_;
 wire _06300_;
 wire _06301_;
 wire _06302_;
 wire _06303_;
 wire _06304_;
 wire _06305_;
 wire _06306_;
 wire _06307_;
 wire _06308_;
 wire _06309_;
 wire _06310_;
 wire _06311_;
 wire _06312_;
 wire _06313_;
 wire _06314_;
 wire _06315_;
 wire _06316_;
 wire _06317_;
 wire _06318_;
 wire _06319_;
 wire _06320_;
 wire _06321_;
 wire _06322_;
 wire _06323_;
 wire _06324_;
 wire _06325_;
 wire _06326_;
 wire _06327_;
 wire _06328_;
 wire _06329_;
 wire _06330_;
 wire _06331_;
 wire _06332_;
 wire _06333_;
 wire _06334_;
 wire _06335_;
 wire _06336_;
 wire _06337_;
 wire _06338_;
 wire _06339_;
 wire _06340_;
 wire _06341_;
 wire _06342_;
 wire _06343_;
 wire _06344_;
 wire _06345_;
 wire _06346_;
 wire _06347_;
 wire _06348_;
 wire _06349_;
 wire _06350_;
 wire _06351_;
 wire _06352_;
 wire _06353_;
 wire _06354_;
 wire _06355_;
 wire _06356_;
 wire _06357_;
 wire _06358_;
 wire _06359_;
 wire _06360_;
 wire _06361_;
 wire _06362_;
 wire _06363_;
 wire _06364_;
 wire _06365_;
 wire _06366_;
 wire _06367_;
 wire _06368_;
 wire _06369_;
 wire _06370_;
 wire _06371_;
 wire _06372_;
 wire _06373_;
 wire _06374_;
 wire _06375_;
 wire _06376_;
 wire _06377_;
 wire _06378_;
 wire _06379_;
 wire _06380_;
 wire _06381_;
 wire _06382_;
 wire _06383_;
 wire _06384_;
 wire _06385_;
 wire _06386_;
 wire _06387_;
 wire _06388_;
 wire _06389_;
 wire _06390_;
 wire _06391_;
 wire _06392_;
 wire _06393_;
 wire _06394_;
 wire _06395_;
 wire _06396_;
 wire _06397_;
 wire _06398_;
 wire _06399_;
 wire _06400_;
 wire _06401_;
 wire _06402_;
 wire _06403_;
 wire _06404_;
 wire _06405_;
 wire _06406_;
 wire _06407_;
 wire _06408_;
 wire _06409_;
 wire _06410_;
 wire _06411_;
 wire _06412_;
 wire _06413_;
 wire _06414_;
 wire _06415_;
 wire _06416_;
 wire _06417_;
 wire _06418_;
 wire _06419_;
 wire _06420_;
 wire _06421_;
 wire _06422_;
 wire _06423_;
 wire _06424_;
 wire _06425_;
 wire _06426_;
 wire _06427_;
 wire _06428_;
 wire _06429_;
 wire _06430_;
 wire _06431_;
 wire _06432_;
 wire _06433_;
 wire _06434_;
 wire _06435_;
 wire _06436_;
 wire _06437_;
 wire _06438_;
 wire _06439_;
 wire _06440_;
 wire _06441_;
 wire _06442_;
 wire _06443_;
 wire _06444_;
 wire _06445_;
 wire _06446_;
 wire _06447_;
 wire _06448_;
 wire _06449_;
 wire _06450_;
 wire _06451_;
 wire _06452_;
 wire _06453_;
 wire _06454_;
 wire _06455_;
 wire _06456_;
 wire _06457_;
 wire _06458_;
 wire _06459_;
 wire _06460_;
 wire _06461_;
 wire _06462_;
 wire _06463_;
 wire _06464_;
 wire _06465_;
 wire _06466_;
 wire _06467_;
 wire _06468_;
 wire _06469_;
 wire _06470_;
 wire _06471_;
 wire _06472_;
 wire _06473_;
 wire _06474_;
 wire _06475_;
 wire _06476_;
 wire _06477_;
 wire _06478_;
 wire _06479_;
 wire _06480_;
 wire _06481_;
 wire _06482_;
 wire _06483_;
 wire _06484_;
 wire _06485_;
 wire _06486_;
 wire _06487_;
 wire _06488_;
 wire _06489_;
 wire _06490_;
 wire _06491_;
 wire _06492_;
 wire _06493_;
 wire _06494_;
 wire _06495_;
 wire _06496_;
 wire _06497_;
 wire _06498_;
 wire _06499_;
 wire _06500_;
 wire _06501_;
 wire _06502_;
 wire _06503_;
 wire _06504_;
 wire _06505_;
 wire _06506_;
 wire _06507_;
 wire _06508_;
 wire _06509_;
 wire _06510_;
 wire _06511_;
 wire _06512_;
 wire _06513_;
 wire _06514_;
 wire _06515_;
 wire _06516_;
 wire _06517_;
 wire _06518_;
 wire _06519_;
 wire _06520_;
 wire _06521_;
 wire _06522_;
 wire _06523_;
 wire _06524_;
 wire _06525_;
 wire _06526_;
 wire _06527_;
 wire _06528_;
 wire _06529_;
 wire _06530_;
 wire _06531_;
 wire _06532_;
 wire _06533_;
 wire _06534_;
 wire _06535_;
 wire _06536_;
 wire _06537_;
 wire _06538_;
 wire _06539_;
 wire _06540_;
 wire _06541_;
 wire _06542_;
 wire _06543_;
 wire _06544_;
 wire _06545_;
 wire _06546_;
 wire _06547_;
 wire _06548_;
 wire _06549_;
 wire _06550_;
 wire _06551_;
 wire _06552_;
 wire _06553_;
 wire _06554_;
 wire _06555_;
 wire _06556_;
 wire _06557_;
 wire _06558_;
 wire _06559_;
 wire _06560_;
 wire _06561_;
 wire _06562_;
 wire _06563_;
 wire _06564_;
 wire _06565_;
 wire _06566_;
 wire _06567_;
 wire _06568_;
 wire _06569_;
 wire _06570_;
 wire _06571_;
 wire _06572_;
 wire _06573_;
 wire _06574_;
 wire _06575_;
 wire _06576_;
 wire _06577_;
 wire _06578_;
 wire _06579_;
 wire _06580_;
 wire _06581_;
 wire _06582_;
 wire _06583_;
 wire _06584_;
 wire _06585_;
 wire _06586_;
 wire _06587_;
 wire _06588_;
 wire _06589_;
 wire _06590_;
 wire _06591_;
 wire _06592_;
 wire _06593_;
 wire _06594_;
 wire _06595_;
 wire _06596_;
 wire _06597_;
 wire _06598_;
 wire _06599_;
 wire _06600_;
 wire _06601_;
 wire _06602_;
 wire _06603_;
 wire _06604_;
 wire _06605_;
 wire _06606_;
 wire _06607_;
 wire _06608_;
 wire _06609_;
 wire _06610_;
 wire _06611_;
 wire _06612_;
 wire _06613_;
 wire _06614_;
 wire _06615_;
 wire _06616_;
 wire _06617_;
 wire _06618_;
 wire _06619_;
 wire _06620_;
 wire _06621_;
 wire _06622_;
 wire _06623_;
 wire _06624_;
 wire _06625_;
 wire _06626_;
 wire _06627_;
 wire _06628_;
 wire _06629_;
 wire _06630_;
 wire _06631_;
 wire _06632_;
 wire _06633_;
 wire _06634_;
 wire _06635_;
 wire _06636_;
 wire _06637_;
 wire _06638_;
 wire _06639_;
 wire _06640_;
 wire _06641_;
 wire _06642_;
 wire _06643_;
 wire _06644_;
 wire _06645_;
 wire _06646_;
 wire _06647_;
 wire _06648_;
 wire _06649_;
 wire _06650_;
 wire _06651_;
 wire _06652_;
 wire _06653_;
 wire _06654_;
 wire _06655_;
 wire _06656_;
 wire _06657_;
 wire _06658_;
 wire _06659_;
 wire _06660_;
 wire _06661_;
 wire _06662_;
 wire _06663_;
 wire _06664_;
 wire _06665_;
 wire _06666_;
 wire _06667_;
 wire _06668_;
 wire _06669_;
 wire _06670_;
 wire _06671_;
 wire _06672_;
 wire _06673_;
 wire _06674_;
 wire _06675_;
 wire _06676_;
 wire _06677_;
 wire _06678_;
 wire _06679_;
 wire _06680_;
 wire _06681_;
 wire _06682_;
 wire _06683_;
 wire _06684_;
 wire _06685_;
 wire _06686_;
 wire _06687_;
 wire _06688_;
 wire _06689_;
 wire _06690_;
 wire _06691_;
 wire _06692_;
 wire _06693_;
 wire _06694_;
 wire _06695_;
 wire _06696_;
 wire _06697_;
 wire _06698_;
 wire _06699_;
 wire _06700_;
 wire _06701_;
 wire _06702_;
 wire _06703_;
 wire _06704_;
 wire _06705_;
 wire _06706_;
 wire _06707_;
 wire _06708_;
 wire _06709_;
 wire _06710_;
 wire _06711_;
 wire _06712_;
 wire _06713_;
 wire _06714_;
 wire _06715_;
 wire _06716_;
 wire _06717_;
 wire _06718_;
 wire _06719_;
 wire _06720_;
 wire _06721_;
 wire _06722_;
 wire _06723_;
 wire _06724_;
 wire _06725_;
 wire _06726_;
 wire _06727_;
 wire _06728_;
 wire _06729_;
 wire _06730_;
 wire _06731_;
 wire _06732_;
 wire _06733_;
 wire _06734_;
 wire _06735_;
 wire _06736_;
 wire _06737_;
 wire _06738_;
 wire _06739_;
 wire _06740_;
 wire _06741_;
 wire _06742_;
 wire _06743_;
 wire _06744_;
 wire _06745_;
 wire _06746_;
 wire _06747_;
 wire _06748_;
 wire _06749_;
 wire _06750_;
 wire _06751_;
 wire _06752_;
 wire _06753_;
 wire _06754_;
 wire _06755_;
 wire _06756_;
 wire _06757_;
 wire _06758_;
 wire _06759_;
 wire _06760_;
 wire _06761_;
 wire _06762_;
 wire _06763_;
 wire _06764_;
 wire _06765_;
 wire _06766_;
 wire _06767_;
 wire _06768_;
 wire _06769_;
 wire _06770_;
 wire _06771_;
 wire _06772_;
 wire _06773_;
 wire _06774_;
 wire _06775_;
 wire _06776_;
 wire _06777_;
 wire _06778_;
 wire _06779_;
 wire _06780_;
 wire _06781_;
 wire _06782_;
 wire _06783_;
 wire _06784_;
 wire _06785_;
 wire _06786_;
 wire _06787_;
 wire _06788_;
 wire _06789_;
 wire _06790_;
 wire _06791_;
 wire _06792_;
 wire _06793_;
 wire _06794_;
 wire _06795_;
 wire _06796_;
 wire _06797_;
 wire _06798_;
 wire _06799_;
 wire _06800_;
 wire _06801_;
 wire clknet_leaf_0_clk_p2c;
 wire aux_enable_p2c;
 wire clk_p2c;
 wire data_in_p2c_1;
 wire data_in_p2c_2;
 wire data_in_p2c_3;
 wire data_in_p2c_4;
 wire data_in_p2c_5;
 wire data_in_p2c_6;
 wire data_in_p2c_7;
 wire data_in_p2c_8;
 wire lfsr_out_c2p;
 wire \median_processor.rst ;
 wire \median_processor.wr_enable ;
 wire out_select_p2c_1;
 wire out_select_p2c_2;
 wire reg_addr_p2c_1;
 wire reg_addr_p2c_2;
 wire reg_addr_p2c_3;
 wire \shift_storage.shreg_in ;
 wire \shift_storage.shreg_out ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net995;
 wire net996;
 wire net997;
 wire net998;
 wire net999;
 wire net1000;
 wire net1001;
 wire net1002;
 wire net1003;
 wire net1004;
 wire net1005;
 wire net1006;
 wire net1007;
 wire net1008;
 wire net1009;
 wire net1010;
 wire net1011;
 wire net1012;
 wire net1013;
 wire net1014;
 wire net1015;
 wire net1016;
 wire net1017;
 wire net1018;
 wire net1019;
 wire net1020;
 wire net1021;
 wire net1022;
 wire net1023;
 wire net1024;
 wire net1025;
 wire net1026;
 wire net1027;
 wire net1028;
 wire net1029;
 wire net1030;
 wire net1031;
 wire net1032;
 wire net1033;
 wire net1034;
 wire net1035;
 wire net1036;
 wire net1037;
 wire net1038;
 wire net1039;
 wire net1040;
 wire net1041;
 wire net1042;
 wire net1043;
 wire net1044;
 wire net1045;
 wire net1046;
 wire net1047;
 wire net1048;
 wire net1049;
 wire net1050;
 wire net1051;
 wire net1052;
 wire net1053;
 wire net1054;
 wire net1055;
 wire net1056;
 wire net1057;
 wire net1058;
 wire net1059;
 wire net1060;
 wire net1061;
 wire net1062;
 wire net1063;
 wire net1064;
 wire net1065;
 wire net1066;
 wire net1067;
 wire net1068;
 wire net1069;
 wire net1070;
 wire net1071;
 wire net1072;
 wire net1073;
 wire net1074;
 wire net1075;
 wire net1076;
 wire net1077;
 wire net1078;
 wire net1079;
 wire net1080;
 wire net1081;
 wire net1082;
 wire net1083;
 wire net1084;
 wire net1085;
 wire net1086;
 wire net1087;
 wire net1088;
 wire net1089;
 wire net1090;
 wire net1091;
 wire net1092;
 wire net1093;
 wire net1094;
 wire net1095;
 wire net1096;
 wire net1097;
 wire net1098;
 wire net1099;
 wire net1100;
 wire net1101;
 wire net1102;
 wire net1103;
 wire net1104;
 wire net1105;
 wire net1106;
 wire net1107;
 wire net1108;
 wire net1109;
 wire net1110;
 wire net1111;
 wire net1112;
 wire net1113;
 wire net1114;
 wire net1115;
 wire net1116;
 wire net1117;
 wire net1118;
 wire net1119;
 wire net1120;
 wire net1121;
 wire net1122;
 wire net1123;
 wire net1124;
 wire net1125;
 wire net1126;
 wire net1127;
 wire net1128;
 wire net1129;
 wire net1130;
 wire net1131;
 wire net1132;
 wire net1133;
 wire net1134;
 wire net1135;
 wire net1136;
 wire net1137;
 wire net1138;
 wire net1139;
 wire net1140;
 wire net1141;
 wire net1142;
 wire net1143;
 wire net1144;
 wire net1145;
 wire net1146;
 wire net1147;
 wire net1148;
 wire net1149;
 wire net1150;
 wire net1151;
 wire net1152;
 wire net1153;
 wire net1154;
 wire net1155;
 wire net1156;
 wire net1157;
 wire net1158;
 wire net1159;
 wire net1160;
 wire net1161;
 wire net1162;
 wire net1163;
 wire net1164;
 wire net1165;
 wire net1166;
 wire net1167;
 wire net1168;
 wire net1169;
 wire net1170;
 wire net1171;
 wire net1172;
 wire net1173;
 wire net1174;
 wire net1175;
 wire net1176;
 wire net1177;
 wire net1178;
 wire net1179;
 wire net1180;
 wire net1181;
 wire net1182;
 wire net1183;
 wire net1184;
 wire net1185;
 wire net1186;
 wire net1187;
 wire net1188;
 wire net1189;
 wire net1190;
 wire net1191;
 wire net1192;
 wire net1193;
 wire net1194;
 wire net1195;
 wire net1196;
 wire net1197;
 wire net1198;
 wire net1199;
 wire net1200;
 wire net1201;
 wire net1202;
 wire net1203;
 wire net1204;
 wire net1205;
 wire net1206;
 wire net1207;
 wire net1208;
 wire net1209;
 wire net1210;
 wire net1211;
 wire net1212;
 wire net1213;
 wire net1214;
 wire net1215;
 wire net1216;
 wire net1217;
 wire net1218;
 wire net1219;
 wire net1220;
 wire net1221;
 wire net1222;
 wire net1223;
 wire net1224;
 wire net1225;
 wire net1226;
 wire net1227;
 wire net1228;
 wire net1229;
 wire net1230;
 wire net1231;
 wire net1232;
 wire net1233;
 wire net1234;
 wire net1235;
 wire net1236;
 wire net1237;
 wire net1238;
 wire net1239;
 wire net1240;
 wire net1241;
 wire net1242;
 wire net1243;
 wire net1244;
 wire net1245;
 wire net1246;
 wire net1247;
 wire net1248;
 wire net1249;
 wire net1250;
 wire net1251;
 wire net1252;
 wire net1253;
 wire net1254;
 wire net1255;
 wire net1256;
 wire net1257;
 wire net1258;
 wire net1259;
 wire net1260;
 wire net1261;
 wire net1262;
 wire net1263;
 wire net1264;
 wire net1265;
 wire net1266;
 wire net1267;
 wire net1268;
 wire net1269;
 wire net1270;
 wire net1271;
 wire net1272;
 wire net1273;
 wire net1274;
 wire net1275;
 wire net1276;
 wire net1277;
 wire net1278;
 wire net1279;
 wire net1280;
 wire net1281;
 wire net1282;
 wire net1283;
 wire net1284;
 wire net1285;
 wire net1286;
 wire net1287;
 wire net1288;
 wire net1289;
 wire net1290;
 wire net1291;
 wire net1292;
 wire net1293;
 wire net1294;
 wire net1295;
 wire net1296;
 wire net1297;
 wire net1298;
 wire net1299;
 wire net1300;
 wire net1301;
 wire net1302;
 wire net1303;
 wire net1304;
 wire net1305;
 wire net1306;
 wire net1307;
 wire net1308;
 wire net1309;
 wire net1310;
 wire net1311;
 wire net1312;
 wire net1313;
 wire net1314;
 wire net1315;
 wire net1316;
 wire net1317;
 wire net1318;
 wire net1319;
 wire net1320;
 wire net1321;
 wire net1322;
 wire net1323;
 wire net1324;
 wire net1325;
 wire net1326;
 wire net1327;
 wire net1328;
 wire net1329;
 wire net1330;
 wire net1331;
 wire net1332;
 wire net1333;
 wire net1334;
 wire net1335;
 wire net1336;
 wire net1337;
 wire net1338;
 wire net1339;
 wire net1340;
 wire net1341;
 wire net1342;
 wire net1343;
 wire net1344;
 wire net1345;
 wire net1346;
 wire net1347;
 wire net1348;
 wire net1349;
 wire net1350;
 wire net1351;
 wire net1352;
 wire net1353;
 wire net1354;
 wire net1355;
 wire net1356;
 wire net1357;
 wire net1358;
 wire net1359;
 wire net1360;
 wire net1361;
 wire net1362;
 wire net1363;
 wire net1364;
 wire net1365;
 wire net1366;
 wire net1367;
 wire net1368;
 wire net1369;
 wire net1370;
 wire net1371;
 wire net1372;
 wire net1373;
 wire net1374;
 wire net1375;
 wire net1376;
 wire net1377;
 wire net1378;
 wire net1379;
 wire net1380;
 wire net1381;
 wire net1382;
 wire net1383;
 wire net1384;
 wire net1385;
 wire net1386;
 wire net1387;
 wire net1388;
 wire net1389;
 wire net1390;
 wire net1391;
 wire net1392;
 wire net1393;
 wire net1394;
 wire net1395;
 wire net1396;
 wire net1397;
 wire net1398;
 wire net1399;
 wire net1400;
 wire net1401;
 wire net1402;
 wire net1403;
 wire net1404;
 wire net1405;
 wire net1406;
 wire net1407;
 wire net1408;
 wire net1409;
 wire net1410;
 wire net1411;
 wire net1412;
 wire net1413;
 wire net1414;
 wire net1415;
 wire net1416;
 wire net1417;
 wire net1418;
 wire net1419;
 wire net1420;
 wire net1421;
 wire net1422;
 wire net1423;
 wire net1424;
 wire net1425;
 wire net1426;
 wire net1427;
 wire net1428;
 wire net1429;
 wire net1430;
 wire net1431;
 wire net1432;
 wire net1433;
 wire net1434;
 wire net1435;
 wire net1436;
 wire net1437;
 wire net1438;
 wire net1439;
 wire net1440;
 wire net1441;
 wire net1442;
 wire net1443;
 wire net1444;
 wire net1445;
 wire net1446;
 wire net1447;
 wire net1448;
 wire net1449;
 wire net1450;
 wire net1451;
 wire net1452;
 wire net1453;
 wire net1454;
 wire net1455;
 wire net1456;
 wire net1457;
 wire net1458;
 wire net1459;
 wire net1460;
 wire net1461;
 wire net1462;
 wire net1463;
 wire net1464;
 wire net1465;
 wire net1466;
 wire net1467;
 wire net1468;
 wire net1469;
 wire net1470;
 wire net1471;
 wire net1472;
 wire net1473;
 wire net1474;
 wire net1475;
 wire net1476;
 wire net1477;
 wire net1478;
 wire net1479;
 wire net1480;
 wire net1481;
 wire net1482;
 wire net1483;
 wire net1484;
 wire net1485;
 wire net1486;
 wire net1487;
 wire net1488;
 wire net1489;
 wire net1490;
 wire net1491;
 wire net1492;
 wire net1493;
 wire net1494;
 wire net1495;
 wire net1496;
 wire net1497;
 wire net1498;
 wire net1499;
 wire net1500;
 wire net1501;
 wire net1502;
 wire net1503;
 wire net1504;
 wire net1505;
 wire net1506;
 wire net1507;
 wire net1508;
 wire net1509;
 wire net1510;
 wire net1511;
 wire net1512;
 wire net1513;
 wire net1514;
 wire net1515;
 wire net1516;
 wire net1517;
 wire net1518;
 wire net1519;
 wire net1520;
 wire net1521;
 wire net1522;
 wire net1523;
 wire net1524;
 wire net1525;
 wire net1526;
 wire net1527;
 wire net1528;
 wire net1529;
 wire net1530;
 wire net1531;
 wire net1532;
 wire net1533;
 wire net1534;
 wire net1535;
 wire net1536;
 wire net1537;
 wire net1538;
 wire net1539;
 wire net1540;
 wire net1541;
 wire net1542;
 wire net1543;
 wire net1544;
 wire net1545;
 wire net1546;
 wire net1547;
 wire net1548;
 wire net1549;
 wire net1550;
 wire net1551;
 wire net1552;
 wire net1553;
 wire net1554;
 wire net1555;
 wire net1556;
 wire net1557;
 wire net1558;
 wire net1559;
 wire net1560;
 wire net1561;
 wire net1562;
 wire net1563;
 wire net1564;
 wire net1565;
 wire net1566;
 wire net1567;
 wire net1568;
 wire net1569;
 wire net1570;
 wire net1571;
 wire net1572;
 wire net1573;
 wire net1574;
 wire net1575;
 wire net1576;
 wire net1577;
 wire net1578;
 wire net1579;
 wire net1580;
 wire net1581;
 wire net1582;
 wire net1583;
 wire net1584;
 wire net1585;
 wire net1586;
 wire net1587;
 wire net1588;
 wire net1589;
 wire net1590;
 wire net1591;
 wire net1592;
 wire net1593;
 wire net1594;
 wire net1595;
 wire net1596;
 wire net1597;
 wire net1598;
 wire net1599;
 wire net1600;
 wire net1601;
 wire net1602;
 wire net1603;
 wire net1604;
 wire net1605;
 wire net1606;
 wire net1607;
 wire net1608;
 wire net1609;
 wire net1610;
 wire net1611;
 wire net1612;
 wire net1613;
 wire net1614;
 wire net1615;
 wire net1616;
 wire net1617;
 wire net1618;
 wire net1619;
 wire net1620;
 wire net1621;
 wire net1622;
 wire net1623;
 wire net1624;
 wire net1625;
 wire net1626;
 wire net1627;
 wire net1628;
 wire net1629;
 wire net1630;
 wire net1631;
 wire net1632;
 wire net1633;
 wire net1634;
 wire net1635;
 wire net1636;
 wire net1637;
 wire net1638;
 wire net1639;
 wire net1640;
 wire net1641;
 wire net1642;
 wire net1643;
 wire net1644;
 wire net1645;
 wire net1646;
 wire net1647;
 wire net1648;
 wire net1649;
 wire net1650;
 wire net1651;
 wire net1652;
 wire net1653;
 wire net1654;
 wire net1655;
 wire net1656;
 wire net1657;
 wire net1658;
 wire net1659;
 wire net1660;
 wire net1661;
 wire net1662;
 wire net1663;
 wire net1664;
 wire net1665;
 wire net1666;
 wire net1667;
 wire net1668;
 wire net1669;
 wire net1670;
 wire net1671;
 wire net1672;
 wire net1673;
 wire net1674;
 wire net1675;
 wire net1676;
 wire net1677;
 wire net1678;
 wire net1679;
 wire net1680;
 wire net1681;
 wire net1682;
 wire net1683;
 wire net1684;
 wire net1685;
 wire net1686;
 wire net1687;
 wire net1688;
 wire net1689;
 wire net1690;
 wire net1691;
 wire net1692;
 wire net1693;
 wire net1694;
 wire net1695;
 wire net1696;
 wire net1697;
 wire net1698;
 wire net1699;
 wire net1700;
 wire net1701;
 wire net1702;
 wire net1703;
 wire net1704;
 wire net1705;
 wire net1706;
 wire net1707;
 wire net1708;
 wire net1709;
 wire net1710;
 wire net1711;
 wire net1712;
 wire net1713;
 wire net1714;
 wire net1715;
 wire net1716;
 wire net1717;
 wire net1718;
 wire net1719;
 wire net1720;
 wire net1721;
 wire net1722;
 wire net1723;
 wire net1724;
 wire net1725;
 wire net1726;
 wire net1727;
 wire net1728;
 wire net1729;
 wire net1730;
 wire net1731;
 wire net1732;
 wire net1733;
 wire net1734;
 wire net1735;
 wire net1736;
 wire net1737;
 wire net1738;
 wire net1739;
 wire net1740;
 wire net1741;
 wire net1742;
 wire net1743;
 wire net1744;
 wire net1745;
 wire net1746;
 wire net1747;
 wire net1748;
 wire net1749;
 wire net1750;
 wire net1751;
 wire net1752;
 wire net1753;
 wire net1754;
 wire net1755;
 wire net1756;
 wire net1757;
 wire net1758;
 wire net1759;
 wire net1760;
 wire net1761;
 wire net1762;
 wire net1763;
 wire net1764;
 wire net1765;
 wire net1766;
 wire net1767;
 wire net1768;
 wire net1769;
 wire net1770;
 wire net1771;
 wire net1772;
 wire net1773;
 wire net1774;
 wire net1775;
 wire net1776;
 wire net1777;
 wire net1778;
 wire net1779;
 wire net1780;
 wire net1781;
 wire net1782;
 wire net1783;
 wire net1784;
 wire net1785;
 wire net1786;
 wire net1787;
 wire net1788;
 wire net1789;
 wire net1790;
 wire net1791;
 wire net1792;
 wire net1793;
 wire net1794;
 wire net1795;
 wire net1796;
 wire net1797;
 wire net1798;
 wire net1799;
 wire net1800;
 wire net1801;
 wire net1802;
 wire net1803;
 wire net1804;
 wire net1805;
 wire net1806;
 wire net1807;
 wire net1808;
 wire net1809;
 wire net1810;
 wire net1811;
 wire net1812;
 wire net1813;
 wire net1814;
 wire net1815;
 wire net1816;
 wire net1817;
 wire net1818;
 wire net1819;
 wire net1820;
 wire net1821;
 wire net1822;
 wire net1823;
 wire net1824;
 wire net1825;
 wire net1826;
 wire net1827;
 wire net1828;
 wire net1829;
 wire net1830;
 wire net1831;
 wire net1832;
 wire net1833;
 wire net1834;
 wire net1835;
 wire net1836;
 wire net1837;
 wire net1838;
 wire net1839;
 wire net1840;
 wire net1841;
 wire net1842;
 wire net1843;
 wire net1844;
 wire net1845;
 wire net1846;
 wire net1847;
 wire net1848;
 wire net1849;
 wire net1850;
 wire net1851;
 wire net1852;
 wire net1853;
 wire net1854;
 wire net1855;
 wire net1856;
 wire net1857;
 wire net1858;
 wire net1859;
 wire net1860;
 wire net1861;
 wire net1862;
 wire net1863;
 wire net1864;
 wire net1865;
 wire net1866;
 wire net1867;
 wire net1868;
 wire net1869;
 wire net1870;
 wire net1871;
 wire net1872;
 wire net1873;
 wire net1874;
 wire net1875;
 wire net1876;
 wire net1877;
 wire net1878;
 wire net1879;
 wire net1880;
 wire net1881;
 wire net1882;
 wire net1883;
 wire net1884;
 wire net1885;
 wire net1886;
 wire net1887;
 wire net1888;
 wire net1889;
 wire net1890;
 wire net1891;
 wire net1892;
 wire net1893;
 wire net1894;
 wire net1895;
 wire net1896;
 wire net1897;
 wire net1898;
 wire net1899;
 wire net1900;
 wire net1901;
 wire net1902;
 wire net1903;
 wire net1904;
 wire net1905;
 wire net1906;
 wire net1907;
 wire net1908;
 wire net1909;
 wire net1910;
 wire net1911;
 wire net1912;
 wire net1913;
 wire net1914;
 wire net1915;
 wire net1916;
 wire net1917;
 wire net1918;
 wire net1919;
 wire net1920;
 wire net1921;
 wire net1922;
 wire net1923;
 wire net1924;
 wire net1925;
 wire net1926;
 wire net1927;
 wire net1928;
 wire net1929;
 wire net1930;
 wire net1931;
 wire net1932;
 wire net1933;
 wire net1934;
 wire net1935;
 wire net1936;
 wire net1937;
 wire net1938;
 wire net1939;
 wire net1940;
 wire net1941;
 wire net1942;
 wire net1943;
 wire net1944;
 wire net1945;
 wire net1946;
 wire net1947;
 wire net1948;
 wire net1949;
 wire net1950;
 wire net1951;
 wire net1952;
 wire net1953;
 wire net1954;
 wire net1955;
 wire net1956;
 wire net1957;
 wire net1958;
 wire net1959;
 wire net1960;
 wire net1961;
 wire net1962;
 wire net1963;
 wire net1964;
 wire net1965;
 wire net1966;
 wire net1967;
 wire net1968;
 wire net1969;
 wire net1970;
 wire net1971;
 wire net1972;
 wire net1973;
 wire net1974;
 wire net1975;
 wire net1976;
 wire net1977;
 wire net1978;
 wire net1979;
 wire net1980;
 wire net1981;
 wire net1982;
 wire net1983;
 wire net1984;
 wire net1985;
 wire net1986;
 wire net1987;
 wire net1988;
 wire net1989;
 wire net1990;
 wire net1991;
 wire net1992;
 wire net1993;
 wire net1994;
 wire net1995;
 wire net1996;
 wire net1997;
 wire net1998;
 wire net1999;
 wire net2000;
 wire net2001;
 wire net2002;
 wire net2003;
 wire net2004;
 wire net2005;
 wire net2006;
 wire net2007;
 wire net2008;
 wire net2009;
 wire net2010;
 wire net2011;
 wire net2012;
 wire net2013;
 wire net2014;
 wire net2015;
 wire net2016;
 wire net2017;
 wire net2018;
 wire net2019;
 wire net2020;
 wire net2021;
 wire net2022;
 wire net2023;
 wire net2024;
 wire net2025;
 wire net2026;
 wire net2027;
 wire net2028;
 wire net2029;
 wire net2030;
 wire net2031;
 wire net2032;
 wire net2033;
 wire net2034;
 wire net2035;
 wire net2036;
 wire net2037;
 wire net2038;
 wire net2039;
 wire net2040;
 wire net2041;
 wire net2042;
 wire net2043;
 wire net2044;
 wire net2045;
 wire net2046;
 wire net2047;
 wire net2048;
 wire net2049;
 wire net2050;
 wire net2051;
 wire net2052;
 wire net2053;
 wire net2054;
 wire net2055;
 wire net2056;
 wire net2057;
 wire net2058;
 wire net2059;
 wire net2060;
 wire net2061;
 wire net2062;
 wire net2063;
 wire net2064;
 wire net2065;
 wire net2066;
 wire net2067;
 wire net2068;
 wire net2069;
 wire net2070;
 wire net2071;
 wire net2072;
 wire net2073;
 wire net2074;
 wire net2075;
 wire net2076;
 wire net2077;
 wire net2078;
 wire net2079;
 wire net2080;
 wire net2081;
 wire net2082;
 wire net2083;
 wire net2084;
 wire net2085;
 wire net2086;
 wire net2087;
 wire net2088;
 wire net2089;
 wire net2090;
 wire net2091;
 wire net2092;
 wire net2093;
 wire net2094;
 wire net2095;
 wire net2096;
 wire net2097;
 wire net2098;
 wire net2099;
 wire net2100;
 wire net2101;
 wire net2102;
 wire net2103;
 wire net2104;
 wire net2105;
 wire net2106;
 wire net2107;
 wire net2108;
 wire net2109;
 wire net2110;
 wire net2111;
 wire net2112;
 wire net2113;
 wire net2114;
 wire net2115;
 wire net2116;
 wire net2117;
 wire net2118;
 wire net2119;
 wire net2120;
 wire net2121;
 wire net2122;
 wire net2123;
 wire net2124;
 wire net2125;
 wire net2126;
 wire net2127;
 wire net2128;
 wire net2129;
 wire net2130;
 wire net2131;
 wire net2132;
 wire net2133;
 wire net2134;
 wire net2135;
 wire net2136;
 wire net2137;
 wire net2138;
 wire net2139;
 wire net2140;
 wire net2141;
 wire net2142;
 wire net2143;
 wire net2144;
 wire net2145;
 wire net2146;
 wire net2147;
 wire net2148;
 wire net2149;
 wire net2150;
 wire net2151;
 wire net2152;
 wire net2153;
 wire net2154;
 wire net2155;
 wire net2156;
 wire net2157;
 wire net2158;
 wire net2159;
 wire net2160;
 wire net2161;
 wire net2162;
 wire net2163;
 wire net2164;
 wire net2165;
 wire net2166;
 wire net2167;
 wire net2168;
 wire net2169;
 wire net2170;
 wire net2171;
 wire net2172;
 wire net2173;
 wire net2174;
 wire net2175;
 wire net2176;
 wire net2177;
 wire net2178;
 wire net2179;
 wire net2180;
 wire net2181;
 wire net2182;
 wire net2183;
 wire net2184;
 wire net2185;
 wire net2186;
 wire net2187;
 wire net2188;
 wire net2189;
 wire net2190;
 wire net2191;
 wire net2192;
 wire net2193;
 wire net2194;
 wire net2195;
 wire net2196;
 wire net2197;
 wire net2198;
 wire clknet_leaf_1_clk_p2c;
 wire clknet_leaf_2_clk_p2c;
 wire clknet_leaf_3_clk_p2c;
 wire clknet_leaf_4_clk_p2c;
 wire clknet_leaf_5_clk_p2c;
 wire clknet_leaf_6_clk_p2c;
 wire clknet_leaf_7_clk_p2c;
 wire clknet_leaf_8_clk_p2c;
 wire clknet_leaf_9_clk_p2c;
 wire clknet_leaf_10_clk_p2c;
 wire clknet_leaf_11_clk_p2c;
 wire clknet_leaf_12_clk_p2c;
 wire clknet_leaf_13_clk_p2c;
 wire clknet_leaf_14_clk_p2c;
 wire clknet_leaf_15_clk_p2c;
 wire clknet_leaf_16_clk_p2c;
 wire clknet_leaf_17_clk_p2c;
 wire clknet_leaf_18_clk_p2c;
 wire clknet_leaf_19_clk_p2c;
 wire clknet_leaf_20_clk_p2c;
 wire clknet_leaf_21_clk_p2c;
 wire clknet_leaf_22_clk_p2c;
 wire clknet_leaf_23_clk_p2c;
 wire clknet_leaf_24_clk_p2c;
 wire clknet_leaf_25_clk_p2c;
 wire clknet_leaf_26_clk_p2c;
 wire clknet_leaf_27_clk_p2c;
 wire clknet_leaf_28_clk_p2c;
 wire clknet_leaf_29_clk_p2c;
 wire clknet_leaf_30_clk_p2c;
 wire clknet_leaf_31_clk_p2c;
 wire clknet_leaf_32_clk_p2c;
 wire clknet_leaf_33_clk_p2c;
 wire clknet_leaf_34_clk_p2c;
 wire clknet_leaf_35_clk_p2c;
 wire clknet_leaf_36_clk_p2c;
 wire clknet_leaf_37_clk_p2c;
 wire clknet_leaf_38_clk_p2c;
 wire clknet_leaf_39_clk_p2c;
 wire clknet_leaf_40_clk_p2c;
 wire clknet_leaf_41_clk_p2c;
 wire clknet_leaf_42_clk_p2c;
 wire clknet_leaf_43_clk_p2c;
 wire clknet_leaf_44_clk_p2c;
 wire clknet_leaf_45_clk_p2c;
 wire clknet_leaf_46_clk_p2c;
 wire clknet_leaf_47_clk_p2c;
 wire clknet_leaf_48_clk_p2c;
 wire clknet_leaf_49_clk_p2c;
 wire clknet_leaf_50_clk_p2c;
 wire clknet_leaf_51_clk_p2c;
 wire clknet_leaf_52_clk_p2c;
 wire clknet_leaf_53_clk_p2c;
 wire clknet_leaf_54_clk_p2c;
 wire clknet_leaf_55_clk_p2c;
 wire clknet_leaf_56_clk_p2c;
 wire clknet_leaf_57_clk_p2c;
 wire clknet_leaf_58_clk_p2c;
 wire clknet_leaf_59_clk_p2c;
 wire clknet_leaf_60_clk_p2c;
 wire clknet_leaf_61_clk_p2c;
 wire clknet_leaf_62_clk_p2c;
 wire clknet_leaf_63_clk_p2c;
 wire clknet_leaf_64_clk_p2c;
 wire clknet_leaf_65_clk_p2c;
 wire clknet_leaf_66_clk_p2c;
 wire clknet_leaf_67_clk_p2c;
 wire clknet_leaf_68_clk_p2c;
 wire clknet_leaf_69_clk_p2c;
 wire clknet_leaf_70_clk_p2c;
 wire clknet_leaf_71_clk_p2c;
 wire clknet_leaf_72_clk_p2c;
 wire clknet_leaf_73_clk_p2c;
 wire clknet_leaf_74_clk_p2c;
 wire clknet_leaf_75_clk_p2c;
 wire clknet_leaf_76_clk_p2c;
 wire clknet_leaf_77_clk_p2c;
 wire clknet_leaf_78_clk_p2c;
 wire clknet_leaf_79_clk_p2c;
 wire clknet_leaf_80_clk_p2c;
 wire clknet_leaf_81_clk_p2c;
 wire clknet_leaf_82_clk_p2c;
 wire clknet_leaf_83_clk_p2c;
 wire clknet_leaf_84_clk_p2c;
 wire clknet_leaf_85_clk_p2c;
 wire clknet_leaf_86_clk_p2c;
 wire clknet_leaf_87_clk_p2c;
 wire clknet_leaf_88_clk_p2c;
 wire clknet_leaf_89_clk_p2c;
 wire clknet_leaf_90_clk_p2c;
 wire clknet_leaf_91_clk_p2c;
 wire clknet_leaf_92_clk_p2c;
 wire clknet_leaf_93_clk_p2c;
 wire clknet_leaf_94_clk_p2c;
 wire clknet_leaf_95_clk_p2c;
 wire clknet_leaf_96_clk_p2c;
 wire clknet_leaf_97_clk_p2c;
 wire clknet_leaf_98_clk_p2c;
 wire clknet_leaf_99_clk_p2c;
 wire clknet_leaf_100_clk_p2c;
 wire clknet_leaf_101_clk_p2c;
 wire clknet_leaf_102_clk_p2c;
 wire clknet_leaf_103_clk_p2c;
 wire clknet_leaf_104_clk_p2c;
 wire clknet_leaf_105_clk_p2c;
 wire clknet_leaf_106_clk_p2c;
 wire clknet_leaf_107_clk_p2c;
 wire clknet_leaf_108_clk_p2c;
 wire clknet_leaf_109_clk_p2c;
 wire clknet_leaf_110_clk_p2c;
 wire clknet_leaf_111_clk_p2c;
 wire clknet_leaf_112_clk_p2c;
 wire clknet_leaf_113_clk_p2c;
 wire clknet_leaf_114_clk_p2c;
 wire clknet_leaf_115_clk_p2c;
 wire clknet_leaf_116_clk_p2c;
 wire clknet_leaf_117_clk_p2c;
 wire clknet_leaf_118_clk_p2c;
 wire clknet_leaf_119_clk_p2c;
 wire clknet_leaf_120_clk_p2c;
 wire clknet_leaf_121_clk_p2c;
 wire clknet_leaf_122_clk_p2c;
 wire clknet_leaf_123_clk_p2c;
 wire clknet_leaf_124_clk_p2c;
 wire clknet_leaf_125_clk_p2c;
 wire clknet_leaf_126_clk_p2c;
 wire clknet_leaf_127_clk_p2c;
 wire clknet_leaf_128_clk_p2c;
 wire clknet_leaf_129_clk_p2c;
 wire clknet_leaf_130_clk_p2c;
 wire clknet_leaf_131_clk_p2c;
 wire clknet_leaf_132_clk_p2c;
 wire clknet_leaf_133_clk_p2c;
 wire clknet_leaf_134_clk_p2c;
 wire clknet_leaf_135_clk_p2c;
 wire clknet_leaf_136_clk_p2c;
 wire clknet_leaf_137_clk_p2c;
 wire clknet_leaf_138_clk_p2c;
 wire clknet_leaf_139_clk_p2c;
 wire clknet_leaf_140_clk_p2c;
 wire clknet_leaf_141_clk_p2c;
 wire clknet_leaf_142_clk_p2c;
 wire clknet_leaf_143_clk_p2c;
 wire clknet_leaf_144_clk_p2c;
 wire clknet_leaf_145_clk_p2c;
 wire clknet_leaf_146_clk_p2c;
 wire clknet_leaf_147_clk_p2c;
 wire clknet_leaf_148_clk_p2c;
 wire clknet_leaf_149_clk_p2c;
 wire clknet_leaf_150_clk_p2c;
 wire clknet_leaf_151_clk_p2c;
 wire clknet_leaf_152_clk_p2c;
 wire clknet_leaf_153_clk_p2c;
 wire clknet_leaf_154_clk_p2c;
 wire clknet_leaf_155_clk_p2c;
 wire clknet_leaf_156_clk_p2c;
 wire clknet_leaf_157_clk_p2c;
 wire clknet_leaf_158_clk_p2c;
 wire clknet_leaf_159_clk_p2c;
 wire clknet_leaf_160_clk_p2c;
 wire clknet_leaf_161_clk_p2c;
 wire clknet_leaf_162_clk_p2c;
 wire clknet_leaf_163_clk_p2c;
 wire clknet_leaf_164_clk_p2c;
 wire clknet_leaf_165_clk_p2c;
 wire clknet_leaf_166_clk_p2c;
 wire clknet_leaf_167_clk_p2c;
 wire clknet_leaf_168_clk_p2c;
 wire clknet_leaf_169_clk_p2c;
 wire clknet_leaf_170_clk_p2c;
 wire clknet_leaf_171_clk_p2c;
 wire clknet_leaf_172_clk_p2c;
 wire clknet_leaf_173_clk_p2c;
 wire clknet_leaf_174_clk_p2c;
 wire clknet_leaf_175_clk_p2c;
 wire clknet_leaf_176_clk_p2c;
 wire clknet_leaf_177_clk_p2c;
 wire clknet_leaf_178_clk_p2c;
 wire clknet_leaf_179_clk_p2c;
 wire clknet_leaf_180_clk_p2c;
 wire clknet_leaf_181_clk_p2c;
 wire clknet_leaf_182_clk_p2c;
 wire clknet_leaf_183_clk_p2c;
 wire clknet_leaf_184_clk_p2c;
 wire clknet_leaf_185_clk_p2c;
 wire clknet_leaf_186_clk_p2c;
 wire clknet_leaf_187_clk_p2c;
 wire clknet_leaf_188_clk_p2c;
 wire clknet_leaf_189_clk_p2c;
 wire clknet_leaf_190_clk_p2c;
 wire clknet_leaf_191_clk_p2c;
 wire clknet_leaf_192_clk_p2c;
 wire clknet_leaf_193_clk_p2c;
 wire clknet_leaf_194_clk_p2c;
 wire clknet_leaf_195_clk_p2c;
 wire clknet_leaf_196_clk_p2c;
 wire clknet_leaf_197_clk_p2c;
 wire clknet_leaf_198_clk_p2c;
 wire clknet_leaf_199_clk_p2c;
 wire clknet_leaf_200_clk_p2c;
 wire clknet_leaf_201_clk_p2c;
 wire clknet_leaf_202_clk_p2c;
 wire clknet_leaf_203_clk_p2c;
 wire clknet_leaf_204_clk_p2c;
 wire clknet_leaf_205_clk_p2c;
 wire clknet_leaf_206_clk_p2c;
 wire clknet_leaf_207_clk_p2c;
 wire clknet_leaf_208_clk_p2c;
 wire clknet_leaf_209_clk_p2c;
 wire clknet_leaf_210_clk_p2c;
 wire clknet_leaf_211_clk_p2c;
 wire clknet_leaf_212_clk_p2c;
 wire clknet_leaf_213_clk_p2c;
 wire clknet_leaf_214_clk_p2c;
 wire clknet_leaf_215_clk_p2c;
 wire clknet_leaf_216_clk_p2c;
 wire clknet_leaf_217_clk_p2c;
 wire clknet_leaf_218_clk_p2c;
 wire clknet_leaf_219_clk_p2c;
 wire clknet_leaf_220_clk_p2c;
 wire clknet_leaf_221_clk_p2c;
 wire clknet_leaf_222_clk_p2c;
 wire clknet_leaf_223_clk_p2c;
 wire clknet_leaf_224_clk_p2c;
 wire clknet_leaf_225_clk_p2c;
 wire clknet_leaf_226_clk_p2c;
 wire clknet_leaf_227_clk_p2c;
 wire clknet_leaf_228_clk_p2c;
 wire clknet_leaf_229_clk_p2c;
 wire clknet_leaf_230_clk_p2c;
 wire clknet_leaf_231_clk_p2c;
 wire clknet_leaf_232_clk_p2c;
 wire clknet_leaf_233_clk_p2c;
 wire clknet_leaf_234_clk_p2c;
 wire clknet_leaf_235_clk_p2c;
 wire clknet_leaf_236_clk_p2c;
 wire clknet_leaf_237_clk_p2c;
 wire clknet_leaf_238_clk_p2c;
 wire clknet_leaf_239_clk_p2c;
 wire clknet_leaf_240_clk_p2c;
 wire clknet_leaf_241_clk_p2c;
 wire clknet_leaf_242_clk_p2c;
 wire clknet_leaf_243_clk_p2c;
 wire clknet_leaf_244_clk_p2c;
 wire clknet_leaf_245_clk_p2c;
 wire clknet_leaf_246_clk_p2c;
 wire clknet_leaf_247_clk_p2c;
 wire clknet_leaf_248_clk_p2c;
 wire clknet_leaf_249_clk_p2c;
 wire clknet_leaf_250_clk_p2c;
 wire clknet_leaf_251_clk_p2c;
 wire clknet_leaf_252_clk_p2c;
 wire clknet_leaf_253_clk_p2c;
 wire clknet_leaf_254_clk_p2c;
 wire clknet_leaf_255_clk_p2c;
 wire clknet_leaf_256_clk_p2c;
 wire clknet_leaf_257_clk_p2c;
 wire clknet_leaf_258_clk_p2c;
 wire clknet_leaf_259_clk_p2c;
 wire clknet_leaf_260_clk_p2c;
 wire clknet_leaf_261_clk_p2c;
 wire clknet_leaf_262_clk_p2c;
 wire clknet_leaf_263_clk_p2c;
 wire clknet_leaf_264_clk_p2c;
 wire clknet_leaf_265_clk_p2c;
 wire clknet_leaf_266_clk_p2c;
 wire clknet_leaf_267_clk_p2c;
 wire clknet_leaf_268_clk_p2c;
 wire clknet_leaf_269_clk_p2c;
 wire clknet_leaf_270_clk_p2c;
 wire clknet_leaf_271_clk_p2c;
 wire clknet_leaf_272_clk_p2c;
 wire clknet_leaf_273_clk_p2c;
 wire clknet_leaf_274_clk_p2c;
 wire clknet_leaf_275_clk_p2c;
 wire clknet_leaf_276_clk_p2c;
 wire clknet_leaf_277_clk_p2c;
 wire clknet_leaf_278_clk_p2c;
 wire clknet_leaf_279_clk_p2c;
 wire clknet_leaf_280_clk_p2c;
 wire clknet_leaf_281_clk_p2c;
 wire clknet_leaf_282_clk_p2c;
 wire clknet_leaf_283_clk_p2c;
 wire clknet_leaf_284_clk_p2c;
 wire clknet_leaf_285_clk_p2c;
 wire clknet_leaf_286_clk_p2c;
 wire clknet_leaf_287_clk_p2c;
 wire clknet_leaf_288_clk_p2c;
 wire clknet_leaf_289_clk_p2c;
 wire clknet_leaf_290_clk_p2c;
 wire clknet_leaf_291_clk_p2c;
 wire clknet_leaf_292_clk_p2c;
 wire clknet_leaf_293_clk_p2c;
 wire clknet_leaf_294_clk_p2c;
 wire clknet_0_clk_p2c;
 wire clknet_4_0_0_clk_p2c;
 wire clknet_4_1_0_clk_p2c;
 wire clknet_4_2_0_clk_p2c;
 wire clknet_4_3_0_clk_p2c;
 wire clknet_4_4_0_clk_p2c;
 wire clknet_4_5_0_clk_p2c;
 wire clknet_4_6_0_clk_p2c;
 wire clknet_4_7_0_clk_p2c;
 wire clknet_4_8_0_clk_p2c;
 wire clknet_4_9_0_clk_p2c;
 wire clknet_4_10_0_clk_p2c;
 wire clknet_4_11_0_clk_p2c;
 wire clknet_4_12_0_clk_p2c;
 wire clknet_4_13_0_clk_p2c;
 wire clknet_4_14_0_clk_p2c;
 wire clknet_4_15_0_clk_p2c;
 wire clknet_5_0__leaf_clk_p2c;
 wire clknet_5_1__leaf_clk_p2c;
 wire clknet_5_2__leaf_clk_p2c;
 wire clknet_5_3__leaf_clk_p2c;
 wire clknet_5_4__leaf_clk_p2c;
 wire clknet_5_5__leaf_clk_p2c;
 wire clknet_5_6__leaf_clk_p2c;
 wire clknet_5_7__leaf_clk_p2c;
 wire clknet_5_8__leaf_clk_p2c;
 wire clknet_5_9__leaf_clk_p2c;
 wire clknet_5_10__leaf_clk_p2c;
 wire clknet_5_11__leaf_clk_p2c;
 wire clknet_5_12__leaf_clk_p2c;
 wire clknet_5_13__leaf_clk_p2c;
 wire clknet_5_14__leaf_clk_p2c;
 wire clknet_5_15__leaf_clk_p2c;
 wire clknet_5_16__leaf_clk_p2c;
 wire clknet_5_17__leaf_clk_p2c;
 wire clknet_5_18__leaf_clk_p2c;
 wire clknet_5_19__leaf_clk_p2c;
 wire clknet_5_20__leaf_clk_p2c;
 wire clknet_5_21__leaf_clk_p2c;
 wire clknet_5_22__leaf_clk_p2c;
 wire clknet_5_23__leaf_clk_p2c;
 wire clknet_5_24__leaf_clk_p2c;
 wire clknet_5_25__leaf_clk_p2c;
 wire clknet_5_26__leaf_clk_p2c;
 wire clknet_5_27__leaf_clk_p2c;
 wire clknet_5_28__leaf_clk_p2c;
 wire clknet_5_29__leaf_clk_p2c;
 wire clknet_5_30__leaf_clk_p2c;
 wire clknet_5_31__leaf_clk_p2c;
 wire [7:0] data_out_c2p;
 wire [63:0] \median_processor.input_storage ;
 wire [7:0] \median_processor.median_processor.median_out ;
 wire [30:0] \rando_generator.lfsr_reg ;
 wire [1598:0] \shift_storage.storage ;

 sg13g2_buf_1 _06803_ (.A(net480),
    .X(_01703_));
 sg13g2_nand2b_1 _06804_ (.Y(_01704_),
    .B(\median_processor.input_storage [28]),
    .A_N(\median_processor.input_storage [20]));
 sg13g2_nand2_1 _06805_ (.Y(_01705_),
    .A(net471),
    .B(_01704_));
 sg13g2_buf_1 _06806_ (.A(\median_processor.input_storage [22]),
    .X(_01706_));
 sg13g2_buf_1 _06807_ (.A(\median_processor.input_storage [31]),
    .X(_01707_));
 sg13g2_nand2b_1 _06808_ (.Y(_01708_),
    .B(net469),
    .A_N(\median_processor.input_storage [23]));
 sg13g2_nand2_1 _06809_ (.Y(_01709_),
    .A(net470),
    .B(_01708_));
 sg13g2_inv_2 _06810_ (.Y(_01710_),
    .A(\median_processor.input_storage [30]));
 sg13g2_nand2_1 _06811_ (.Y(_01711_),
    .A(_01710_),
    .B(_01708_));
 sg13g2_nor2_1 _06812_ (.A(net471),
    .B(_01704_),
    .Y(_01712_));
 sg13g2_a221oi_1 _06813_ (.B2(_01711_),
    .C1(_01712_),
    .B1(_01709_),
    .A1(\median_processor.input_storage [29]),
    .Y(_01713_),
    .A2(_01705_));
 sg13g2_inv_1 _06814_ (.Y(_01714_),
    .A(\median_processor.input_storage [23]));
 sg13g2_nand3_1 _06815_ (.B(net470),
    .C(_01708_),
    .A(_01710_),
    .Y(_01715_));
 sg13g2_o21ai_1 _06816_ (.B1(_01715_),
    .Y(_01716_),
    .A1(net469),
    .A2(_01714_));
 sg13g2_nor2_1 _06817_ (.A(_01713_),
    .B(_01716_),
    .Y(_01717_));
 sg13g2_inv_1 _06818_ (.Y(_01718_),
    .A(\median_processor.input_storage [19]));
 sg13g2_buf_1 _06819_ (.A(_01718_),
    .X(_01719_));
 sg13g2_nand2b_1 _06820_ (.Y(_01720_),
    .B(\median_processor.input_storage [18]),
    .A_N(\median_processor.input_storage [26]));
 sg13g2_buf_8 _06821_ (.A(\median_processor.input_storage [17]),
    .X(_01721_));
 sg13g2_nand3b_1 _06822_ (.B(net468),
    .C(\median_processor.input_storage [16]),
    .Y(_01722_),
    .A_N(\median_processor.input_storage [24]));
 sg13g2_and3_1 _06823_ (.X(_01723_),
    .A(net396),
    .B(_01720_),
    .C(_01722_));
 sg13g2_and3_1 _06824_ (.X(_01724_),
    .A(\median_processor.input_storage [27]),
    .B(_01720_),
    .C(_01722_));
 sg13g2_buf_1 _06825_ (.A(\median_processor.input_storage [24]),
    .X(_01725_));
 sg13g2_nor2b_1 _06826_ (.A(net467),
    .B_N(\median_processor.input_storage [16]),
    .Y(_01726_));
 sg13g2_inv_2 _06827_ (.Y(_01727_),
    .A(net479));
 sg13g2_o21ai_1 _06828_ (.B1(_01727_),
    .Y(_01728_),
    .A1(net468),
    .A2(_01726_));
 sg13g2_o21ai_1 _06829_ (.B1(_01728_),
    .Y(_01729_),
    .A1(_01723_),
    .A2(_01724_));
 sg13g2_buf_1 _06830_ (.A(\median_processor.input_storage [27]),
    .X(_01730_));
 sg13g2_inv_1 _06831_ (.Y(_01731_),
    .A(\median_processor.input_storage [27]));
 sg13g2_buf_1 _06832_ (.A(\median_processor.input_storage [19]),
    .X(_01732_));
 sg13g2_nand2b_1 _06833_ (.Y(_01733_),
    .B(\median_processor.input_storage [26]),
    .A_N(\median_processor.input_storage [18]));
 sg13g2_a21oi_1 _06834_ (.A1(net465),
    .A2(net464),
    .Y(_01734_),
    .B1(_01733_));
 sg13g2_a21oi_1 _06835_ (.A1(_01730_),
    .A2(net396),
    .Y(_01735_),
    .B1(_01734_));
 sg13g2_xnor2_1 _06836_ (.Y(_01736_),
    .A(\median_processor.input_storage [25]),
    .B(net468));
 sg13g2_nand3_1 _06837_ (.B(_01720_),
    .C(_01733_),
    .A(_01736_),
    .Y(_01737_));
 sg13g2_buf_1 _06838_ (.A(\median_processor.input_storage [16]),
    .X(_01738_));
 sg13g2_nand2b_1 _06839_ (.Y(_01739_),
    .B(net467),
    .A_N(net463));
 sg13g2_xnor2_1 _06840_ (.Y(_01740_),
    .A(\median_processor.input_storage [27]),
    .B(net464));
 sg13g2_nand3b_1 _06841_ (.B(_01739_),
    .C(_01740_),
    .Y(_01741_),
    .A_N(_01726_));
 sg13g2_xor2_1 _06842_ (.B(\median_processor.input_storage [20]),
    .A(\median_processor.input_storage [28]),
    .X(_01742_));
 sg13g2_xor2_1 _06843_ (.B(\median_processor.input_storage [23]),
    .A(\median_processor.input_storage [31]),
    .X(_01743_));
 sg13g2_xor2_1 _06844_ (.B(net480),
    .A(\median_processor.input_storage [29]),
    .X(_01744_));
 sg13g2_xor2_1 _06845_ (.B(\median_processor.input_storage [22]),
    .A(\median_processor.input_storage [30]),
    .X(_01745_));
 sg13g2_nor4_1 _06846_ (.A(_01742_),
    .B(_01743_),
    .C(_01744_),
    .D(_01745_),
    .Y(_01746_));
 sg13g2_o21ai_1 _06847_ (.B1(_01746_),
    .Y(_01747_),
    .A1(_01737_),
    .A2(_01741_));
 sg13g2_a21oi_2 _06848_ (.B1(_01747_),
    .Y(_01748_),
    .A2(_01735_),
    .A1(_01729_));
 sg13g2_nor2_2 _06849_ (.A(_01717_),
    .B(_01748_),
    .Y(_01749_));
 sg13g2_inv_1 _06850_ (.Y(_01750_),
    .A(_01749_));
 sg13g2_inv_1 _06851_ (.Y(_01751_),
    .A(\median_processor.input_storage [6]));
 sg13g2_buf_1 _06852_ (.A(\median_processor.input_storage [3]),
    .X(_01752_));
 sg13g2_nor2b_1 _06853_ (.A(\median_processor.input_storage [18]),
    .B_N(net478),
    .Y(_01753_));
 sg13g2_a21oi_1 _06854_ (.A1(net461),
    .A2(net396),
    .Y(_01754_),
    .B1(_01753_));
 sg13g2_inv_1 _06855_ (.Y(_01755_),
    .A(\median_processor.input_storage [17]));
 sg13g2_nand2b_1 _06856_ (.Y(_01756_),
    .B(\median_processor.input_storage [18]),
    .A_N(net478));
 sg13g2_nand2b_1 _06857_ (.Y(_01757_),
    .B(\median_processor.input_storage [16]),
    .A_N(net484));
 sg13g2_nand3_1 _06858_ (.B(_01756_),
    .C(_01757_),
    .A(_01755_),
    .Y(_01758_));
 sg13g2_nand3b_1 _06859_ (.B(net468),
    .C(\median_processor.input_storage [16]),
    .Y(_01759_),
    .A_N(net484));
 sg13g2_nand3_1 _06860_ (.B(_01756_),
    .C(_01759_),
    .A(\median_processor.input_storage [1]),
    .Y(_01760_));
 sg13g2_nand3_1 _06861_ (.B(_01758_),
    .C(_01760_),
    .A(_01754_),
    .Y(_01761_));
 sg13g2_inv_2 _06862_ (.Y(_01762_),
    .A(\median_processor.input_storage [5]));
 sg13g2_inv_2 _06863_ (.Y(_01763_),
    .A(\median_processor.input_storage [3]));
 sg13g2_inv_1 _06864_ (.Y(_01764_),
    .A(\median_processor.input_storage [4]));
 sg13g2_a221oi_1 _06865_ (.B2(_01763_),
    .C1(_01764_),
    .B1(net464),
    .A1(_01762_),
    .Y(_01765_),
    .A2(net480));
 sg13g2_nand2_1 _06866_ (.Y(_01766_),
    .A(\median_processor.input_storage [1]),
    .B(_01759_));
 sg13g2_a221oi_1 _06867_ (.B2(_01757_),
    .C1(_01753_),
    .B1(_01755_),
    .A1(net461),
    .Y(_01767_),
    .A2(_01718_));
 sg13g2_o21ai_1 _06868_ (.B1(net461),
    .Y(_01768_),
    .A1(net396),
    .A2(_01756_));
 sg13g2_nand2_1 _06869_ (.Y(_01769_),
    .A(net396),
    .B(_01756_));
 sg13g2_a22oi_1 _06870_ (.Y(_01770_),
    .B1(_01768_),
    .B2(_01769_),
    .A2(_01767_),
    .A1(_01766_));
 sg13g2_a21oi_1 _06871_ (.A1(_01762_),
    .A2(net480),
    .Y(_01771_),
    .B1(\median_processor.input_storage [20]));
 sg13g2_inv_1 _06872_ (.Y(_01772_),
    .A(net480));
 sg13g2_nor2b_1 _06873_ (.A(\median_processor.input_storage [20]),
    .B_N(\median_processor.input_storage [4]),
    .Y(_01773_));
 sg13g2_a21oi_1 _06874_ (.A1(_01772_),
    .A2(_01773_),
    .Y(_01774_),
    .B1(\median_processor.input_storage [5]));
 sg13g2_nor2_1 _06875_ (.A(_01772_),
    .B(_01773_),
    .Y(_01775_));
 sg13g2_nor2_1 _06876_ (.A(_01774_),
    .B(_01775_),
    .Y(_01776_));
 sg13g2_a221oi_1 _06877_ (.B2(_01771_),
    .C1(_01776_),
    .B1(_01770_),
    .A1(_01761_),
    .Y(_01777_),
    .A2(_01765_));
 sg13g2_a21oi_1 _06878_ (.A1(net462),
    .A2(_01777_),
    .Y(_01778_),
    .B1(net470));
 sg13g2_nor2b_1 _06879_ (.A(net483),
    .B_N(\median_processor.input_storage [20]),
    .Y(_01779_));
 sg13g2_nor2_1 _06880_ (.A(net480),
    .B(_01779_),
    .Y(_01780_));
 sg13g2_inv_1 _06881_ (.Y(_01781_),
    .A(net482));
 sg13g2_a21oi_1 _06882_ (.A1(net480),
    .A2(_01779_),
    .Y(_01782_),
    .B1(_01781_));
 sg13g2_nor2_1 _06883_ (.A(_01780_),
    .B(_01782_),
    .Y(_01783_));
 sg13g2_nand2b_1 _06884_ (.Y(_01784_),
    .B(\median_processor.input_storage [14]),
    .A_N(\median_processor.input_storage [22]));
 sg13g2_nand2b_1 _06885_ (.Y(_01785_),
    .B(\median_processor.input_storage [10]),
    .A_N(\median_processor.input_storage [18]));
 sg13g2_inv_1 _06886_ (.Y(_01786_),
    .A(\median_processor.input_storage [11]));
 sg13g2_a21oi_1 _06887_ (.A1(\median_processor.input_storage [19]),
    .A2(_01785_),
    .Y(_01787_),
    .B1(_01786_));
 sg13g2_nor2_1 _06888_ (.A(_01781_),
    .B(net480),
    .Y(_01788_));
 sg13g2_inv_1 _06889_ (.Y(_01789_),
    .A(net483));
 sg13g2_o21ai_1 _06890_ (.B1(_01784_),
    .Y(_01790_),
    .A1(_01789_),
    .A2(\median_processor.input_storage [20]));
 sg13g2_nor2_1 _06891_ (.A(\median_processor.input_storage [19]),
    .B(_01785_),
    .Y(_01791_));
 sg13g2_nor4_1 _06892_ (.A(_01787_),
    .B(_01788_),
    .C(_01790_),
    .D(_01791_),
    .Y(_01792_));
 sg13g2_inv_1 _06893_ (.Y(_01793_),
    .A(\median_processor.input_storage [8]));
 sg13g2_a21oi_1 _06894_ (.A1(_01793_),
    .A2(\median_processor.input_storage [16]),
    .Y(_01794_),
    .B1(net468));
 sg13g2_and2_1 _06895_ (.A(\median_processor.input_storage [17]),
    .B(\median_processor.input_storage [16]),
    .X(_01795_));
 sg13g2_nor2b_1 _06896_ (.A(\median_processor.input_storage [10]),
    .B_N(\median_processor.input_storage [18]),
    .Y(_01796_));
 sg13g2_a221oi_1 _06897_ (.B2(_01793_),
    .C1(_01796_),
    .B1(_01795_),
    .A1(_01786_),
    .Y(_01797_),
    .A2(\median_processor.input_storage [19]));
 sg13g2_o21ai_1 _06898_ (.B1(_01797_),
    .Y(_01798_),
    .A1(\median_processor.input_storage [9]),
    .A2(_01794_));
 sg13g2_inv_2 _06899_ (.Y(_01799_),
    .A(\median_processor.input_storage [22]));
 sg13g2_inv_2 _06900_ (.Y(_01800_),
    .A(net481));
 sg13g2_buf_1 _06901_ (.A(\median_processor.input_storage [23]),
    .X(_01801_));
 sg13g2_nand2_1 _06902_ (.Y(_01802_),
    .A(_01800_),
    .B(net460));
 sg13g2_o21ai_1 _06903_ (.B1(_01802_),
    .Y(_01803_),
    .A1(\median_processor.input_storage [14]),
    .A2(_01799_));
 sg13g2_a221oi_1 _06904_ (.B2(_01798_),
    .C1(_01803_),
    .B1(_01792_),
    .A1(_01783_),
    .Y(_01804_),
    .A2(_01784_));
 sg13g2_buf_1 _06905_ (.A(_01804_),
    .X(_01805_));
 sg13g2_nand3_1 _06906_ (.B(_01761_),
    .C(_01765_),
    .A(\median_processor.input_storage [6]),
    .Y(_01806_));
 sg13g2_and2_1 _06907_ (.A(\median_processor.input_storage [6]),
    .B(_01771_),
    .X(_01807_));
 sg13g2_inv_2 _06908_ (.Y(_01808_),
    .A(net472));
 sg13g2_a21oi_1 _06909_ (.A1(_01808_),
    .A2(_01800_),
    .Y(_01809_),
    .B1(net460));
 sg13g2_a221oi_1 _06910_ (.B2(_01770_),
    .C1(_01809_),
    .B1(_01807_),
    .A1(\median_processor.input_storage [6]),
    .Y(_01810_),
    .A2(_01776_));
 sg13g2_nand3b_1 _06911_ (.B(_01806_),
    .C(_01810_),
    .Y(_01811_),
    .A_N(_01805_));
 sg13g2_or3_1 _06912_ (.A(net472),
    .B(_01714_),
    .C(_01805_),
    .X(_01812_));
 sg13g2_o21ai_1 _06913_ (.B1(_01812_),
    .Y(_01813_),
    .A1(_01778_),
    .A2(_01811_));
 sg13g2_inv_2 _06914_ (.Y(_01814_),
    .A(\median_processor.input_storage [58]));
 sg13g2_buf_1 _06915_ (.A(\median_processor.input_storage [18]),
    .X(_01815_));
 sg13g2_nor2_1 _06916_ (.A(_01814_),
    .B(net459),
    .Y(_01816_));
 sg13g2_inv_2 _06917_ (.Y(_01817_),
    .A(\median_processor.input_storage [57]));
 sg13g2_buf_1 _06918_ (.A(\median_processor.input_storage [56]),
    .X(_01818_));
 sg13g2_nand2b_1 _06919_ (.Y(_01819_),
    .B(net457),
    .A_N(net463));
 sg13g2_nand3b_1 _06920_ (.B(net457),
    .C(\median_processor.input_storage [57]),
    .Y(_01820_),
    .A_N(net463));
 sg13g2_a22oi_1 _06921_ (.Y(_01821_),
    .B1(_01820_),
    .B2(net468),
    .A2(_01819_),
    .A1(net458));
 sg13g2_buf_1 _06922_ (.A(\median_processor.input_storage [20]),
    .X(_01822_));
 sg13g2_buf_1 _06923_ (.A(\median_processor.input_storage [61]),
    .X(_01823_));
 sg13g2_nor2b_1 _06924_ (.A(net455),
    .B_N(net471),
    .Y(_01824_));
 sg13g2_buf_1 _06925_ (.A(\median_processor.input_storage [58]),
    .X(_01825_));
 sg13g2_nor2b_1 _06926_ (.A(net454),
    .B_N(net459),
    .Y(_01826_));
 sg13g2_nor2b_1 _06927_ (.A(\median_processor.input_storage [59]),
    .B_N(net464),
    .Y(_01827_));
 sg13g2_nor4_1 _06928_ (.A(net456),
    .B(_01824_),
    .C(_01826_),
    .D(_01827_),
    .Y(_01828_));
 sg13g2_o21ai_1 _06929_ (.B1(_01828_),
    .Y(_01829_),
    .A1(_01816_),
    .A2(_01821_));
 sg13g2_inv_1 _06930_ (.Y(_01830_),
    .A(\median_processor.input_storage [60]));
 sg13g2_nor4_1 _06931_ (.A(_01830_),
    .B(_01824_),
    .C(_01826_),
    .D(_01827_),
    .Y(_01831_));
 sg13g2_o21ai_1 _06932_ (.B1(_01831_),
    .Y(_01832_),
    .A1(_01816_),
    .A2(_01821_));
 sg13g2_inv_2 _06933_ (.Y(_01833_),
    .A(net455));
 sg13g2_buf_1 _06934_ (.A(\median_processor.input_storage [59]),
    .X(_01834_));
 sg13g2_nand2b_1 _06935_ (.Y(_01835_),
    .B(net453),
    .A_N(net464));
 sg13g2_a221oi_1 _06936_ (.B2(_01830_),
    .C1(_01835_),
    .B1(net456),
    .A1(net395),
    .Y(_01836_),
    .A2(net471));
 sg13g2_nor3_1 _06937_ (.A(_01830_),
    .B(net456),
    .C(_01824_),
    .Y(_01837_));
 sg13g2_nor2_1 _06938_ (.A(_01836_),
    .B(_01837_),
    .Y(_01838_));
 sg13g2_nor2b_1 _06939_ (.A(net460),
    .B_N(net473),
    .Y(_01839_));
 sg13g2_a21oi_1 _06940_ (.A1(net455),
    .A2(_01772_),
    .Y(_01840_),
    .B1(_01839_));
 sg13g2_and2_1 _06941_ (.A(net470),
    .B(_01840_),
    .X(_01841_));
 sg13g2_nand4_1 _06942_ (.B(_01832_),
    .C(_01838_),
    .A(_01829_),
    .Y(_01842_),
    .D(_01841_));
 sg13g2_buf_1 _06943_ (.A(\median_processor.input_storage [62]),
    .X(_01843_));
 sg13g2_nor2b_1 _06944_ (.A(net452),
    .B_N(_01840_),
    .Y(_01844_));
 sg13g2_nand4_1 _06945_ (.B(_01832_),
    .C(_01838_),
    .A(_01829_),
    .Y(_01845_),
    .D(_01844_));
 sg13g2_inv_1 _06946_ (.Y(_01846_),
    .A(net473));
 sg13g2_buf_1 _06947_ (.A(_01846_),
    .X(_01847_));
 sg13g2_buf_1 _06948_ (.A(net460),
    .X(_01848_));
 sg13g2_nor3_1 _06949_ (.A(net452),
    .B(_01799_),
    .C(_01839_),
    .Y(_01849_));
 sg13g2_a21oi_1 _06950_ (.A1(net394),
    .A2(net393),
    .Y(_01850_),
    .B1(_01849_));
 sg13g2_nand3_1 _06951_ (.B(_01845_),
    .C(_01850_),
    .A(_01842_),
    .Y(_01851_));
 sg13g2_buf_1 _06952_ (.A(_01851_),
    .X(_01852_));
 sg13g2_buf_1 _06953_ (.A(\median_processor.input_storage [51]),
    .X(_01853_));
 sg13g2_xor2_1 _06954_ (.B(net464),
    .A(net451),
    .X(_01854_));
 sg13g2_buf_1 _06955_ (.A(\median_processor.input_storage [52]),
    .X(_01855_));
 sg13g2_nand2b_1 _06956_ (.Y(_01856_),
    .B(net450),
    .A_N(net456));
 sg13g2_buf_1 _06957_ (.A(\median_processor.input_storage [53]),
    .X(_01857_));
 sg13g2_nand2b_1 _06958_ (.Y(_01858_),
    .B(net449),
    .A_N(\median_processor.input_storage [21]));
 sg13g2_buf_1 _06959_ (.A(\median_processor.input_storage [48]),
    .X(_01859_));
 sg13g2_xnor2_1 _06960_ (.Y(_01860_),
    .A(net448),
    .B(net463));
 sg13g2_xnor2_1 _06961_ (.Y(_01861_),
    .A(\median_processor.input_storage [50]),
    .B(\median_processor.input_storage [18]));
 sg13g2_nand4_1 _06962_ (.B(_01858_),
    .C(_01860_),
    .A(_01856_),
    .Y(_01862_),
    .D(_01861_));
 sg13g2_buf_1 _06963_ (.A(\median_processor.input_storage [54]),
    .X(_01863_));
 sg13g2_nand2b_1 _06964_ (.Y(_01864_),
    .B(net447),
    .A_N(net470));
 sg13g2_inv_2 _06965_ (.Y(_01865_),
    .A(\median_processor.input_storage [54]));
 sg13g2_nand2_1 _06966_ (.Y(_01866_),
    .A(_01865_),
    .B(net470));
 sg13g2_inv_1 _06967_ (.Y(_01867_),
    .A(\median_processor.input_storage [55]));
 sg13g2_nand2_1 _06968_ (.Y(_01868_),
    .A(net446),
    .B(net460));
 sg13g2_inv_2 _06969_ (.Y(_01869_),
    .A(net449));
 sg13g2_a22oi_1 _06970_ (.Y(_01870_),
    .B1(net471),
    .B2(_01869_),
    .A2(_01714_),
    .A1(\median_processor.input_storage [55]));
 sg13g2_nand4_1 _06971_ (.B(_01866_),
    .C(_01868_),
    .A(_01864_),
    .Y(_01871_),
    .D(_01870_));
 sg13g2_inv_1 _06972_ (.Y(_01872_),
    .A(net456));
 sg13g2_xnor2_1 _06973_ (.Y(_01873_),
    .A(net474),
    .B(net468));
 sg13g2_o21ai_1 _06974_ (.B1(_01873_),
    .Y(_01874_),
    .A1(net450),
    .A2(_01872_));
 sg13g2_or4_1 _06975_ (.A(_01854_),
    .B(_01862_),
    .C(_01871_),
    .D(_01874_),
    .X(_01875_));
 sg13g2_inv_1 _06976_ (.Y(_01876_),
    .A(net448));
 sg13g2_nand2_1 _06977_ (.Y(_01877_),
    .A(_01876_),
    .B(net463));
 sg13g2_nand2b_1 _06978_ (.Y(_01878_),
    .B(net451),
    .A_N(net464));
 sg13g2_nand2_1 _06979_ (.Y(_01879_),
    .A(net459),
    .B(_01878_));
 sg13g2_inv_1 _06980_ (.Y(_01880_),
    .A(\median_processor.input_storage [50]));
 sg13g2_nand2_1 _06981_ (.Y(_01881_),
    .A(_01880_),
    .B(_01878_));
 sg13g2_inv_2 _06982_ (.Y(_01882_),
    .A(net474));
 sg13g2_a21oi_1 _06983_ (.A1(_01876_),
    .A2(_01795_),
    .Y(_01883_),
    .B1(_01882_));
 sg13g2_a221oi_1 _06984_ (.B2(_01881_),
    .C1(_01883_),
    .B1(_01879_),
    .A1(_01755_),
    .Y(_01884_),
    .A2(_01877_));
 sg13g2_nand3_1 _06985_ (.B(net459),
    .C(_01878_),
    .A(_01880_),
    .Y(_01885_));
 sg13g2_o21ai_1 _06986_ (.B1(_01885_),
    .Y(_01886_),
    .A1(net451),
    .A2(net396));
 sg13g2_nand2_1 _06987_ (.Y(_01887_),
    .A(net460),
    .B(_01864_));
 sg13g2_o21ai_1 _06988_ (.B1(net446),
    .Y(_01888_),
    .A1(net460),
    .A2(_01864_));
 sg13g2_nand2_1 _06989_ (.Y(_01889_),
    .A(_01856_),
    .B(_01858_));
 sg13g2_a21oi_1 _06990_ (.A1(_01887_),
    .A2(_01888_),
    .Y(_01890_),
    .B1(_01889_));
 sg13g2_o21ai_1 _06991_ (.B1(_01890_),
    .Y(_01891_),
    .A1(_01884_),
    .A2(_01886_));
 sg13g2_nor3_1 _06992_ (.A(net450),
    .B(_01872_),
    .C(_01889_),
    .Y(_01892_));
 sg13g2_nand2_1 _06993_ (.Y(_01893_),
    .A(_01887_),
    .B(_01888_));
 sg13g2_o21ai_1 _06994_ (.B1(_01893_),
    .Y(_01894_),
    .A1(_01871_),
    .A2(_01892_));
 sg13g2_nand3_1 _06995_ (.B(_01891_),
    .C(_01894_),
    .A(_01875_),
    .Y(_01895_));
 sg13g2_buf_1 _06996_ (.A(_01895_),
    .X(_01896_));
 sg13g2_buf_1 _06997_ (.A(\median_processor.input_storage [38]),
    .X(_01897_));
 sg13g2_nand2b_1 _06998_ (.Y(_01898_),
    .B(net445),
    .A_N(net470));
 sg13g2_nor2_1 _06999_ (.A(net460),
    .B(_01898_),
    .Y(_01899_));
 sg13g2_buf_1 _07000_ (.A(\median_processor.input_storage [39]),
    .X(_01900_));
 sg13g2_inv_2 _07001_ (.Y(_01901_),
    .A(net444));
 sg13g2_buf_1 _07002_ (.A(_01901_),
    .X(_01902_));
 sg13g2_a21oi_1 _07003_ (.A1(_01801_),
    .A2(_01898_),
    .Y(_01903_),
    .B1(net222));
 sg13g2_inv_1 _07004_ (.Y(_01904_),
    .A(net476));
 sg13g2_nand2b_1 _07005_ (.Y(_01905_),
    .B(\median_processor.input_storage [36]),
    .A_N(net456));
 sg13g2_o21ai_1 _07006_ (.B1(_01905_),
    .Y(_01906_),
    .A1(net443),
    .A2(net471));
 sg13g2_inv_1 _07007_ (.Y(_01907_),
    .A(net477));
 sg13g2_inv_1 _07008_ (.Y(_01908_),
    .A(\median_processor.input_storage [33]));
 sg13g2_a21o_1 _07009_ (.A2(_01795_),
    .A1(_01907_),
    .B1(_01908_),
    .X(_01909_));
 sg13g2_buf_1 _07010_ (.A(\median_processor.input_storage [35]),
    .X(_01910_));
 sg13g2_nand2b_1 _07011_ (.Y(_01911_),
    .B(net463),
    .A_N(net477));
 sg13g2_buf_1 _07012_ (.A(\median_processor.input_storage [34]),
    .X(_01912_));
 sg13g2_nor2b_1 _07013_ (.A(net459),
    .B_N(net441),
    .Y(_01913_));
 sg13g2_a221oi_1 _07014_ (.B2(_01911_),
    .C1(_01913_),
    .B1(_01755_),
    .A1(net442),
    .Y(_01914_),
    .A2(net396));
 sg13g2_nand2b_1 _07015_ (.Y(_01915_),
    .B(net459),
    .A_N(net441));
 sg13g2_o21ai_1 _07016_ (.B1(_01719_),
    .Y(_01916_),
    .A1(net442),
    .A2(_01915_));
 sg13g2_nand2_1 _07017_ (.Y(_01917_),
    .A(net442),
    .B(_01915_));
 sg13g2_nor2b_1 _07018_ (.A(\median_processor.input_storage [36]),
    .B_N(net456),
    .Y(_01918_));
 sg13g2_a221oi_1 _07019_ (.B2(_01917_),
    .C1(_01918_),
    .B1(_01916_),
    .A1(_01909_),
    .Y(_01919_),
    .A2(_01914_));
 sg13g2_nor4_2 _07020_ (.A(_01899_),
    .B(_01903_),
    .C(_01906_),
    .Y(_01920_),
    .D(_01919_));
 sg13g2_nor2_1 _07021_ (.A(_01899_),
    .B(_01903_),
    .Y(_01921_));
 sg13g2_nand2b_1 _07022_ (.Y(_01922_),
    .B(_01915_),
    .A_N(_01913_));
 sg13g2_nand2b_1 _07023_ (.Y(_01923_),
    .B(net477),
    .A_N(net463));
 sg13g2_xnor2_1 _07024_ (.Y(_01924_),
    .A(\median_processor.input_storage [35]),
    .B(_01732_));
 sg13g2_nand3_1 _07025_ (.B(_01923_),
    .C(_01924_),
    .A(_01911_),
    .Y(_01925_));
 sg13g2_xnor2_1 _07026_ (.Y(_01926_),
    .A(\median_processor.input_storage [33]),
    .B(_01721_));
 sg13g2_nand2b_1 _07027_ (.Y(_01927_),
    .B(_01926_),
    .A_N(_01918_));
 sg13g2_nor4_1 _07028_ (.A(_01906_),
    .B(_01922_),
    .C(_01925_),
    .D(_01927_),
    .Y(_01928_));
 sg13g2_inv_1 _07029_ (.Y(_01929_),
    .A(net445));
 sg13g2_nand2_1 _07030_ (.Y(_01930_),
    .A(net392),
    .B(_01799_));
 sg13g2_nand2_1 _07031_ (.Y(_01931_),
    .A(net445),
    .B(_01706_));
 sg13g2_xor2_1 _07032_ (.B(_01801_),
    .A(net444),
    .X(_01932_));
 sg13g2_a221oi_1 _07033_ (.B2(_01931_),
    .C1(_01932_),
    .B1(_01930_),
    .A1(net443),
    .Y(_01933_),
    .A2(net471));
 sg13g2_mux2_1 _07034_ (.A0(_01921_),
    .A1(_01928_),
    .S(_01933_),
    .X(_01934_));
 sg13g2_or2_2 _07035_ (.X(_01935_),
    .B(_01934_),
    .A(_01920_));
 sg13g2_nor3_1 _07036_ (.A(net25),
    .B(net24),
    .C(_01935_),
    .Y(_01936_));
 sg13g2_a21oi_1 _07037_ (.A1(net25),
    .A2(net24),
    .Y(_01937_),
    .B1(_01936_));
 sg13g2_and2_1 _07038_ (.A(_01851_),
    .B(_01935_),
    .X(_01938_));
 sg13g2_nand2_1 _07039_ (.Y(_01939_),
    .A(net24),
    .B(_01938_));
 sg13g2_nor2_1 _07040_ (.A(_01813_),
    .B(_01939_),
    .Y(_01940_));
 sg13g2_a21oi_1 _07041_ (.A1(_01813_),
    .A2(_01937_),
    .Y(_01941_),
    .B1(_01940_));
 sg13g2_and3_1 _07042_ (.X(_01942_),
    .A(_01750_),
    .B(net25),
    .C(net24));
 sg13g2_nor2_2 _07043_ (.A(_01920_),
    .B(_01934_),
    .Y(_01943_));
 sg13g2_buf_1 _07044_ (.A(_01808_),
    .X(_01944_));
 sg13g2_inv_1 _07045_ (.Y(_01945_),
    .A(net28));
 sg13g2_buf_1 _07046_ (.A(\median_processor.input_storage [6]),
    .X(_01946_));
 sg13g2_nand2_1 _07047_ (.Y(_01947_),
    .A(net440),
    .B(_01799_));
 sg13g2_nor2_1 _07048_ (.A(net440),
    .B(_01799_),
    .Y(_01948_));
 sg13g2_a21o_1 _07049_ (.A2(_01947_),
    .A1(_01777_),
    .B1(_01948_),
    .X(_01949_));
 sg13g2_nor3_2 _07050_ (.A(net391),
    .B(_01945_),
    .C(_01949_),
    .Y(_01950_));
 sg13g2_a221oi_1 _07051_ (.B2(net391),
    .C1(net393),
    .B1(_01949_),
    .A1(_01800_),
    .Y(_01951_),
    .A2(_01945_));
 sg13g2_or3_1 _07052_ (.A(_01813_),
    .B(_01950_),
    .C(_01951_),
    .X(_01952_));
 sg13g2_nor2_1 _07053_ (.A(_01778_),
    .B(_01811_),
    .Y(_01953_));
 sg13g2_nor2b_1 _07054_ (.A(_01953_),
    .B_N(_01812_),
    .Y(_01954_));
 sg13g2_o21ai_1 _07055_ (.B1(_01954_),
    .Y(_01955_),
    .A1(_01943_),
    .A2(_01952_));
 sg13g2_nor4_2 _07056_ (.A(_01750_),
    .B(_01813_),
    .C(_01950_),
    .Y(_01956_),
    .D(_01951_));
 sg13g2_or2_1 _07057_ (.X(_01957_),
    .B(_01956_),
    .A(_01813_));
 sg13g2_xnor2_1 _07058_ (.Y(_01958_),
    .A(net25),
    .B(_01943_));
 sg13g2_mux2_1 _07059_ (.A0(_01938_),
    .A1(_01958_),
    .S(net24),
    .X(_01959_));
 sg13g2_a22oi_1 _07060_ (.Y(_01960_),
    .B1(_01957_),
    .B2(_01959_),
    .A2(_01955_),
    .A1(_01942_));
 sg13g2_o21ai_1 _07061_ (.B1(_01960_),
    .Y(_01961_),
    .A1(_01750_),
    .A2(_01941_));
 sg13g2_inv_1 _07062_ (.Y(_01962_),
    .A(\median_processor.input_storage [47]));
 sg13g2_nor2_1 _07063_ (.A(\median_processor.input_storage [45]),
    .B(\median_processor.input_storage [44]),
    .Y(_01963_));
 sg13g2_a21oi_1 _07064_ (.A1(_01822_),
    .A2(_01963_),
    .Y(_01964_),
    .B1(_01706_));
 sg13g2_inv_2 _07065_ (.Y(_01965_),
    .A(\median_processor.input_storage [46]));
 sg13g2_a21oi_1 _07066_ (.A1(_01822_),
    .A2(_01963_),
    .Y(_01966_),
    .B1(_01965_));
 sg13g2_buf_1 _07067_ (.A(\median_processor.input_storage [44]),
    .X(_01967_));
 sg13g2_buf_1 _07068_ (.A(\median_processor.input_storage [45]),
    .X(_01968_));
 sg13g2_o21ai_1 _07069_ (.B1(net437),
    .Y(_01969_),
    .A1(_01872_),
    .A2(net438));
 sg13g2_nand2_1 _07070_ (.Y(_01970_),
    .A(_01703_),
    .B(_01969_));
 sg13g2_o21ai_1 _07071_ (.B1(_01970_),
    .Y(_01971_),
    .A1(_01964_),
    .A2(_01966_));
 sg13g2_buf_1 _07072_ (.A(\median_processor.input_storage [46]),
    .X(_01972_));
 sg13g2_nor2b_1 _07073_ (.A(_01848_),
    .B_N(\median_processor.input_storage [47]),
    .Y(_01973_));
 sg13g2_a21oi_1 _07074_ (.A1(_01799_),
    .A2(net436),
    .Y(_01974_),
    .B1(_01973_));
 sg13g2_nand2_1 _07075_ (.Y(_01975_),
    .A(net475),
    .B(\median_processor.input_storage [40]));
 sg13g2_o21ai_1 _07076_ (.B1(_01721_),
    .Y(_01976_),
    .A1(_01738_),
    .A2(_01975_));
 sg13g2_inv_2 _07077_ (.Y(_01977_),
    .A(\median_processor.input_storage [43]));
 sg13g2_buf_1 _07078_ (.A(\median_processor.input_storage [42]),
    .X(_01978_));
 sg13g2_inv_1 _07079_ (.Y(_01979_),
    .A(net435));
 sg13g2_inv_1 _07080_ (.Y(_01980_),
    .A(_01738_));
 sg13g2_buf_1 _07081_ (.A(\median_processor.input_storage [40]),
    .X(_01981_));
 sg13g2_a21oi_1 _07082_ (.A1(_01980_),
    .A2(net434),
    .Y(_01982_),
    .B1(net475));
 sg13g2_a221oi_1 _07083_ (.B2(net459),
    .C1(_01982_),
    .B1(_01979_),
    .A1(_01732_),
    .Y(_01983_),
    .A2(_01977_));
 sg13g2_buf_1 _07084_ (.A(\median_processor.input_storage [43]),
    .X(_01984_));
 sg13g2_nor2b_1 _07085_ (.A(_01815_),
    .B_N(net435),
    .Y(_01985_));
 sg13g2_o21ai_1 _07086_ (.B1(_01719_),
    .Y(_01986_),
    .A1(net433),
    .A2(_01985_));
 sg13g2_nand2_1 _07087_ (.Y(_01987_),
    .A(net433),
    .B(_01985_));
 sg13g2_nor2b_1 _07088_ (.A(_01703_),
    .B_N(net437),
    .Y(_01988_));
 sg13g2_a221oi_1 _07089_ (.B2(net436),
    .C1(_01973_),
    .B1(_01988_),
    .A1(_01872_),
    .Y(_01989_),
    .A2(net438));
 sg13g2_o21ai_1 _07090_ (.B1(_01799_),
    .Y(_01990_),
    .A1(net436),
    .A2(_01988_));
 sg13g2_nand4_1 _07091_ (.B(_01987_),
    .C(_01989_),
    .A(_01986_),
    .Y(_01991_),
    .D(_01990_));
 sg13g2_a21oi_1 _07092_ (.A1(_01976_),
    .A2(_01983_),
    .Y(_01992_),
    .B1(_01991_));
 sg13g2_a221oi_1 _07093_ (.B2(_01974_),
    .C1(_01992_),
    .B1(_01971_),
    .A1(_01848_),
    .Y(_01993_),
    .A2(net439));
 sg13g2_buf_2 _07094_ (.A(_01993_),
    .X(_01994_));
 sg13g2_xor2_1 _07095_ (.B(_01895_),
    .A(_01749_),
    .X(_01995_));
 sg13g2_xnor2_1 _07096_ (.Y(_01996_),
    .A(_01952_),
    .B(_01995_));
 sg13g2_xnor2_1 _07097_ (.Y(_01997_),
    .A(_01958_),
    .B(_01996_));
 sg13g2_and2_1 _07098_ (.A(_01994_),
    .B(_01997_),
    .X(_01998_));
 sg13g2_nor3_1 _07099_ (.A(_01813_),
    .B(_01950_),
    .C(_01951_),
    .Y(_01999_));
 sg13g2_nor4_1 _07100_ (.A(_01749_),
    .B(_01851_),
    .C(_01935_),
    .D(_01999_),
    .Y(_02000_));
 sg13g2_a21oi_1 _07101_ (.A1(_01750_),
    .A2(_01952_),
    .Y(_02001_),
    .B1(_01939_));
 sg13g2_nor4_1 _07102_ (.A(_01749_),
    .B(net24),
    .C(_01935_),
    .D(_01999_),
    .Y(_02002_));
 sg13g2_nor4_1 _07103_ (.A(_01749_),
    .B(net25),
    .C(net24),
    .D(_01999_),
    .Y(_02003_));
 sg13g2_or4_1 _07104_ (.A(_02000_),
    .B(_02001_),
    .C(_02002_),
    .D(_02003_),
    .X(_02004_));
 sg13g2_and2_1 _07105_ (.A(_01938_),
    .B(_01956_),
    .X(_02005_));
 sg13g2_and3_1 _07106_ (.X(_02006_),
    .A(net24),
    .B(_01935_),
    .C(_01956_));
 sg13g2_and3_1 _07107_ (.X(_02007_),
    .A(_01852_),
    .B(_01896_),
    .C(_01956_));
 sg13g2_nor4_1 _07108_ (.A(_01852_),
    .B(_01896_),
    .C(_01935_),
    .D(_01956_),
    .Y(_02008_));
 sg13g2_or4_1 _07109_ (.A(_02005_),
    .B(_02006_),
    .C(_02007_),
    .D(_02008_),
    .X(_02009_));
 sg13g2_or2_1 _07110_ (.X(_02010_),
    .B(_02009_),
    .A(_02004_));
 sg13g2_nor3_1 _07111_ (.A(_01954_),
    .B(_01994_),
    .C(_01997_),
    .Y(_02011_));
 sg13g2_inv_1 _07112_ (.Y(_02012_),
    .A(_01994_));
 sg13g2_nand2_1 _07113_ (.Y(_02013_),
    .A(_01954_),
    .B(_02012_));
 sg13g2_nor4_1 _07114_ (.A(_01997_),
    .B(_02004_),
    .C(_02009_),
    .D(_02013_),
    .Y(_02014_));
 sg13g2_a221oi_1 _07115_ (.B2(_02011_),
    .C1(_02014_),
    .B1(_02010_),
    .A1(_01961_),
    .Y(_02015_),
    .A2(_01998_));
 sg13g2_buf_1 _07116_ (.A(_02015_),
    .X(_02016_));
 sg13g2_inv_1 _07117_ (.Y(_02017_),
    .A(net484));
 sg13g2_buf_1 _07118_ (.A(\median_processor.input_storage [47]),
    .X(_02018_));
 sg13g2_buf_1 _07119_ (.A(net483),
    .X(_02019_));
 sg13g2_inv_1 _07120_ (.Y(_02020_),
    .A(net438));
 sg13g2_buf_1 _07121_ (.A(\median_processor.input_storage [11]),
    .X(_02021_));
 sg13g2_inv_1 _07122_ (.Y(_02022_),
    .A(net475));
 sg13g2_buf_1 _07123_ (.A(\median_processor.input_storage [8]),
    .X(_02023_));
 sg13g2_nand2b_1 _07124_ (.Y(_02024_),
    .B(net434),
    .A_N(net429));
 sg13g2_nand3b_1 _07125_ (.B(net475),
    .C(net434),
    .Y(_02025_),
    .A_N(net429));
 sg13g2_buf_1 _07126_ (.A(\median_processor.input_storage [9]),
    .X(_02026_));
 sg13g2_a22oi_1 _07127_ (.Y(_02027_),
    .B1(_02025_),
    .B2(net428),
    .A2(_02024_),
    .A1(_02022_));
 sg13g2_inv_1 _07128_ (.Y(_02028_),
    .A(\median_processor.input_storage [10]));
 sg13g2_o21ai_1 _07129_ (.B1(_02028_),
    .Y(_02029_),
    .A1(net435),
    .A2(_02027_));
 sg13g2_nand2_1 _07130_ (.Y(_02030_),
    .A(net435),
    .B(_02027_));
 sg13g2_a22oi_1 _07131_ (.Y(_02031_),
    .B1(_02029_),
    .B2(_02030_),
    .A2(_01977_),
    .A1(net430));
 sg13g2_a21oi_1 _07132_ (.A1(_01786_),
    .A2(net433),
    .Y(_02032_),
    .B1(_02031_));
 sg13g2_o21ai_1 _07133_ (.B1(_02032_),
    .Y(_02033_),
    .A1(net431),
    .A2(net390));
 sg13g2_buf_1 _07134_ (.A(net482),
    .X(_02034_));
 sg13g2_inv_1 _07135_ (.Y(_02035_),
    .A(net437));
 sg13g2_inv_2 _07136_ (.Y(_02036_),
    .A(\median_processor.input_storage [14]));
 sg13g2_nor2_1 _07137_ (.A(_02036_),
    .B(net436),
    .Y(_02037_));
 sg13g2_buf_1 _07138_ (.A(net481),
    .X(_02038_));
 sg13g2_a21oi_1 _07139_ (.A1(net439),
    .A2(_02037_),
    .Y(_02039_),
    .B1(_02038_));
 sg13g2_nor2_1 _07140_ (.A(net439),
    .B(_02037_),
    .Y(_02040_));
 sg13g2_nor2_1 _07141_ (.A(_02039_),
    .B(_02040_),
    .Y(_02041_));
 sg13g2_a221oi_1 _07142_ (.B2(net431),
    .C1(_02041_),
    .B1(_02020_),
    .A1(net427),
    .Y(_02042_),
    .A2(net389));
 sg13g2_nor2_1 _07143_ (.A(_02034_),
    .B(net389),
    .Y(_02043_));
 sg13g2_nand2_1 _07144_ (.Y(_02044_),
    .A(net436),
    .B(_02043_));
 sg13g2_o21ai_1 _07145_ (.B1(_02036_),
    .Y(_02045_),
    .A1(net436),
    .A2(_02043_));
 sg13g2_a22oi_1 _07146_ (.Y(_02046_),
    .B1(_02044_),
    .B2(_02045_),
    .A2(net439),
    .A1(_02038_));
 sg13g2_a221oi_1 _07147_ (.B2(_02042_),
    .C1(_02046_),
    .B1(_02033_),
    .A1(_01800_),
    .Y(_02047_),
    .A2(net432));
 sg13g2_buf_1 _07148_ (.A(_02047_),
    .X(_02048_));
 sg13g2_nor2_1 _07149_ (.A(net391),
    .B(net426),
    .Y(_02049_));
 sg13g2_inv_1 _07150_ (.Y(_02050_),
    .A(net478));
 sg13g2_buf_1 _07151_ (.A(\median_processor.input_storage [10]),
    .X(_02051_));
 sg13g2_nor2b_1 _07152_ (.A(net461),
    .B_N(net430),
    .Y(_02052_));
 sg13g2_a21oi_1 _07153_ (.A1(net425),
    .A2(net424),
    .Y(_02053_),
    .B1(_02052_));
 sg13g2_nor2_1 _07154_ (.A(net425),
    .B(net424),
    .Y(_02054_));
 sg13g2_inv_1 _07155_ (.Y(_02055_),
    .A(\median_processor.input_storage [1]));
 sg13g2_nor2b_1 _07156_ (.A(net484),
    .B_N(net429),
    .Y(_02056_));
 sg13g2_o21ai_1 _07157_ (.B1(net428),
    .Y(_02057_),
    .A1(_02055_),
    .A2(_02056_));
 sg13g2_a221oi_1 _07158_ (.B2(_02055_),
    .C1(_02052_),
    .B1(_02056_),
    .A1(net425),
    .Y(_02058_),
    .A2(net424));
 sg13g2_buf_1 _07159_ (.A(\median_processor.input_storage [4]),
    .X(_02059_));
 sg13g2_nand2b_1 _07160_ (.Y(_02060_),
    .B(net423),
    .A_N(net431));
 sg13g2_buf_1 _07161_ (.A(\median_processor.input_storage [5]),
    .X(_02061_));
 sg13g2_nand2b_1 _07162_ (.Y(_02062_),
    .B(net422),
    .A_N(net427));
 sg13g2_nand2b_1 _07163_ (.Y(_02063_),
    .B(net461),
    .A_N(net430));
 sg13g2_nand3_1 _07164_ (.B(_02062_),
    .C(_02063_),
    .A(_02060_),
    .Y(_02064_));
 sg13g2_a221oi_1 _07165_ (.B2(_02058_),
    .C1(_02064_),
    .B1(_02057_),
    .A1(_02053_),
    .Y(_02065_),
    .A2(_02054_));
 sg13g2_nor2b_1 _07166_ (.A(net423),
    .B_N(net431),
    .Y(_02066_));
 sg13g2_nand2_1 _07167_ (.Y(_02067_),
    .A(net427),
    .B(_02066_));
 sg13g2_o21ai_1 _07168_ (.B1(_01762_),
    .Y(_02068_),
    .A1(net427),
    .A2(_02066_));
 sg13g2_nand2_1 _07169_ (.Y(_02069_),
    .A(_02067_),
    .B(_02068_));
 sg13g2_nand2_1 _07170_ (.Y(_02070_),
    .A(net440),
    .B(_02036_));
 sg13g2_o21ai_1 _07171_ (.B1(_02070_),
    .Y(_02071_),
    .A1(_02065_),
    .A2(_02069_));
 sg13g2_buf_1 _07172_ (.A(\median_processor.input_storage [14]),
    .X(_02072_));
 sg13g2_nand2_1 _07173_ (.Y(_02073_),
    .A(net462),
    .B(net421));
 sg13g2_and2_1 _07174_ (.A(_02071_),
    .B(_02073_),
    .X(_02074_));
 sg13g2_nand2_1 _07175_ (.Y(_02075_),
    .A(net391),
    .B(net426));
 sg13g2_and2_1 _07176_ (.A(net28),
    .B(_02075_),
    .X(_02076_));
 sg13g2_o21ai_1 _07177_ (.B1(_02076_),
    .Y(_02077_),
    .A1(_02049_),
    .A2(_02074_));
 sg13g2_nor2_1 _07178_ (.A(net462),
    .B(net421),
    .Y(_02078_));
 sg13g2_or2_1 _07179_ (.X(_02079_),
    .B(_02066_),
    .A(net427));
 sg13g2_nand2_1 _07180_ (.Y(_02080_),
    .A(net422),
    .B(_02067_));
 sg13g2_a221oi_1 _07181_ (.B2(_02080_),
    .C1(_02065_),
    .B1(_02079_),
    .A1(net462),
    .Y(_02081_),
    .A2(net421));
 sg13g2_nand2_1 _07182_ (.Y(_02082_),
    .A(net426),
    .B(net393));
 sg13g2_nor4_1 _07183_ (.A(net28),
    .B(_02078_),
    .C(_02081_),
    .D(_02082_),
    .Y(_02083_));
 sg13g2_nor3_1 _07184_ (.A(_01714_),
    .B(net28),
    .C(_02075_),
    .Y(_02084_));
 sg13g2_nor2_1 _07185_ (.A(_01800_),
    .B(net393),
    .Y(_02085_));
 sg13g2_and4_1 _07186_ (.A(net472),
    .B(_02085_),
    .C(_02071_),
    .D(_02073_),
    .X(_02086_));
 sg13g2_nand2_1 _07187_ (.Y(_02087_),
    .A(net391),
    .B(_01800_));
 sg13g2_nor4_1 _07188_ (.A(net28),
    .B(_02087_),
    .C(_02078_),
    .D(_02081_),
    .Y(_02088_));
 sg13g2_nor4_1 _07189_ (.A(_02083_),
    .B(_02084_),
    .C(_02086_),
    .D(_02088_),
    .Y(_02089_));
 sg13g2_nand2_1 _07190_ (.Y(_02090_),
    .A(_02077_),
    .B(_02089_));
 sg13g2_nand2_1 _07191_ (.Y(_02091_),
    .A(_02071_),
    .B(_02073_));
 sg13g2_a21oi_1 _07192_ (.A1(net426),
    .A2(_02091_),
    .Y(_02092_),
    .B1(net391));
 sg13g2_nand2_1 _07193_ (.Y(_02093_),
    .A(net393),
    .B(_01945_));
 sg13g2_a22oi_1 _07194_ (.Y(_02094_),
    .B1(_02091_),
    .B2(net28),
    .A2(_02093_),
    .A1(net426));
 sg13g2_nor3_1 _07195_ (.A(net14),
    .B(_02092_),
    .C(_02094_),
    .Y(_02095_));
 sg13g2_a21o_1 _07196_ (.A2(_02090_),
    .A1(net14),
    .B1(_02095_),
    .X(_02096_));
 sg13g2_nor2_1 _07197_ (.A(_01869_),
    .B(net482),
    .Y(_02097_));
 sg13g2_nand2b_1 _07198_ (.Y(_02098_),
    .B(\median_processor.input_storage [51]),
    .A_N(\median_processor.input_storage [11]));
 sg13g2_inv_2 _07199_ (.Y(_02099_),
    .A(net450));
 sg13g2_a221oi_1 _07200_ (.B2(_02098_),
    .C1(_02099_),
    .B1(net483),
    .A1(_01869_),
    .Y(_02100_),
    .A2(net482));
 sg13g2_nor2b_1 _07201_ (.A(net449),
    .B_N(net482),
    .Y(_02101_));
 sg13g2_nor3_1 _07202_ (.A(net483),
    .B(_02101_),
    .C(_02098_),
    .Y(_02102_));
 sg13g2_nor3_1 _07203_ (.A(_02097_),
    .B(_02100_),
    .C(_02102_),
    .Y(_02103_));
 sg13g2_buf_1 _07204_ (.A(\median_processor.input_storage [50]),
    .X(_02104_));
 sg13g2_nand2b_1 _07205_ (.Y(_02105_),
    .B(\median_processor.input_storage [8]),
    .A_N(net448));
 sg13g2_inv_1 _07206_ (.Y(_02106_),
    .A(\median_processor.input_storage [9]));
 sg13g2_a221oi_1 _07207_ (.B2(net474),
    .C1(_02106_),
    .B1(_02105_),
    .A1(net420),
    .Y(_02107_),
    .A2(_02028_));
 sg13g2_xor2_1 _07208_ (.B(\median_processor.input_storage [12]),
    .A(\median_processor.input_storage [52]),
    .X(_02108_));
 sg13g2_nor2b_1 _07209_ (.A(\median_processor.input_storage [51]),
    .B_N(\median_processor.input_storage [11]),
    .Y(_02109_));
 sg13g2_nor2b_1 _07210_ (.A(\median_processor.input_storage [50]),
    .B_N(\median_processor.input_storage [10]),
    .Y(_02110_));
 sg13g2_nor4_2 _07211_ (.A(_02101_),
    .B(_02108_),
    .C(_02109_),
    .Y(_02111_),
    .D(_02110_));
 sg13g2_nand2b_1 _07212_ (.Y(_02112_),
    .B(\median_processor.input_storage [50]),
    .A_N(\median_processor.input_storage [10]));
 sg13g2_nand4_1 _07213_ (.B(_01876_),
    .C(\median_processor.input_storage [8]),
    .A(_01882_),
    .Y(_02113_),
    .D(_02112_));
 sg13g2_nand3b_1 _07214_ (.B(_02111_),
    .C(_02113_),
    .Y(_02114_),
    .A_N(_02107_));
 sg13g2_xnor2_1 _07215_ (.Y(_02115_),
    .A(net474),
    .B(\median_processor.input_storage [9]));
 sg13g2_nand2b_1 _07216_ (.Y(_02116_),
    .B(net448),
    .A_N(\median_processor.input_storage [8]));
 sg13g2_xnor2_1 _07217_ (.Y(_02117_),
    .A(\median_processor.input_storage [54]),
    .B(\median_processor.input_storage [14]));
 sg13g2_nand4_1 _07218_ (.B(_02115_),
    .C(_02116_),
    .A(_02105_),
    .Y(_02118_),
    .D(_02117_));
 sg13g2_nand2_1 _07219_ (.Y(_02119_),
    .A(_02098_),
    .B(_02112_));
 sg13g2_nor3_1 _07220_ (.A(_02097_),
    .B(_02118_),
    .C(_02119_),
    .Y(_02120_));
 sg13g2_nand2_1 _07221_ (.Y(_02121_),
    .A(net446),
    .B(net481));
 sg13g2_nand2_1 _07222_ (.Y(_02122_),
    .A(_02036_),
    .B(_02121_));
 sg13g2_a221oi_1 _07223_ (.B2(_02111_),
    .C1(_02122_),
    .B1(_02120_),
    .A1(_02103_),
    .Y(_02123_),
    .A2(_02114_));
 sg13g2_nand2_1 _07224_ (.Y(_02124_),
    .A(net447),
    .B(_02121_));
 sg13g2_a221oi_1 _07225_ (.B2(_02111_),
    .C1(_02124_),
    .B1(_02120_),
    .A1(_02103_),
    .Y(_02125_),
    .A2(_02114_));
 sg13g2_nand3_1 _07226_ (.B(_02036_),
    .C(_02121_),
    .A(net447),
    .Y(_02126_));
 sg13g2_o21ai_1 _07227_ (.B1(_02126_),
    .Y(_02127_),
    .A1(net446),
    .A2(net481));
 sg13g2_or3_1 _07228_ (.A(_02123_),
    .B(_02125_),
    .C(_02127_),
    .X(_02128_));
 sg13g2_buf_2 _07229_ (.A(_02128_),
    .X(_02129_));
 sg13g2_nand2_1 _07230_ (.Y(_02130_),
    .A(net469),
    .B(_01800_));
 sg13g2_inv_2 _07231_ (.Y(_02131_),
    .A(net469));
 sg13g2_nand2_1 _07232_ (.Y(_02132_),
    .A(_02131_),
    .B(\median_processor.input_storage [15]));
 sg13g2_buf_1 _07233_ (.A(\median_processor.input_storage [28]),
    .X(_02133_));
 sg13g2_nor2_1 _07234_ (.A(_02034_),
    .B(net431),
    .Y(_02134_));
 sg13g2_nand2_1 _07235_ (.Y(_02135_),
    .A(net419),
    .B(_02134_));
 sg13g2_nor2b_1 _07236_ (.A(net431),
    .B_N(net419),
    .Y(_02136_));
 sg13g2_buf_1 _07237_ (.A(\median_processor.input_storage [29]),
    .X(_02137_));
 sg13g2_o21ai_1 _07238_ (.B1(net418),
    .Y(_02138_),
    .A1(_01781_),
    .A2(_02136_));
 sg13g2_a21oi_1 _07239_ (.A1(_02135_),
    .A2(_02138_),
    .Y(_02139_),
    .B1(net421));
 sg13g2_nand2_1 _07240_ (.Y(_02140_),
    .A(_02132_),
    .B(_02139_));
 sg13g2_buf_1 _07241_ (.A(\median_processor.input_storage [30]),
    .X(_02141_));
 sg13g2_nand3_1 _07242_ (.B(_02135_),
    .C(_02138_),
    .A(net421),
    .Y(_02142_));
 sg13g2_nand3_1 _07243_ (.B(_02132_),
    .C(_02142_),
    .A(net417),
    .Y(_02143_));
 sg13g2_xnor2_1 _07244_ (.Y(_02144_),
    .A(net419),
    .B(_02019_));
 sg13g2_xor2_1 _07245_ (.B(\median_processor.input_storage [13]),
    .A(\median_processor.input_storage [29]),
    .X(_02145_));
 sg13g2_xor2_1 _07246_ (.B(net421),
    .A(net417),
    .X(_02146_));
 sg13g2_nor2_1 _07247_ (.A(_02145_),
    .B(_02146_),
    .Y(_02147_));
 sg13g2_nand4_1 _07248_ (.B(_02132_),
    .C(_02130_),
    .A(_02144_),
    .Y(_02148_),
    .D(_02147_));
 sg13g2_xor2_1 _07249_ (.B(net428),
    .A(net479),
    .X(_02149_));
 sg13g2_inv_1 _07250_ (.Y(_02150_),
    .A(\median_processor.input_storage [26]));
 sg13g2_nor2_1 _07251_ (.A(net416),
    .B(net424),
    .Y(_02151_));
 sg13g2_nor2b_1 _07252_ (.A(\median_processor.input_storage [26]),
    .B_N(net424),
    .Y(_02152_));
 sg13g2_nor2b_1 _07253_ (.A(net467),
    .B_N(net429),
    .Y(_02153_));
 sg13g2_nand2b_1 _07254_ (.Y(_02154_),
    .B(net467),
    .A_N(net429));
 sg13g2_xnor2_1 _07255_ (.Y(_02155_),
    .A(net466),
    .B(\median_processor.input_storage [11]));
 sg13g2_nand3b_1 _07256_ (.B(_02154_),
    .C(_02155_),
    .Y(_02156_),
    .A_N(_02153_));
 sg13g2_nor4_1 _07257_ (.A(_02149_),
    .B(_02151_),
    .C(_02152_),
    .D(_02156_),
    .Y(_02157_));
 sg13g2_o21ai_1 _07258_ (.B1(_01727_),
    .Y(_02158_),
    .A1(net428),
    .A2(_02153_));
 sg13g2_inv_1 _07259_ (.Y(_02159_),
    .A(\median_processor.input_storage [24]));
 sg13g2_nand3_1 _07260_ (.B(net428),
    .C(net429),
    .A(_02159_),
    .Y(_02160_));
 sg13g2_a221oi_1 _07261_ (.B2(_02160_),
    .C1(_02151_),
    .B1(_02158_),
    .A1(net466),
    .Y(_02161_),
    .A2(_01786_));
 sg13g2_o21ai_1 _07262_ (.B1(_02152_),
    .Y(_02162_),
    .A1(net465),
    .A2(net430));
 sg13g2_o21ai_1 _07263_ (.B1(_02162_),
    .Y(_02163_),
    .A1(net466),
    .A2(_01786_));
 sg13g2_or4_1 _07264_ (.A(_02148_),
    .B(_02157_),
    .C(_02161_),
    .D(_02163_),
    .X(_02164_));
 sg13g2_nand4_1 _07265_ (.B(_02140_),
    .C(_02143_),
    .A(_02130_),
    .Y(_02165_),
    .D(_02164_));
 sg13g2_buf_1 _07266_ (.A(_02165_),
    .X(_02166_));
 sg13g2_and2_1 _07267_ (.A(_02129_),
    .B(net23),
    .X(_02167_));
 sg13g2_buf_1 _07268_ (.A(\median_processor.input_storage [36]),
    .X(_02168_));
 sg13g2_nand2_1 _07269_ (.Y(_02169_),
    .A(net415),
    .B(_02134_));
 sg13g2_nor2b_1 _07270_ (.A(_02019_),
    .B_N(\median_processor.input_storage [36]),
    .Y(_02170_));
 sg13g2_o21ai_1 _07271_ (.B1(net476),
    .Y(_02171_),
    .A1(_01781_),
    .A2(_02170_));
 sg13g2_a21oi_1 _07272_ (.A1(_02169_),
    .A2(_02171_),
    .Y(_02172_),
    .B1(_02072_));
 sg13g2_a21oi_1 _07273_ (.A1(net415),
    .A2(_02134_),
    .Y(_02173_),
    .B1(_02036_));
 sg13g2_a21oi_1 _07274_ (.A1(_02171_),
    .A2(_02173_),
    .Y(_02174_),
    .B1(net392));
 sg13g2_nand2_1 _07275_ (.Y(_02175_),
    .A(net222),
    .B(net481));
 sg13g2_o21ai_1 _07276_ (.B1(_02175_),
    .Y(_02176_),
    .A1(_02172_),
    .A2(_02174_));
 sg13g2_buf_1 _07277_ (.A(\median_processor.input_storage [33]),
    .X(_02177_));
 sg13g2_nand2b_1 _07278_ (.Y(_02178_),
    .B(net429),
    .A_N(net477));
 sg13g2_a21oi_1 _07279_ (.A1(net414),
    .A2(_02178_),
    .Y(_02179_),
    .B1(_02106_));
 sg13g2_nor2_1 _07280_ (.A(net414),
    .B(_02178_),
    .Y(_02180_));
 sg13g2_nor2b_1 _07281_ (.A(net424),
    .B_N(net441),
    .Y(_02181_));
 sg13g2_a21oi_1 _07282_ (.A1(net442),
    .A2(_01786_),
    .Y(_02182_),
    .B1(_02181_));
 sg13g2_o21ai_1 _07283_ (.B1(_02182_),
    .Y(_02183_),
    .A1(_02179_),
    .A2(_02180_));
 sg13g2_xor2_1 _07284_ (.B(net481),
    .A(net444),
    .X(_02184_));
 sg13g2_xor2_1 _07285_ (.B(net483),
    .A(\median_processor.input_storage [36]),
    .X(_02185_));
 sg13g2_xor2_1 _07286_ (.B(net482),
    .A(net476),
    .X(_02186_));
 sg13g2_xor2_1 _07287_ (.B(_02072_),
    .A(net445),
    .X(_02187_));
 sg13g2_nor4_1 _07288_ (.A(_02184_),
    .B(_02185_),
    .C(_02186_),
    .D(_02187_),
    .Y(_02188_));
 sg13g2_inv_2 _07289_ (.Y(_02189_),
    .A(\median_processor.input_storage [35]));
 sg13g2_nand2_1 _07290_ (.Y(_02190_),
    .A(_02189_),
    .B(net430));
 sg13g2_nor2b_1 _07291_ (.A(net441),
    .B_N(_02051_),
    .Y(_02191_));
 sg13g2_o21ai_1 _07292_ (.B1(_02191_),
    .Y(_02192_),
    .A1(_02189_),
    .A2(_02021_));
 sg13g2_and3_1 _07293_ (.X(_02193_),
    .A(_02188_),
    .B(_02190_),
    .C(_02192_));
 sg13g2_a22oi_1 _07294_ (.Y(_02194_),
    .B1(_02183_),
    .B2(_02193_),
    .A2(_01800_),
    .A1(net444));
 sg13g2_xor2_1 _07295_ (.B(net428),
    .A(net414),
    .X(_02195_));
 sg13g2_nor3_1 _07296_ (.A(_02195_),
    .B(_02191_),
    .C(_02181_),
    .Y(_02196_));
 sg13g2_xnor2_1 _07297_ (.Y(_02197_),
    .A(net477),
    .B(_02023_));
 sg13g2_xnor2_1 _07298_ (.Y(_02198_),
    .A(net442),
    .B(_02021_));
 sg13g2_nand4_1 _07299_ (.B(_02196_),
    .C(_02197_),
    .A(_02188_),
    .Y(_02199_),
    .D(_02198_));
 sg13g2_inv_1 _07300_ (.Y(_02200_),
    .A(_02199_));
 sg13g2_a21oi_1 _07301_ (.A1(_02176_),
    .A2(_02194_),
    .Y(_02201_),
    .B1(_02200_));
 sg13g2_nor2_1 _07302_ (.A(_01846_),
    .B(net481),
    .Y(_02202_));
 sg13g2_nand2b_1 _07303_ (.Y(_02203_),
    .B(net457),
    .A_N(_02023_));
 sg13g2_o21ai_1 _07304_ (.B1(_02203_),
    .Y(_02204_),
    .A1(net458),
    .A2(_02026_));
 sg13g2_a22oi_1 _07305_ (.Y(_02205_),
    .B1(_02026_),
    .B2(net458),
    .A2(_02051_),
    .A1(_01814_));
 sg13g2_nand2b_1 _07306_ (.Y(_02206_),
    .B(\median_processor.input_storage [60]),
    .A_N(net483));
 sg13g2_nand2b_1 _07307_ (.Y(_02207_),
    .B(\median_processor.input_storage [61]),
    .A_N(net482));
 sg13g2_nand2b_1 _07308_ (.Y(_02208_),
    .B(net454),
    .A_N(\median_processor.input_storage [10]));
 sg13g2_nand4_1 _07309_ (.B(_02206_),
    .C(_02207_),
    .A(net430),
    .Y(_02209_),
    .D(_02208_));
 sg13g2_inv_1 _07310_ (.Y(_02210_),
    .A(\median_processor.input_storage [59]));
 sg13g2_nand4_1 _07311_ (.B(_02206_),
    .C(_02207_),
    .A(_02210_),
    .Y(_02211_),
    .D(_02208_));
 sg13g2_a22oi_1 _07312_ (.Y(_02212_),
    .B1(_02209_),
    .B2(_02211_),
    .A2(_02205_),
    .A1(_02204_));
 sg13g2_nor2b_1 _07313_ (.A(\median_processor.input_storage [60]),
    .B_N(net483),
    .Y(_02213_));
 sg13g2_nand2_1 _07314_ (.Y(_02214_),
    .A(net427),
    .B(_02213_));
 sg13g2_o21ai_1 _07315_ (.B1(net395),
    .Y(_02215_),
    .A1(net482),
    .A2(_02213_));
 sg13g2_nand4_1 _07316_ (.B(\median_processor.input_storage [11]),
    .C(_02206_),
    .A(_02210_),
    .Y(_02216_),
    .D(_02207_));
 sg13g2_nand3_1 _07317_ (.B(_02215_),
    .C(_02216_),
    .A(_02214_),
    .Y(_02217_));
 sg13g2_nand2_1 _07318_ (.Y(_02218_),
    .A(_01846_),
    .B(net481));
 sg13g2_nand2_1 _07319_ (.Y(_02219_),
    .A(_02036_),
    .B(_02218_));
 sg13g2_nor3_1 _07320_ (.A(_02212_),
    .B(_02217_),
    .C(_02219_),
    .Y(_02220_));
 sg13g2_nand2_1 _07321_ (.Y(_02221_),
    .A(net452),
    .B(_02218_));
 sg13g2_nor3_1 _07322_ (.A(_02212_),
    .B(_02217_),
    .C(_02221_),
    .Y(_02222_));
 sg13g2_buf_1 _07323_ (.A(net452),
    .X(_02223_));
 sg13g2_and3_1 _07324_ (.X(_02224_),
    .A(net388),
    .B(_02036_),
    .C(_02218_));
 sg13g2_or4_1 _07325_ (.A(_02202_),
    .B(_02220_),
    .C(_02222_),
    .D(_02224_),
    .X(_02225_));
 sg13g2_buf_1 _07326_ (.A(_02225_),
    .X(_02226_));
 sg13g2_nor2_1 _07327_ (.A(net26),
    .B(net22),
    .Y(_02227_));
 sg13g2_nor2_1 _07328_ (.A(_02129_),
    .B(net23),
    .Y(_02228_));
 sg13g2_and2_1 _07329_ (.A(net26),
    .B(net22),
    .X(_02229_));
 sg13g2_a22oi_1 _07330_ (.Y(_02230_),
    .B1(_02228_),
    .B2(_02229_),
    .A2(_02227_),
    .A1(_02167_));
 sg13g2_xnor2_1 _07331_ (.Y(_02231_),
    .A(_02129_),
    .B(_02165_));
 sg13g2_or3_1 _07332_ (.A(_02229_),
    .B(_02227_),
    .C(_02231_),
    .X(_02232_));
 sg13g2_nand2_1 _07333_ (.Y(_02233_),
    .A(_02230_),
    .B(_02232_));
 sg13g2_nor2_1 _07334_ (.A(net23),
    .B(net22),
    .Y(_02234_));
 sg13g2_a21oi_1 _07335_ (.A1(_02077_),
    .A2(_02089_),
    .Y(_02235_),
    .B1(net26));
 sg13g2_o21ai_1 _07336_ (.B1(_02235_),
    .Y(_02236_),
    .A1(_02228_),
    .A2(_02234_));
 sg13g2_nor2_1 _07337_ (.A(_02129_),
    .B(net22),
    .Y(_02237_));
 sg13g2_nand2_1 _07338_ (.Y(_02238_),
    .A(_02235_),
    .B(_02237_));
 sg13g2_inv_2 _07339_ (.Y(_02239_),
    .A(net26));
 sg13g2_nor3_1 _07340_ (.A(_02129_),
    .B(net23),
    .C(net22),
    .Y(_02240_));
 sg13g2_o21ai_1 _07341_ (.B1(_02240_),
    .Y(_02241_),
    .A1(_02239_),
    .A2(_02090_));
 sg13g2_nand3_1 _07342_ (.B(_02238_),
    .C(_02241_),
    .A(_02236_),
    .Y(_02242_));
 sg13g2_o21ai_1 _07343_ (.B1(_02075_),
    .Y(_02243_),
    .A1(_02049_),
    .A2(_02074_));
 sg13g2_nor3_1 _07344_ (.A(net28),
    .B(_02085_),
    .C(_02243_),
    .Y(_02244_));
 sg13g2_xor2_1 _07345_ (.B(net22),
    .A(net26),
    .X(_02245_));
 sg13g2_xnor2_1 _07346_ (.Y(_02246_),
    .A(_02245_),
    .B(_02231_));
 sg13g2_mux2_1 _07347_ (.A0(_02244_),
    .A1(_02090_),
    .S(_02246_),
    .X(_02247_));
 sg13g2_nor2b_1 _07348_ (.A(net14),
    .B_N(_02247_),
    .Y(_02248_));
 sg13g2_nand2_1 _07349_ (.Y(_02249_),
    .A(net26),
    .B(net23));
 sg13g2_o21ai_1 _07350_ (.B1(net22),
    .Y(_02250_),
    .A1(_02201_),
    .A2(_02165_));
 sg13g2_nor3_1 _07351_ (.A(_02123_),
    .B(_02125_),
    .C(_02127_),
    .Y(_02251_));
 sg13g2_a21o_1 _07352_ (.A2(_02250_),
    .A1(_02249_),
    .B1(_02251_),
    .X(_02252_));
 sg13g2_nand3_1 _07353_ (.B(net23),
    .C(net22),
    .A(_02201_),
    .Y(_02253_));
 sg13g2_nand4_1 _07354_ (.B(net14),
    .C(_02244_),
    .A(_02252_),
    .Y(_02254_),
    .D(_02253_));
 sg13g2_a21o_1 _07355_ (.A2(net23),
    .A1(net26),
    .B1(_02129_),
    .X(_02255_));
 sg13g2_nor2_1 _07356_ (.A(net26),
    .B(net23),
    .Y(_02256_));
 sg13g2_a21oi_1 _07357_ (.A1(net28),
    .A2(_02091_),
    .Y(_02257_),
    .B1(net426));
 sg13g2_nor3_1 _07358_ (.A(_02256_),
    .B(_02092_),
    .C(_02257_),
    .Y(_02258_));
 sg13g2_nand4_1 _07359_ (.B(net14),
    .C(_02255_),
    .A(_02093_),
    .Y(_02259_),
    .D(_02258_));
 sg13g2_nand2_1 _07360_ (.Y(_02260_),
    .A(_02245_),
    .B(_02231_));
 sg13g2_nor2_1 _07361_ (.A(_02251_),
    .B(_02229_),
    .Y(_02261_));
 sg13g2_or2_1 _07362_ (.X(_02262_),
    .B(_02231_),
    .A(_02245_));
 sg13g2_a21o_1 _07363_ (.A2(_02261_),
    .A1(_02090_),
    .B1(_02262_),
    .X(_02263_));
 sg13g2_a22oi_1 _07364_ (.Y(_02264_),
    .B1(_02260_),
    .B2(_02263_),
    .A2(_02259_),
    .A1(_02254_));
 sg13g2_a221oi_1 _07365_ (.B2(_02248_),
    .C1(_02264_),
    .B1(_02242_),
    .A1(_02096_),
    .Y(_02265_),
    .A2(_02233_));
 sg13g2_mux2_1 _07366_ (.A0(_01793_),
    .A1(_02017_),
    .S(_02265_),
    .X(_02266_));
 sg13g2_nand2_1 _07367_ (.Y(_02267_),
    .A(net7),
    .B(_02266_));
 sg13g2_or2_1 _07368_ (.X(_02268_),
    .B(net7),
    .A(net463));
 sg13g2_a22oi_1 _07369_ (.Y(_02269_),
    .B1(_01968_),
    .B2(_01762_),
    .A2(net432),
    .A1(_01808_));
 sg13g2_o21ai_1 _07370_ (.B1(_02269_),
    .Y(_02270_),
    .A1(net440),
    .A2(_01965_));
 sg13g2_inv_1 _07371_ (.Y(_02271_),
    .A(_02270_));
 sg13g2_a21o_1 _07372_ (.A2(net434),
    .A1(_02017_),
    .B1(net475),
    .X(_02272_));
 sg13g2_o21ai_1 _07373_ (.B1(\median_processor.input_storage [1]),
    .Y(_02273_),
    .A1(net484),
    .A2(_01975_));
 sg13g2_nor2_1 _07374_ (.A(net461),
    .B(_01977_),
    .Y(_02274_));
 sg13g2_a221oi_1 _07375_ (.B2(_02273_),
    .C1(_02274_),
    .B1(_02272_),
    .A1(net425),
    .Y(_02275_),
    .A2(net435));
 sg13g2_nand2_1 _07376_ (.Y(_02276_),
    .A(net478),
    .B(_01979_));
 sg13g2_nand2_1 _07377_ (.Y(_02277_),
    .A(net461),
    .B(_01977_));
 sg13g2_o21ai_1 _07378_ (.B1(_02277_),
    .Y(_02278_),
    .A1(_02274_),
    .A2(_02276_));
 sg13g2_nor3_1 _07379_ (.A(net390),
    .B(_02275_),
    .C(_02278_),
    .Y(_02279_));
 sg13g2_o21ai_1 _07380_ (.B1(net390),
    .Y(_02280_),
    .A1(_02275_),
    .A2(_02278_));
 sg13g2_o21ai_1 _07381_ (.B1(_02280_),
    .Y(_02281_),
    .A1(_01764_),
    .A2(_02279_));
 sg13g2_nand2_1 _07382_ (.Y(_02282_),
    .A(net422),
    .B(_02035_));
 sg13g2_a21oi_1 _07383_ (.A1(net436),
    .A2(_02282_),
    .Y(_02283_),
    .B1(_01751_));
 sg13g2_nor2_1 _07384_ (.A(_01972_),
    .B(_02282_),
    .Y(_02284_));
 sg13g2_nand2_1 _07385_ (.Y(_02285_),
    .A(_01808_),
    .B(net432));
 sg13g2_o21ai_1 _07386_ (.B1(_02285_),
    .Y(_02286_),
    .A1(_02283_),
    .A2(_02284_));
 sg13g2_o21ai_1 _07387_ (.B1(_02286_),
    .Y(_02287_),
    .A1(net391),
    .A2(net432));
 sg13g2_a21o_1 _07388_ (.A2(_02281_),
    .A1(_02271_),
    .B1(_02287_),
    .X(_02288_));
 sg13g2_buf_1 _07389_ (.A(_02288_),
    .X(_02289_));
 sg13g2_nor2_1 _07390_ (.A(net388),
    .B(_01965_),
    .Y(_02290_));
 sg13g2_nor2b_1 _07391_ (.A(net454),
    .B_N(net435),
    .Y(_02291_));
 sg13g2_nor2b_1 _07392_ (.A(net457),
    .B_N(net434),
    .Y(_02292_));
 sg13g2_nor3_1 _07393_ (.A(net458),
    .B(_02291_),
    .C(_02292_),
    .Y(_02293_));
 sg13g2_a221oi_1 _07394_ (.B2(net458),
    .C1(net475),
    .B1(_02292_),
    .A1(_01814_),
    .Y(_02294_),
    .A2(net435));
 sg13g2_nand2b_1 _07395_ (.Y(_02295_),
    .B(net454),
    .A_N(net435));
 sg13g2_nand2b_1 _07396_ (.Y(_02296_),
    .B(net453),
    .A_N(net433));
 sg13g2_nand2b_1 _07397_ (.Y(_02297_),
    .B(net455),
    .A_N(net437));
 sg13g2_nand2b_1 _07398_ (.Y(_02298_),
    .B(\median_processor.input_storage [60]),
    .A_N(net438));
 sg13g2_nand4_1 _07399_ (.B(_02296_),
    .C(_02297_),
    .A(_02295_),
    .Y(_02299_),
    .D(_02298_));
 sg13g2_nor4_1 _07400_ (.A(net388),
    .B(_02293_),
    .C(_02294_),
    .D(_02299_),
    .Y(_02300_));
 sg13g2_nor3_1 _07401_ (.A(net432),
    .B(_02290_),
    .C(_02300_),
    .Y(_02301_));
 sg13g2_nor3_1 _07402_ (.A(net394),
    .B(_02290_),
    .C(_02300_),
    .Y(_02302_));
 sg13g2_nor2b_1 _07403_ (.A(net453),
    .B_N(net433),
    .Y(_02303_));
 sg13g2_a21oi_1 _07404_ (.A1(net438),
    .A2(_02303_),
    .Y(_02304_),
    .B1(net395));
 sg13g2_a21oi_1 _07405_ (.A1(net438),
    .A2(_02303_),
    .Y(_02305_),
    .B1(net437));
 sg13g2_buf_1 _07406_ (.A(_01830_),
    .X(_02306_));
 sg13g2_o21ai_1 _07407_ (.B1(net387),
    .Y(_02307_),
    .A1(net438),
    .A2(_02303_));
 sg13g2_o21ai_1 _07408_ (.B1(_02307_),
    .Y(_02308_),
    .A1(_02304_),
    .A2(_02305_));
 sg13g2_a22oi_1 _07409_ (.Y(_02309_),
    .B1(net389),
    .B2(net455),
    .A2(_01965_),
    .A1(net388));
 sg13g2_xnor2_1 _07410_ (.Y(_02310_),
    .A(net457),
    .B(net434));
 sg13g2_xnor2_1 _07411_ (.Y(_02311_),
    .A(\median_processor.input_storage [57]),
    .B(net475));
 sg13g2_xnor2_1 _07412_ (.Y(_02312_),
    .A(net452),
    .B(\median_processor.input_storage [46]));
 sg13g2_a22oi_1 _07413_ (.Y(_02313_),
    .B1(net438),
    .B2(net387),
    .A2(net437),
    .A1(net395));
 sg13g2_and4_1 _07414_ (.A(_02310_),
    .B(_02311_),
    .C(_02312_),
    .D(_02313_),
    .X(_02314_));
 sg13g2_nor2_1 _07415_ (.A(net473),
    .B(net439),
    .Y(_02315_));
 sg13g2_nor4_1 _07416_ (.A(_02291_),
    .B(_02299_),
    .C(_02303_),
    .D(_02315_),
    .Y(_02316_));
 sg13g2_nor4_1 _07417_ (.A(_01965_),
    .B(_02293_),
    .C(_02294_),
    .D(_02299_),
    .Y(_02317_));
 sg13g2_a221oi_1 _07418_ (.B2(_02316_),
    .C1(_02317_),
    .B1(_02314_),
    .A1(_02308_),
    .Y(_02318_),
    .A2(_02309_));
 sg13g2_o21ai_1 _07419_ (.B1(_02318_),
    .Y(_02319_),
    .A1(_02301_),
    .A2(_02302_));
 sg13g2_nand2_1 _07420_ (.Y(_02320_),
    .A(net473),
    .B(net439));
 sg13g2_and2_1 _07421_ (.A(_02319_),
    .B(_02320_),
    .X(_02321_));
 sg13g2_xnor2_1 _07422_ (.Y(_02322_),
    .A(net17),
    .B(_02321_));
 sg13g2_a22oi_1 _07423_ (.Y(_02323_),
    .B1(_01972_),
    .B2(net392),
    .A2(net432),
    .A1(net222));
 sg13g2_nand2_1 _07424_ (.Y(_02324_),
    .A(_02035_),
    .B(_02323_));
 sg13g2_nand2_1 _07425_ (.Y(_02325_),
    .A(net476),
    .B(_02323_));
 sg13g2_inv_2 _07426_ (.Y(_02326_),
    .A(\median_processor.input_storage [34]));
 sg13g2_a21o_1 _07427_ (.A2(net434),
    .A1(_01907_),
    .B1(net475),
    .X(_02327_));
 sg13g2_o21ai_1 _07428_ (.B1(net414),
    .Y(_02328_),
    .A1(\median_processor.input_storage [32]),
    .A2(_01975_));
 sg13g2_a22oi_1 _07429_ (.Y(_02329_),
    .B1(_02327_),
    .B2(_02328_),
    .A2(_01978_),
    .A1(_02326_));
 sg13g2_a21o_1 _07430_ (.A2(_01979_),
    .A1(net441),
    .B1(_02329_),
    .X(_02330_));
 sg13g2_nor2_1 _07431_ (.A(net415),
    .B(net390),
    .Y(_02331_));
 sg13g2_a21oi_1 _07432_ (.A1(_02189_),
    .A2(net433),
    .Y(_02332_),
    .B1(_02331_));
 sg13g2_nor3_1 _07433_ (.A(_02189_),
    .B(net433),
    .C(_02331_),
    .Y(_02333_));
 sg13g2_a221oi_1 _07434_ (.B2(_02332_),
    .C1(_02333_),
    .B1(_02330_),
    .A1(net415),
    .Y(_02334_),
    .A2(net390));
 sg13g2_a21o_1 _07435_ (.A2(_02325_),
    .A1(_02324_),
    .B1(_02334_),
    .X(_02335_));
 sg13g2_nand2_1 _07436_ (.Y(_02336_),
    .A(net445),
    .B(_01965_));
 sg13g2_nand2_1 _07437_ (.Y(_02337_),
    .A(net432),
    .B(_02336_));
 sg13g2_o21ai_1 _07438_ (.B1(net222),
    .Y(_02338_),
    .A1(_02018_),
    .A2(_02336_));
 sg13g2_nor2_1 _07439_ (.A(net443),
    .B(_01968_),
    .Y(_02339_));
 sg13g2_a22oi_1 _07440_ (.Y(_02340_),
    .B1(_02323_),
    .B2(_02339_),
    .A2(_02338_),
    .A1(_02337_));
 sg13g2_nand2_2 _07441_ (.Y(_02341_),
    .A(_02335_),
    .B(_02340_));
 sg13g2_nand2_1 _07442_ (.Y(_02342_),
    .A(_02322_),
    .B(_02341_));
 sg13g2_nand2_2 _07443_ (.Y(_02343_),
    .A(_02319_),
    .B(_02320_));
 sg13g2_and2_1 _07444_ (.A(_02335_),
    .B(_02340_),
    .X(_02344_));
 sg13g2_nand3_1 _07445_ (.B(_02343_),
    .C(_02344_),
    .A(net17),
    .Y(_02345_));
 sg13g2_nand2_2 _07446_ (.Y(_02346_),
    .A(_02131_),
    .B(_02018_));
 sg13g2_nand2_1 _07447_ (.Y(_02347_),
    .A(net469),
    .B(net439));
 sg13g2_nand2b_1 _07448_ (.Y(_02348_),
    .B(_01981_),
    .A_N(net467));
 sg13g2_o21ai_1 _07449_ (.B1(_02348_),
    .Y(_02349_),
    .A1(net479),
    .A2(_02022_));
 sg13g2_a22oi_1 _07450_ (.Y(_02350_),
    .B1(_02022_),
    .B2(net479),
    .A2(_01979_),
    .A1(\median_processor.input_storage [26]));
 sg13g2_nand2_1 _07451_ (.Y(_02351_),
    .A(_02349_),
    .B(_02350_));
 sg13g2_nor2_1 _07452_ (.A(net418),
    .B(net389),
    .Y(_02352_));
 sg13g2_nand2b_1 _07453_ (.Y(_02353_),
    .B(net433),
    .A_N(net466));
 sg13g2_nand2b_1 _07454_ (.Y(_02354_),
    .B(_01967_),
    .A_N(net419));
 sg13g2_nand2b_1 _07455_ (.Y(_02355_),
    .B(_01978_),
    .A_N(\median_processor.input_storage [26]));
 sg13g2_nand3_1 _07456_ (.B(_02354_),
    .C(_02355_),
    .A(_02353_),
    .Y(_02356_));
 sg13g2_nor3_1 _07457_ (.A(\median_processor.input_storage [46]),
    .B(_02352_),
    .C(_02356_),
    .Y(_02357_));
 sg13g2_a221oi_1 _07458_ (.B2(net466),
    .C1(net419),
    .B1(_01977_),
    .A1(net418),
    .Y(_02358_),
    .A2(net389));
 sg13g2_nor2b_1 _07459_ (.A(_01984_),
    .B_N(net466),
    .Y(_02359_));
 sg13g2_a221oi_1 _07460_ (.B2(net419),
    .C1(net390),
    .B1(_02359_),
    .A1(net418),
    .Y(_02360_),
    .A2(net389));
 sg13g2_nor4_1 _07461_ (.A(\median_processor.input_storage [46]),
    .B(_02352_),
    .C(_02358_),
    .D(_02360_),
    .Y(_02361_));
 sg13g2_a21oi_1 _07462_ (.A1(_02351_),
    .A2(_02357_),
    .Y(_02362_),
    .B1(_02361_));
 sg13g2_a21oi_1 _07463_ (.A1(_02349_),
    .A2(_02350_),
    .Y(_02363_),
    .B1(_02356_));
 sg13g2_o21ai_1 _07464_ (.B1(\median_processor.input_storage [46]),
    .Y(_02364_),
    .A1(_02358_),
    .A2(_02360_));
 sg13g2_a21oi_1 _07465_ (.A1(net436),
    .A2(_02352_),
    .Y(_02365_),
    .B1(_01710_));
 sg13g2_o21ai_1 _07466_ (.B1(_02365_),
    .Y(_02366_),
    .A1(_02363_),
    .A2(_02364_));
 sg13g2_nand3_1 _07467_ (.B(_02362_),
    .C(_02366_),
    .A(_02347_),
    .Y(_02367_));
 sg13g2_nand2_2 _07468_ (.Y(_02368_),
    .A(_02346_),
    .B(_02367_));
 sg13g2_and2_1 _07469_ (.A(_02346_),
    .B(_02367_),
    .X(_02369_));
 sg13g2_buf_1 _07470_ (.A(_02369_),
    .X(_02370_));
 sg13g2_nand2_1 _07471_ (.Y(_02371_),
    .A(net446),
    .B(net432));
 sg13g2_nand2b_1 _07472_ (.Y(_02372_),
    .B(net448),
    .A_N(\median_processor.input_storage [40]));
 sg13g2_o21ai_1 _07473_ (.B1(_02372_),
    .Y(_02373_),
    .A1(_01882_),
    .A2(\median_processor.input_storage [41]));
 sg13g2_a22oi_1 _07474_ (.Y(_02374_),
    .B1(\median_processor.input_storage [41]),
    .B2(_01882_),
    .A2(\median_processor.input_storage [42]),
    .A1(_01880_));
 sg13g2_inv_1 _07475_ (.Y(_02375_),
    .A(net451));
 sg13g2_nand2b_1 _07476_ (.Y(_02376_),
    .B(net420),
    .A_N(\median_processor.input_storage [42]));
 sg13g2_nand2_1 _07477_ (.Y(_02377_),
    .A(_02375_),
    .B(_02376_));
 sg13g2_nand2_1 _07478_ (.Y(_02378_),
    .A(_01984_),
    .B(_02376_));
 sg13g2_a22oi_1 _07479_ (.Y(_02379_),
    .B1(_02377_),
    .B2(_02378_),
    .A2(_02374_),
    .A1(_02373_));
 sg13g2_a22oi_1 _07480_ (.Y(_02380_),
    .B1(_01967_),
    .B2(_02099_),
    .A2(net437),
    .A1(_01869_));
 sg13g2_o21ai_1 _07481_ (.B1(_02380_),
    .Y(_02381_),
    .A1(_01853_),
    .A2(_01977_));
 sg13g2_and2_1 _07482_ (.A(net450),
    .B(_01963_),
    .X(_02382_));
 sg13g2_nand2b_1 _07483_ (.Y(_02383_),
    .B(net450),
    .A_N(\median_processor.input_storage [44]));
 sg13g2_a21oi_1 _07484_ (.A1(net437),
    .A2(_02383_),
    .Y(_02384_),
    .B1(_01869_));
 sg13g2_nand2b_1 _07485_ (.Y(_02385_),
    .B(\median_processor.input_storage [55]),
    .A_N(\median_processor.input_storage [47]));
 sg13g2_nand2_1 _07486_ (.Y(_02386_),
    .A(\median_processor.input_storage [46]),
    .B(_02385_));
 sg13g2_nor3_1 _07487_ (.A(_02382_),
    .B(_02384_),
    .C(_02386_),
    .Y(_02387_));
 sg13g2_o21ai_1 _07488_ (.B1(_02387_),
    .Y(_02388_),
    .A1(_02379_),
    .A2(_02381_));
 sg13g2_nand2_1 _07489_ (.Y(_02389_),
    .A(_01865_),
    .B(_02385_));
 sg13g2_nor3_1 _07490_ (.A(_02382_),
    .B(_02384_),
    .C(_02389_),
    .Y(_02390_));
 sg13g2_o21ai_1 _07491_ (.B1(_02390_),
    .Y(_02391_),
    .A1(_02379_),
    .A2(_02381_));
 sg13g2_nand3_1 _07492_ (.B(\median_processor.input_storage [46]),
    .C(_02385_),
    .A(_01865_),
    .Y(_02392_));
 sg13g2_nand4_1 _07493_ (.B(_02388_),
    .C(_02391_),
    .A(_02371_),
    .Y(_02393_),
    .D(_02392_));
 sg13g2_buf_1 _07494_ (.A(_02393_),
    .X(_02394_));
 sg13g2_inv_1 _07495_ (.Y(_02395_),
    .A(net21));
 sg13g2_o21ai_1 _07496_ (.B1(_02395_),
    .Y(_02396_),
    .A1(_02012_),
    .A2(net16));
 sg13g2_o21ai_1 _07497_ (.B1(_02396_),
    .Y(_02397_),
    .A1(_01994_),
    .A2(_02368_));
 sg13g2_a21o_1 _07498_ (.A2(_02345_),
    .A1(_02342_),
    .B1(_02397_),
    .X(_02398_));
 sg13g2_nor3_1 _07499_ (.A(net17),
    .B(_02343_),
    .C(_02341_),
    .Y(_02399_));
 sg13g2_nand2_1 _07500_ (.Y(_02400_),
    .A(_02397_),
    .B(_02399_));
 sg13g2_xor2_1 _07501_ (.B(net21),
    .A(_01994_),
    .X(_02401_));
 sg13g2_xnor2_1 _07502_ (.Y(_02402_),
    .A(net14),
    .B(_02401_));
 sg13g2_nand2_1 _07503_ (.Y(_02403_),
    .A(net16),
    .B(_02402_));
 sg13g2_nand2b_1 _07504_ (.Y(_02404_),
    .B(_02368_),
    .A_N(_02402_));
 sg13g2_a22oi_1 _07505_ (.Y(_02405_),
    .B1(_02403_),
    .B2(_02404_),
    .A2(_02400_),
    .A1(_02398_));
 sg13g2_nand3_1 _07506_ (.B(_02289_),
    .C(_02341_),
    .A(net21),
    .Y(_02406_));
 sg13g2_nand2_1 _07507_ (.Y(_02407_),
    .A(_01994_),
    .B(_02343_));
 sg13g2_nor4_1 _07508_ (.A(net14),
    .B(net16),
    .C(_02406_),
    .D(_02407_),
    .Y(_02408_));
 sg13g2_and2_1 _07509_ (.A(net474),
    .B(\median_processor.input_storage [48]),
    .X(_02409_));
 sg13g2_nor2b_1 _07510_ (.A(\median_processor.input_storage [27]),
    .B_N(\median_processor.input_storage [51]),
    .Y(_02410_));
 sg13g2_a221oi_1 _07511_ (.B2(_02159_),
    .C1(_02410_),
    .B1(_02409_),
    .A1(net416),
    .Y(_02411_),
    .A2(\median_processor.input_storage [50]));
 sg13g2_nor2b_1 _07512_ (.A(_01725_),
    .B_N(_01859_),
    .Y(_02412_));
 sg13g2_o21ai_1 _07513_ (.B1(_01727_),
    .Y(_02413_),
    .A1(net474),
    .A2(_02412_));
 sg13g2_nor2_1 _07514_ (.A(net416),
    .B(net420),
    .Y(_02414_));
 sg13g2_nand2_1 _07515_ (.Y(_02415_),
    .A(net465),
    .B(\median_processor.input_storage [51]));
 sg13g2_nor2b_1 _07516_ (.A(\median_processor.input_storage [55]),
    .B_N(\median_processor.input_storage [31]),
    .Y(_02416_));
 sg13g2_nor2b_1 _07517_ (.A(\median_processor.input_storage [53]),
    .B_N(\median_processor.input_storage [29]),
    .Y(_02417_));
 sg13g2_nor2b_1 _07518_ (.A(\median_processor.input_storage [51]),
    .B_N(\median_processor.input_storage [27]),
    .Y(_02418_));
 sg13g2_nor2b_1 _07519_ (.A(\median_processor.input_storage [52]),
    .B_N(\median_processor.input_storage [28]),
    .Y(_02419_));
 sg13g2_or4_1 _07520_ (.A(_02416_),
    .B(_02417_),
    .C(_02418_),
    .D(_02419_),
    .X(_02420_));
 sg13g2_a221oi_1 _07521_ (.B2(_02415_),
    .C1(_02420_),
    .B1(_02414_),
    .A1(_02411_),
    .Y(_02421_),
    .A2(_02413_));
 sg13g2_buf_1 _07522_ (.A(\median_processor.input_storage [55]),
    .X(_02422_));
 sg13g2_nand2b_1 _07523_ (.Y(_02423_),
    .B(net450),
    .A_N(\median_processor.input_storage [28]));
 sg13g2_nand2b_1 _07524_ (.Y(_02424_),
    .B(_01857_),
    .A_N(\median_processor.input_storage [29]));
 sg13g2_a221oi_1 _07525_ (.B2(_02424_),
    .C1(_02417_),
    .B1(_02423_),
    .A1(_01707_),
    .Y(_02425_),
    .A2(net446));
 sg13g2_a21o_1 _07526_ (.A2(net447),
    .A1(net413),
    .B1(_02425_),
    .X(_02426_));
 sg13g2_o21ai_1 _07527_ (.B1(_01710_),
    .Y(_02427_),
    .A1(_02421_),
    .A2(_02426_));
 sg13g2_o21ai_1 _07528_ (.B1(_01867_),
    .Y(_02428_),
    .A1(net417),
    .A2(_01865_));
 sg13g2_and2_1 _07529_ (.A(net447),
    .B(_02425_),
    .X(_02429_));
 sg13g2_a221oi_1 _07530_ (.B2(_02131_),
    .C1(_02429_),
    .B1(_02428_),
    .A1(_01863_),
    .Y(_02430_),
    .A2(_02421_));
 sg13g2_nand2_2 _07531_ (.Y(_02431_),
    .A(_02427_),
    .B(_02430_));
 sg13g2_xnor2_1 _07532_ (.Y(_02432_),
    .A(_01895_),
    .B(_02431_));
 sg13g2_and2_1 _07533_ (.A(net21),
    .B(_02432_),
    .X(_02433_));
 sg13g2_and2_1 _07534_ (.A(_02427_),
    .B(_02430_),
    .X(_02434_));
 sg13g2_buf_2 _07535_ (.A(_02434_),
    .X(_02435_));
 sg13g2_nand2_1 _07536_ (.Y(_02436_),
    .A(_01895_),
    .B(_02435_));
 sg13g2_nor2_1 _07537_ (.A(net21),
    .B(_02436_),
    .Y(_02437_));
 sg13g2_nand2b_1 _07538_ (.Y(_02438_),
    .B(_01900_),
    .A_N(\median_processor.input_storage [55]));
 sg13g2_nand2b_1 _07539_ (.Y(_02439_),
    .B(\median_processor.input_storage [36]),
    .A_N(_01855_));
 sg13g2_nand2b_1 _07540_ (.Y(_02440_),
    .B(_01897_),
    .A_N(\median_processor.input_storage [54]));
 sg13g2_nand2b_1 _07541_ (.Y(_02441_),
    .B(net476),
    .A_N(\median_processor.input_storage [53]));
 sg13g2_nand4_1 _07542_ (.B(_02439_),
    .C(_02440_),
    .A(_02438_),
    .Y(_02442_),
    .D(_02441_));
 sg13g2_nor2_1 _07543_ (.A(_02326_),
    .B(_02104_),
    .Y(_02443_));
 sg13g2_nor3_1 _07544_ (.A(_02375_),
    .B(_02442_),
    .C(_02443_),
    .Y(_02444_));
 sg13g2_nor3_1 _07545_ (.A(_01910_),
    .B(_02442_),
    .C(_02443_),
    .Y(_02445_));
 sg13g2_a21oi_1 _07546_ (.A1(_01907_),
    .A2(_01859_),
    .Y(_02446_),
    .B1(\median_processor.input_storage [49]));
 sg13g2_a21oi_1 _07547_ (.A1(_01907_),
    .A2(_02409_),
    .Y(_02447_),
    .B1(_01908_));
 sg13g2_nand2_1 _07548_ (.Y(_02448_),
    .A(_02326_),
    .B(_02104_));
 sg13g2_o21ai_1 _07549_ (.B1(_02448_),
    .Y(_02449_),
    .A1(_02446_),
    .A2(_02447_));
 sg13g2_o21ai_1 _07550_ (.B1(_02449_),
    .Y(_02450_),
    .A1(_02444_),
    .A2(_02445_));
 sg13g2_nor2b_1 _07551_ (.A(\median_processor.input_storage [36]),
    .B_N(_01855_),
    .Y(_02451_));
 sg13g2_nand3_1 _07552_ (.B(_02440_),
    .C(_02451_),
    .A(net222),
    .Y(_02452_));
 sg13g2_nand2_1 _07553_ (.Y(_02453_),
    .A(_02189_),
    .B(_01853_));
 sg13g2_a21o_1 _07554_ (.A2(_02453_),
    .A1(_02452_),
    .B1(_02442_),
    .X(_02454_));
 sg13g2_nand2_1 _07555_ (.Y(_02455_),
    .A(net413),
    .B(_02440_));
 sg13g2_o21ai_1 _07556_ (.B1(_01901_),
    .Y(_02456_),
    .A1(net413),
    .A2(_02440_));
 sg13g2_nand2_1 _07557_ (.Y(_02457_),
    .A(_02455_),
    .B(_02456_));
 sg13g2_nand3_1 _07558_ (.B(_02441_),
    .C(_02451_),
    .A(_02422_),
    .Y(_02458_));
 sg13g2_a22oi_1 _07559_ (.Y(_02459_),
    .B1(_01857_),
    .B2(net443),
    .A2(_01863_),
    .A1(net392));
 sg13g2_nand2_1 _07560_ (.Y(_02460_),
    .A(_01901_),
    .B(_02422_));
 sg13g2_nand3_1 _07561_ (.B(_02459_),
    .C(_02460_),
    .A(_02458_),
    .Y(_02461_));
 sg13g2_nand2_1 _07562_ (.Y(_02462_),
    .A(_02457_),
    .B(_02461_));
 sg13g2_and3_1 _07563_ (.X(_02463_),
    .A(_02450_),
    .B(_02454_),
    .C(_02462_));
 sg13g2_buf_1 _07564_ (.A(_02463_),
    .X(_02464_));
 sg13g2_nor2_2 _07565_ (.A(net413),
    .B(net394),
    .Y(_02465_));
 sg13g2_nand2_1 _07566_ (.Y(_02466_),
    .A(\median_processor.input_storage [57]),
    .B(\median_processor.input_storage [56]));
 sg13g2_o21ai_1 _07567_ (.B1(net474),
    .Y(_02467_),
    .A1(net448),
    .A2(_02466_));
 sg13g2_nand2b_1 _07568_ (.Y(_02468_),
    .B(\median_processor.input_storage [56]),
    .A_N(net448));
 sg13g2_a221oi_1 _07569_ (.B2(_02468_),
    .C1(_02210_),
    .B1(net458),
    .A1(net420),
    .Y(_02469_),
    .A2(_01814_));
 sg13g2_nand2b_1 _07570_ (.Y(_02470_),
    .B(net454),
    .A_N(net420));
 sg13g2_a21oi_1 _07571_ (.A1(net451),
    .A2(_02210_),
    .Y(_02471_),
    .B1(_02470_));
 sg13g2_a21oi_1 _07572_ (.A1(_02467_),
    .A2(_02469_),
    .Y(_02472_),
    .B1(_02471_));
 sg13g2_a221oi_1 _07573_ (.B2(_02468_),
    .C1(net451),
    .B1(net458),
    .A1(net420),
    .Y(_02473_),
    .A2(_01814_));
 sg13g2_a22oi_1 _07574_ (.Y(_02474_),
    .B1(_02467_),
    .B2(_02473_),
    .A2(net453),
    .A1(_02375_));
 sg13g2_nand2_1 _07575_ (.Y(_02475_),
    .A(net449),
    .B(net395));
 sg13g2_nand2_1 _07576_ (.Y(_02476_),
    .A(\median_processor.input_storage [60]),
    .B(_02475_));
 sg13g2_nand2_1 _07577_ (.Y(_02477_),
    .A(_02099_),
    .B(_02475_));
 sg13g2_a22oi_1 _07578_ (.Y(_02478_),
    .B1(_02476_),
    .B2(_02477_),
    .A2(_02474_),
    .A1(_02472_));
 sg13g2_nand3_1 _07579_ (.B(\median_processor.input_storage [60]),
    .C(_02475_),
    .A(_02099_),
    .Y(_02479_));
 sg13g2_o21ai_1 _07580_ (.B1(_02479_),
    .Y(_02480_),
    .A1(net449),
    .A2(net395));
 sg13g2_o21ai_1 _07581_ (.B1(net388),
    .Y(_02481_),
    .A1(_02478_),
    .A2(_02480_));
 sg13g2_nor3_1 _07582_ (.A(_02223_),
    .B(_02478_),
    .C(_02480_),
    .Y(_02482_));
 sg13g2_a221oi_1 _07583_ (.B2(net447),
    .C1(_02482_),
    .B1(_02481_),
    .A1(net413),
    .Y(_02483_),
    .A2(net394));
 sg13g2_nor3_1 _07584_ (.A(net20),
    .B(_02465_),
    .C(_02483_),
    .Y(_02484_));
 sg13g2_o21ai_1 _07585_ (.B1(_02484_),
    .Y(_02485_),
    .A1(_02433_),
    .A2(_02437_));
 sg13g2_nand2b_1 _07586_ (.Y(_02486_),
    .B(_02431_),
    .A_N(_01895_));
 sg13g2_o21ai_1 _07587_ (.B1(net20),
    .Y(_02487_),
    .A1(_02465_),
    .A2(_02483_));
 sg13g2_or3_1 _07588_ (.A(net21),
    .B(_02486_),
    .C(_02487_),
    .X(_02488_));
 sg13g2_nand2_1 _07589_ (.Y(_02489_),
    .A(net423),
    .B(_02099_));
 sg13g2_nand2_1 _07590_ (.Y(_02490_),
    .A(net478),
    .B(_01880_));
 sg13g2_nand3_1 _07591_ (.B(_02489_),
    .C(_02490_),
    .A(net451),
    .Y(_02491_));
 sg13g2_nand3_1 _07592_ (.B(_02489_),
    .C(_02490_),
    .A(_01763_),
    .Y(_02492_));
 sg13g2_nand2b_1 _07593_ (.Y(_02493_),
    .B(net448),
    .A_N(net484));
 sg13g2_o21ai_1 _07594_ (.B1(_01882_),
    .Y(_02494_),
    .A1(\median_processor.input_storage [1]),
    .A2(_02493_));
 sg13g2_nand2_1 _07595_ (.Y(_02495_),
    .A(\median_processor.input_storage [1]),
    .B(_02493_));
 sg13g2_a22oi_1 _07596_ (.Y(_02496_),
    .B1(_02494_),
    .B2(_02495_),
    .A2(net420),
    .A1(net425));
 sg13g2_a21o_1 _07597_ (.A2(_02492_),
    .A1(_02491_),
    .B1(_02496_),
    .X(_02497_));
 sg13g2_nor2_1 _07598_ (.A(net461),
    .B(_02375_),
    .Y(_02498_));
 sg13g2_nor2_1 _07599_ (.A(net423),
    .B(_02099_),
    .Y(_02499_));
 sg13g2_a21oi_1 _07600_ (.A1(_02489_),
    .A2(_02498_),
    .Y(_02500_),
    .B1(_02499_));
 sg13g2_a22oi_1 _07601_ (.Y(_02501_),
    .B1(_01865_),
    .B2(net440),
    .A2(net446),
    .A1(net472));
 sg13g2_nand2_1 _07602_ (.Y(_02502_),
    .A(net449),
    .B(_02501_));
 sg13g2_nand2_1 _07603_ (.Y(_02503_),
    .A(_01762_),
    .B(_02501_));
 sg13g2_a22oi_1 _07604_ (.Y(_02504_),
    .B1(_02502_),
    .B2(_02503_),
    .A2(_02500_),
    .A1(_02497_));
 sg13g2_nor2_1 _07605_ (.A(_01946_),
    .B(_01865_),
    .Y(_02505_));
 sg13g2_nand2_1 _07606_ (.Y(_02506_),
    .A(net413),
    .B(_02505_));
 sg13g2_o21ai_1 _07607_ (.B1(_01808_),
    .Y(_02507_),
    .A1(net413),
    .A2(_02505_));
 sg13g2_nand3_1 _07608_ (.B(net449),
    .C(_02501_),
    .A(_01762_),
    .Y(_02508_));
 sg13g2_nand3_1 _07609_ (.B(_02507_),
    .C(_02508_),
    .A(_02506_),
    .Y(_02509_));
 sg13g2_o21ai_1 _07610_ (.B1(_02129_),
    .Y(_02510_),
    .A1(_02504_),
    .A2(_02509_));
 sg13g2_nor2_2 _07611_ (.A(_02504_),
    .B(_02509_),
    .Y(_02511_));
 sg13g2_nand2_1 _07612_ (.Y(_02512_),
    .A(_02251_),
    .B(_02511_));
 sg13g2_nand2_1 _07613_ (.Y(_02513_),
    .A(_02510_),
    .B(_02512_));
 sg13g2_a21oi_1 _07614_ (.A1(_02485_),
    .A2(_02488_),
    .Y(_02514_),
    .B1(_02513_));
 sg13g2_o21ai_1 _07615_ (.B1(net21),
    .Y(_02515_),
    .A1(_01895_),
    .A2(_02435_));
 sg13g2_nand2_1 _07616_ (.Y(_02516_),
    .A(_02436_),
    .B(_02515_));
 sg13g2_mux2_1 _07617_ (.A0(_02512_),
    .A1(_02510_),
    .S(_02516_),
    .X(_02517_));
 sg13g2_or2_1 _07618_ (.X(_02518_),
    .B(_02465_),
    .A(net20));
 sg13g2_nor2_1 _07619_ (.A(net446),
    .B(net473),
    .Y(_02519_));
 sg13g2_nand2b_1 _07620_ (.Y(_02520_),
    .B(net20),
    .A_N(_02519_));
 sg13g2_a21oi_1 _07621_ (.A1(net447),
    .A2(_02481_),
    .Y(_02521_),
    .B1(_02482_));
 sg13g2_mux2_1 _07622_ (.A0(_02518_),
    .A1(_02520_),
    .S(_02521_),
    .X(_02522_));
 sg13g2_nand3_1 _07623_ (.B(_02454_),
    .C(_02462_),
    .A(_02450_),
    .Y(_02523_));
 sg13g2_mux2_1 _07624_ (.A0(_02465_),
    .A1(_02519_),
    .S(_02523_),
    .X(_02524_));
 sg13g2_inv_1 _07625_ (.Y(_02525_),
    .A(_02524_));
 sg13g2_xnor2_1 _07626_ (.Y(_02526_),
    .A(_02395_),
    .B(_02432_));
 sg13g2_a21oi_1 _07627_ (.A1(_02522_),
    .A2(_02525_),
    .Y(_02527_),
    .B1(_02526_));
 sg13g2_nor2b_1 _07628_ (.A(_02484_),
    .B_N(_02526_),
    .Y(_02528_));
 sg13g2_nor3_1 _07629_ (.A(_02517_),
    .B(_02527_),
    .C(_02528_),
    .Y(_02529_));
 sg13g2_nand2_1 _07630_ (.Y(_02530_),
    .A(_02395_),
    .B(_02432_));
 sg13g2_or2_1 _07631_ (.X(_02531_),
    .B(_02486_),
    .A(_02395_));
 sg13g2_or2_1 _07632_ (.X(_02532_),
    .B(_02487_),
    .A(_02510_));
 sg13g2_nand4_1 _07633_ (.B(_02512_),
    .C(_02522_),
    .A(_02510_),
    .Y(_02533_),
    .D(_02525_));
 sg13g2_a22oi_1 _07634_ (.Y(_02534_),
    .B1(_02532_),
    .B2(_02533_),
    .A2(_02531_),
    .A1(_02530_));
 sg13g2_or3_1 _07635_ (.A(_02514_),
    .B(_02529_),
    .C(_02534_),
    .X(_02535_));
 sg13g2_buf_2 _07636_ (.A(_02535_),
    .X(_02536_));
 sg13g2_nand2_1 _07637_ (.Y(_02537_),
    .A(_02322_),
    .B(_02344_));
 sg13g2_nand3b_1 _07638_ (.B(_02321_),
    .C(_02341_),
    .Y(_02538_),
    .A_N(_02289_));
 sg13g2_and3_1 _07639_ (.X(_02539_),
    .A(_01994_),
    .B(net14),
    .C(net16));
 sg13g2_xnor2_1 _07640_ (.Y(_02540_),
    .A(_02048_),
    .B(_02368_));
 sg13g2_nor4_1 _07641_ (.A(_01994_),
    .B(_02048_),
    .C(net21),
    .D(net16),
    .Y(_02541_));
 sg13g2_a221oi_1 _07642_ (.B2(_02401_),
    .C1(_02541_),
    .B1(_02540_),
    .A1(_02394_),
    .Y(_02542_),
    .A2(_02539_));
 sg13g2_a21oi_1 _07643_ (.A1(_02537_),
    .A2(_02538_),
    .Y(_02543_),
    .B1(_02542_));
 sg13g2_or4_1 _07644_ (.A(_02405_),
    .B(_02408_),
    .C(_02536_),
    .D(_02543_),
    .X(_02544_));
 sg13g2_buf_1 _07645_ (.A(_02544_),
    .X(_02545_));
 sg13g2_buf_1 _07646_ (.A(net4),
    .X(_02546_));
 sg13g2_nor2_1 _07647_ (.A(net434),
    .B(_02536_),
    .Y(_02547_));
 sg13g2_a21oi_1 _07648_ (.A1(_01876_),
    .A2(_02536_),
    .Y(_02548_),
    .B1(_02547_));
 sg13g2_nand2b_1 _07649_ (.Y(_02549_),
    .B(_02017_),
    .A_N(_02466_));
 sg13g2_nor2b_1 _07650_ (.A(net484),
    .B_N(_01818_),
    .Y(_02550_));
 sg13g2_o21ai_1 _07651_ (.B1(_02055_),
    .Y(_02551_),
    .A1(\median_processor.input_storage [57]),
    .A2(_02550_));
 sg13g2_nor2_1 _07652_ (.A(_01763_),
    .B(net453),
    .Y(_02552_));
 sg13g2_a221oi_1 _07653_ (.B2(_02551_),
    .C1(_02552_),
    .B1(_02549_),
    .A1(net478),
    .Y(_02553_),
    .A2(_01814_));
 sg13g2_nand2_1 _07654_ (.Y(_02554_),
    .A(net425),
    .B(net454));
 sg13g2_nand2_1 _07655_ (.Y(_02555_),
    .A(_01763_),
    .B(net453));
 sg13g2_o21ai_1 _07656_ (.B1(_02555_),
    .Y(_02556_),
    .A1(_02552_),
    .A2(_02554_));
 sg13g2_nand2b_1 _07657_ (.Y(_02557_),
    .B(net472),
    .A_N(net473));
 sg13g2_nand2b_1 _07658_ (.Y(_02558_),
    .B(net440),
    .A_N(net452));
 sg13g2_nand2b_1 _07659_ (.Y(_02559_),
    .B(net422),
    .A_N(net455));
 sg13g2_nand3_1 _07660_ (.B(_02558_),
    .C(_02559_),
    .A(_02557_),
    .Y(_02560_));
 sg13g2_nor2_1 _07661_ (.A(net387),
    .B(_02560_),
    .Y(_02561_));
 sg13g2_o21ai_1 _07662_ (.B1(_02561_),
    .Y(_02562_),
    .A1(_02553_),
    .A2(_02556_));
 sg13g2_nor2_1 _07663_ (.A(net423),
    .B(_02560_),
    .Y(_02563_));
 sg13g2_o21ai_1 _07664_ (.B1(_02563_),
    .Y(_02564_),
    .A1(_02553_),
    .A2(_02556_));
 sg13g2_nor2b_1 _07665_ (.A(net422),
    .B_N(net455),
    .Y(_02565_));
 sg13g2_o21ai_1 _07666_ (.B1(net388),
    .Y(_02566_),
    .A1(net462),
    .A2(_02565_));
 sg13g2_nand2_1 _07667_ (.Y(_02567_),
    .A(net462),
    .B(_02565_));
 sg13g2_a22oi_1 _07668_ (.Y(_02568_),
    .B1(_02566_),
    .B2(_02567_),
    .A2(net394),
    .A1(net472));
 sg13g2_nor2_1 _07669_ (.A(net472),
    .B(net394),
    .Y(_02569_));
 sg13g2_nor3_1 _07670_ (.A(net423),
    .B(net387),
    .C(_02560_),
    .Y(_02570_));
 sg13g2_nor3_1 _07671_ (.A(_02568_),
    .B(_02569_),
    .C(_02570_),
    .Y(_02571_));
 sg13g2_nand3_1 _07672_ (.B(_02564_),
    .C(_02571_),
    .A(_02562_),
    .Y(_02572_));
 sg13g2_and2_1 _07673_ (.A(_02226_),
    .B(_02572_),
    .X(_02573_));
 sg13g2_nor2_1 _07674_ (.A(_02226_),
    .B(_02572_),
    .Y(_02574_));
 sg13g2_or2_1 _07675_ (.X(_02575_),
    .B(_02574_),
    .A(_02573_));
 sg13g2_nor2_1 _07676_ (.A(net476),
    .B(net395),
    .Y(_02576_));
 sg13g2_nand2_1 _07677_ (.Y(_02577_),
    .A(net452),
    .B(_01823_));
 sg13g2_o21ai_1 _07678_ (.B1(net445),
    .Y(_02578_),
    .A1(net476),
    .A2(_02577_));
 sg13g2_o21ai_1 _07679_ (.B1(_02578_),
    .Y(_02579_),
    .A1(_02223_),
    .A2(_02576_));
 sg13g2_o21ai_1 _07680_ (.B1(_02579_),
    .Y(_02580_),
    .A1(net444),
    .A2(net394));
 sg13g2_nand2_1 _07681_ (.Y(_02581_),
    .A(net444),
    .B(_01847_));
 sg13g2_nand2b_1 _07682_ (.Y(_02582_),
    .B(_01818_),
    .A_N(net477));
 sg13g2_a21oi_1 _07683_ (.A1(net414),
    .A2(_02582_),
    .Y(_02583_),
    .B1(_01817_));
 sg13g2_nor2_1 _07684_ (.A(net414),
    .B(_02582_),
    .Y(_02584_));
 sg13g2_nand2_1 _07685_ (.Y(_02585_),
    .A(net441),
    .B(_01814_));
 sg13g2_o21ai_1 _07686_ (.B1(_02585_),
    .Y(_02586_),
    .A1(_02583_),
    .A2(_02584_));
 sg13g2_nor2_1 _07687_ (.A(net415),
    .B(net387),
    .Y(_02587_));
 sg13g2_a221oi_1 _07688_ (.B2(_02326_),
    .C1(_02587_),
    .B1(net454),
    .A1(_02189_),
    .Y(_02588_),
    .A2(net453));
 sg13g2_nand2b_1 _07689_ (.Y(_02589_),
    .B(net476),
    .A_N(_01823_));
 sg13g2_nand2b_1 _07690_ (.Y(_02590_),
    .B(net445),
    .A_N(\median_processor.input_storage [62]));
 sg13g2_nand3_1 _07691_ (.B(_02589_),
    .C(_02590_),
    .A(net473),
    .Y(_02591_));
 sg13g2_a21oi_1 _07692_ (.A1(net392),
    .A2(net452),
    .Y(_02592_),
    .B1(_02589_));
 sg13g2_o21ai_1 _07693_ (.B1(net222),
    .Y(_02593_),
    .A1(\median_processor.input_storage [63]),
    .A2(_02590_));
 sg13g2_a21o_1 _07694_ (.A2(_02592_),
    .A1(_01846_),
    .B1(_02593_),
    .X(_02594_));
 sg13g2_nor2b_1 _07695_ (.A(_01834_),
    .B_N(net442),
    .Y(_02595_));
 sg13g2_nor2_1 _07696_ (.A(net387),
    .B(_02595_),
    .Y(_02596_));
 sg13g2_a21oi_1 _07697_ (.A1(net387),
    .A2(_02595_),
    .Y(_02597_),
    .B1(net415));
 sg13g2_nor2_1 _07698_ (.A(_02596_),
    .B(_02597_),
    .Y(_02598_));
 sg13g2_a221oi_1 _07699_ (.B2(_02594_),
    .C1(_02598_),
    .B1(_02591_),
    .A1(_02586_),
    .Y(_02599_),
    .A2(_02588_));
 sg13g2_a21oi_2 _07700_ (.B1(_02599_),
    .Y(_02600_),
    .A2(_02581_),
    .A1(_02580_));
 sg13g2_nor2_1 _07701_ (.A(_02343_),
    .B(_02600_),
    .Y(_02601_));
 sg13g2_a21o_2 _07702_ (.A2(_02581_),
    .A1(_02580_),
    .B1(_02599_),
    .X(_02602_));
 sg13g2_nor2_1 _07703_ (.A(_02321_),
    .B(_02602_),
    .Y(_02603_));
 sg13g2_nor2_1 _07704_ (.A(_02601_),
    .B(_02603_),
    .Y(_02604_));
 sg13g2_nor2_1 _07705_ (.A(_02321_),
    .B(_02600_),
    .Y(_02605_));
 sg13g2_nor2_1 _07706_ (.A(_02343_),
    .B(_02602_),
    .Y(_02606_));
 sg13g2_a22oi_1 _07707_ (.Y(_02607_),
    .B1(_02606_),
    .B2(_02573_),
    .A2(_02574_),
    .A1(_02605_));
 sg13g2_o21ai_1 _07708_ (.B1(_02607_),
    .Y(_02608_),
    .A1(_02575_),
    .A2(_02604_));
 sg13g2_nand2_1 _07709_ (.Y(_02609_),
    .A(net469),
    .B(_01846_));
 sg13g2_nor2_1 _07710_ (.A(net418),
    .B(_01833_),
    .Y(_02610_));
 sg13g2_o21ai_1 _07711_ (.B1(net417),
    .Y(_02611_),
    .A1(net418),
    .A2(_02577_));
 sg13g2_o21ai_1 _07712_ (.B1(_02611_),
    .Y(_02612_),
    .A1(_01843_),
    .A2(_02610_));
 sg13g2_o21ai_1 _07713_ (.B1(_02612_),
    .Y(_02613_),
    .A1(net469),
    .A2(net394));
 sg13g2_nor2_1 _07714_ (.A(net416),
    .B(_01825_),
    .Y(_02614_));
 sg13g2_inv_1 _07715_ (.Y(_02615_),
    .A(net457));
 sg13g2_o21ai_1 _07716_ (.B1(net479),
    .Y(_02616_),
    .A1(net467),
    .A2(_02615_));
 sg13g2_or2_1 _07717_ (.X(_02617_),
    .B(net467),
    .A(net479));
 sg13g2_o21ai_1 _07718_ (.B1(_01817_),
    .Y(_02618_),
    .A1(_02615_),
    .A2(_02617_));
 sg13g2_a22oi_1 _07719_ (.Y(_02619_),
    .B1(_02616_),
    .B2(_02618_),
    .A2(_01825_),
    .A1(net416));
 sg13g2_nand2_1 _07720_ (.Y(_02620_),
    .A(net465),
    .B(_01834_));
 sg13g2_o21ai_1 _07721_ (.B1(_02620_),
    .Y(_02621_),
    .A1(_02614_),
    .A2(_02619_));
 sg13g2_nand2b_1 _07722_ (.Y(_02622_),
    .B(net417),
    .A_N(_01843_));
 sg13g2_nand2_1 _07723_ (.Y(_02623_),
    .A(net418),
    .B(_01833_));
 sg13g2_nand3_1 _07724_ (.B(_02622_),
    .C(_02623_),
    .A(_02609_),
    .Y(_02624_));
 sg13g2_a221oi_1 _07725_ (.B2(net466),
    .C1(_02624_),
    .B1(_02210_),
    .A1(net419),
    .Y(_02625_),
    .A2(_02306_));
 sg13g2_nor3_1 _07726_ (.A(net419),
    .B(_02306_),
    .C(_02624_),
    .Y(_02626_));
 sg13g2_a221oi_1 _07727_ (.B2(_02625_),
    .C1(_02626_),
    .B1(_02621_),
    .A1(_02609_),
    .Y(_02627_),
    .A2(_02613_));
 sg13g2_buf_1 _07728_ (.A(_02627_),
    .X(_02628_));
 sg13g2_nor2_1 _07729_ (.A(net25),
    .B(net19),
    .Y(_02629_));
 sg13g2_nand2_1 _07730_ (.Y(_02630_),
    .A(_02608_),
    .B(_02629_));
 sg13g2_or2_1 _07731_ (.X(_02631_),
    .B(_02483_),
    .A(_02465_));
 sg13g2_o21ai_1 _07732_ (.B1(_02573_),
    .Y(_02632_),
    .A1(_02601_),
    .A2(_02603_));
 sg13g2_nor2_1 _07733_ (.A(_02573_),
    .B(_02574_),
    .Y(_02633_));
 sg13g2_nand2_1 _07734_ (.Y(_02634_),
    .A(_02605_),
    .B(_02633_));
 sg13g2_xnor2_1 _07735_ (.Y(_02635_),
    .A(net25),
    .B(net19));
 sg13g2_a21oi_1 _07736_ (.A1(_02632_),
    .A2(_02634_),
    .Y(_02636_),
    .B1(_02635_));
 sg13g2_and2_1 _07737_ (.A(net25),
    .B(net19),
    .X(_02637_));
 sg13g2_nand2_1 _07738_ (.Y(_02638_),
    .A(_02573_),
    .B(_02637_));
 sg13g2_nor3_1 _07739_ (.A(_02321_),
    .B(_02600_),
    .C(_02638_),
    .Y(_02639_));
 sg13g2_nor3_1 _07740_ (.A(_02631_),
    .B(_02636_),
    .C(_02639_),
    .Y(_02640_));
 sg13g2_a22oi_1 _07741_ (.Y(_02641_),
    .B1(_02637_),
    .B2(_02605_),
    .A2(_02629_),
    .A1(_02606_));
 sg13g2_o21ai_1 _07742_ (.B1(_02641_),
    .Y(_02642_),
    .A1(_02635_),
    .A2(_02604_));
 sg13g2_nand2_1 _07743_ (.Y(_02643_),
    .A(_02633_),
    .B(_02642_));
 sg13g2_nand2_1 _07744_ (.Y(_02644_),
    .A(_02574_),
    .B(_02629_));
 sg13g2_a21oi_1 _07745_ (.A1(_02638_),
    .A2(_02644_),
    .Y(_02645_),
    .B1(_02604_));
 sg13g2_o21ai_1 _07746_ (.B1(_02631_),
    .Y(_02646_),
    .A1(_02635_),
    .A2(_02607_));
 sg13g2_nor2_1 _07747_ (.A(_02645_),
    .B(_02646_),
    .Y(_02647_));
 sg13g2_a22oi_1 _07748_ (.Y(_02648_),
    .B1(_02643_),
    .B2(_02647_),
    .A2(_02640_),
    .A1(_02630_));
 sg13g2_a21oi_1 _07749_ (.A1(_02017_),
    .A2(net477),
    .Y(_02649_),
    .B1(net414));
 sg13g2_nand2b_1 _07750_ (.Y(_02650_),
    .B(net478),
    .A_N(net441));
 sg13g2_nand2_1 _07751_ (.Y(_02651_),
    .A(_02055_),
    .B(_02650_));
 sg13g2_nand4_1 _07752_ (.B(net414),
    .C(net477),
    .A(_02017_),
    .Y(_02652_),
    .D(_02650_));
 sg13g2_o21ai_1 _07753_ (.B1(_02652_),
    .Y(_02653_),
    .A1(_02649_),
    .A2(_02651_));
 sg13g2_a221oi_1 _07754_ (.B2(net425),
    .C1(_02653_),
    .B1(net441),
    .A1(_01763_),
    .Y(_02654_),
    .A2(net442));
 sg13g2_inv_1 _07755_ (.Y(_02655_),
    .A(net415));
 sg13g2_a22oi_1 _07756_ (.Y(_02656_),
    .B1(_02655_),
    .B2(net423),
    .A2(net443),
    .A1(net422));
 sg13g2_o21ai_1 _07757_ (.B1(_02656_),
    .Y(_02657_),
    .A1(_01763_),
    .A2(net442));
 sg13g2_nand2_1 _07758_ (.Y(_02658_),
    .A(_01808_),
    .B(net444));
 sg13g2_nand2b_1 _07759_ (.Y(_02659_),
    .B(net415),
    .A_N(_02059_));
 sg13g2_nor2_1 _07760_ (.A(net443),
    .B(_02659_),
    .Y(_02660_));
 sg13g2_a21oi_1 _07761_ (.A1(net443),
    .A2(_02659_),
    .Y(_02661_),
    .B1(net422));
 sg13g2_nor2_1 _07762_ (.A(_02660_),
    .B(_02661_),
    .Y(_02662_));
 sg13g2_and3_1 _07763_ (.X(_02663_),
    .A(net392),
    .B(_02658_),
    .C(_02662_));
 sg13g2_o21ai_1 _07764_ (.B1(_02663_),
    .Y(_02664_),
    .A1(_02654_),
    .A2(_02657_));
 sg13g2_and3_1 _07765_ (.X(_02665_),
    .A(net440),
    .B(_02658_),
    .C(_02662_));
 sg13g2_o21ai_1 _07766_ (.B1(_02665_),
    .Y(_02666_),
    .A1(_02654_),
    .A2(_02657_));
 sg13g2_nor2_1 _07767_ (.A(net462),
    .B(net445),
    .Y(_02667_));
 sg13g2_nor2_1 _07768_ (.A(_01944_),
    .B(net444),
    .Y(_02668_));
 sg13g2_a21oi_1 _07769_ (.A1(_02658_),
    .A2(_02667_),
    .Y(_02669_),
    .B1(_02668_));
 sg13g2_nand3_1 _07770_ (.B(_02666_),
    .C(_02669_),
    .A(_02664_),
    .Y(_02670_));
 sg13g2_buf_1 _07771_ (.A(_02670_),
    .X(_02671_));
 sg13g2_o21ai_1 _07772_ (.B1(net222),
    .Y(_02672_),
    .A1(_02141_),
    .A2(net392));
 sg13g2_nor2_1 _07773_ (.A(_02141_),
    .B(_01929_),
    .Y(_02673_));
 sg13g2_a21o_1 _07774_ (.A2(_02673_),
    .A1(_01900_),
    .B1(_02131_),
    .X(_02674_));
 sg13g2_nor2b_1 _07775_ (.A(_01897_),
    .B_N(\median_processor.input_storage [30]),
    .Y(_02675_));
 sg13g2_a221oi_1 _07776_ (.B2(\median_processor.input_storage [29]),
    .C1(_02675_),
    .B1(_01904_),
    .A1(_01707_),
    .Y(_02676_),
    .A2(_01902_));
 sg13g2_nand2b_1 _07777_ (.Y(_02677_),
    .B(\median_processor.input_storage [26]),
    .A_N(_01912_));
 sg13g2_o21ai_1 _07778_ (.B1(_01910_),
    .Y(_02678_),
    .A1(net465),
    .A2(_02677_));
 sg13g2_nand2_1 _07779_ (.Y(_02679_),
    .A(net465),
    .B(_02677_));
 sg13g2_nor2b_1 _07780_ (.A(_01725_),
    .B_N(\median_processor.input_storage [32]),
    .Y(_02680_));
 sg13g2_nor2b_1 _07781_ (.A(_01730_),
    .B_N(\median_processor.input_storage [35]),
    .Y(_02681_));
 sg13g2_a221oi_1 _07782_ (.B2(_02680_),
    .C1(_02681_),
    .B1(_02177_),
    .A1(net416),
    .Y(_02682_),
    .A2(_01912_));
 sg13g2_o21ai_1 _07783_ (.B1(_01727_),
    .Y(_02683_),
    .A1(_02177_),
    .A2(_02680_));
 sg13g2_inv_1 _07784_ (.Y(_02684_),
    .A(_02133_));
 sg13g2_nor2_1 _07785_ (.A(_02684_),
    .B(_02168_),
    .Y(_02685_));
 sg13g2_a221oi_1 _07786_ (.B2(_02683_),
    .C1(_02685_),
    .B1(_02682_),
    .A1(_02678_),
    .Y(_02686_),
    .A2(_02679_));
 sg13g2_inv_1 _07787_ (.Y(_02687_),
    .A(net418));
 sg13g2_a22oi_1 _07788_ (.Y(_02688_),
    .B1(_02168_),
    .B2(_02684_),
    .A2(\median_processor.input_storage [37]),
    .A1(_02687_));
 sg13g2_nor2b_1 _07789_ (.A(_02688_),
    .B_N(_02676_),
    .Y(_02689_));
 sg13g2_a221oi_1 _07790_ (.B2(_02686_),
    .C1(_02689_),
    .B1(_02676_),
    .A1(_02672_),
    .Y(_02690_),
    .A2(_02674_));
 sg13g2_and2_1 _07791_ (.A(_01935_),
    .B(_02690_),
    .X(_02691_));
 sg13g2_nor2_1 _07792_ (.A(_02523_),
    .B(_02602_),
    .Y(_02692_));
 sg13g2_xnor2_1 _07793_ (.Y(_02693_),
    .A(_01943_),
    .B(_02690_));
 sg13g2_xnor2_1 _07794_ (.Y(_02694_),
    .A(_02523_),
    .B(_02600_));
 sg13g2_or3_1 _07795_ (.A(_01920_),
    .B(_01934_),
    .C(_02690_),
    .X(_02695_));
 sg13g2_nor3_1 _07796_ (.A(net20),
    .B(_02600_),
    .C(_02695_),
    .Y(_02696_));
 sg13g2_a221oi_1 _07797_ (.B2(_02694_),
    .C1(_02696_),
    .B1(_02693_),
    .A1(_02691_),
    .Y(_02697_),
    .A2(_02692_));
 sg13g2_nor2_1 _07798_ (.A(net15),
    .B(_02697_),
    .Y(_02698_));
 sg13g2_nor2_1 _07799_ (.A(_02239_),
    .B(_02697_),
    .Y(_02699_));
 sg13g2_nor2_1 _07800_ (.A(net20),
    .B(_02600_),
    .Y(_02700_));
 sg13g2_nor2_1 _07801_ (.A(net20),
    .B(_02602_),
    .Y(_02701_));
 sg13g2_and4_1 _07802_ (.A(_01935_),
    .B(_02464_),
    .C(_02602_),
    .D(_02690_),
    .X(_02702_));
 sg13g2_a221oi_1 _07803_ (.B2(_02691_),
    .C1(_02702_),
    .B1(_02701_),
    .A1(_02700_),
    .Y(_02703_),
    .A2(_02693_));
 sg13g2_nor3_1 _07804_ (.A(_02239_),
    .B(net15),
    .C(_02703_),
    .Y(_02704_));
 sg13g2_a221oi_1 _07805_ (.B2(net15),
    .C1(_02704_),
    .B1(_02699_),
    .A1(_02239_),
    .Y(_02705_),
    .A2(_02698_));
 sg13g2_nor2_1 _07806_ (.A(_02602_),
    .B(_02695_),
    .Y(_02706_));
 sg13g2_nor3_1 _07807_ (.A(_02523_),
    .B(_02600_),
    .C(_02695_),
    .Y(_02707_));
 sg13g2_a221oi_1 _07808_ (.B2(_02523_),
    .C1(_02707_),
    .B1(_02706_),
    .A1(_02692_),
    .Y(_02708_),
    .A2(_02693_));
 sg13g2_nand2_1 _07809_ (.Y(_02709_),
    .A(_02239_),
    .B(_02671_));
 sg13g2_nor3_1 _07810_ (.A(_02344_),
    .B(_02708_),
    .C(_02709_),
    .Y(_02710_));
 sg13g2_xnor2_1 _07811_ (.Y(_02711_),
    .A(_02239_),
    .B(_02670_));
 sg13g2_nor3_1 _07812_ (.A(_02341_),
    .B(_02708_),
    .C(_02711_),
    .Y(_02712_));
 sg13g2_nor4_1 _07813_ (.A(_02239_),
    .B(_02341_),
    .C(_02671_),
    .D(_02697_),
    .Y(_02713_));
 sg13g2_nand2_1 _07814_ (.Y(_02714_),
    .A(net20),
    .B(_02600_));
 sg13g2_nor4_1 _07815_ (.A(_02341_),
    .B(_02714_),
    .C(_02695_),
    .D(_02709_),
    .Y(_02715_));
 sg13g2_nor4_1 _07816_ (.A(_02710_),
    .B(_02712_),
    .C(_02713_),
    .D(_02715_),
    .Y(_02716_));
 sg13g2_o21ai_1 _07817_ (.B1(_02716_),
    .Y(_02717_),
    .A1(_02344_),
    .A2(_02705_));
 sg13g2_buf_1 _07818_ (.A(_02717_),
    .X(_02718_));
 sg13g2_xor2_1 _07819_ (.B(_02690_),
    .A(_01749_),
    .X(_02719_));
 sg13g2_xnor2_1 _07820_ (.Y(_02720_),
    .A(_02435_),
    .B(_02719_));
 sg13g2_nor2b_1 _07821_ (.A(_01946_),
    .B_N(net417),
    .Y(_02721_));
 sg13g2_nor2b_1 _07822_ (.A(_02061_),
    .B_N(_02137_),
    .Y(_02722_));
 sg13g2_a221oi_1 _07823_ (.B2(_01808_),
    .C1(_02722_),
    .B1(_02721_),
    .A1(_02133_),
    .Y(_02723_),
    .A2(_01764_));
 sg13g2_o21ai_1 _07824_ (.B1(net469),
    .Y(_02724_),
    .A1(_01808_),
    .A2(_02721_));
 sg13g2_and2_1 _07825_ (.A(_02723_),
    .B(_02724_),
    .X(_02725_));
 sg13g2_nor2b_1 _07826_ (.A(\median_processor.input_storage [0]),
    .B_N(net467),
    .Y(_02726_));
 sg13g2_a21oi_1 _07827_ (.A1(net479),
    .A2(_02726_),
    .Y(_02727_),
    .B1(_02055_));
 sg13g2_nor2_1 _07828_ (.A(net479),
    .B(_02726_),
    .Y(_02728_));
 sg13g2_nand2_1 _07829_ (.Y(_02729_),
    .A(_02050_),
    .B(\median_processor.input_storage [26]));
 sg13g2_o21ai_1 _07830_ (.B1(_02729_),
    .Y(_02730_),
    .A1(_02727_),
    .A2(_02728_));
 sg13g2_a22oi_1 _07831_ (.Y(_02731_),
    .B1(\median_processor.input_storage [2]),
    .B2(net416),
    .A2(net465),
    .A1(_01752_));
 sg13g2_a22oi_1 _07832_ (.Y(_02732_),
    .B1(_02730_),
    .B2(_02731_),
    .A2(net466),
    .A1(_01763_));
 sg13g2_nor2_1 _07833_ (.A(_02131_),
    .B(\median_processor.input_storage [7]),
    .Y(_02733_));
 sg13g2_nand2b_1 _07834_ (.Y(_02734_),
    .B(_02061_),
    .A_N(_02137_));
 sg13g2_nand2_1 _07835_ (.Y(_02735_),
    .A(net417),
    .B(_02734_));
 sg13g2_o21ai_1 _07836_ (.B1(_01751_),
    .Y(_02736_),
    .A1(net417),
    .A2(_02734_));
 sg13g2_a22oi_1 _07837_ (.Y(_02737_),
    .B1(_02735_),
    .B2(_02736_),
    .A2(\median_processor.input_storage [7]),
    .A1(_02131_));
 sg13g2_nand4_1 _07838_ (.B(_02059_),
    .C(_02723_),
    .A(_02684_),
    .Y(_02738_),
    .D(_02724_));
 sg13g2_o21ai_1 _07839_ (.B1(_02738_),
    .Y(_02739_),
    .A1(_02733_),
    .A2(_02737_));
 sg13g2_a21o_2 _07840_ (.A2(_02732_),
    .A1(_02725_),
    .B1(_02739_),
    .X(_02740_));
 sg13g2_and2_1 _07841_ (.A(net19),
    .B(_02740_),
    .X(_02741_));
 sg13g2_nor3_1 _07842_ (.A(_01717_),
    .B(_01748_),
    .C(_02690_),
    .Y(_02742_));
 sg13g2_o21ai_1 _07843_ (.B1(_02690_),
    .Y(_02743_),
    .A1(_01717_),
    .A2(_01748_));
 sg13g2_o21ai_1 _07844_ (.B1(_02743_),
    .Y(_02744_),
    .A1(_02431_),
    .A2(_02742_));
 sg13g2_nand3_1 _07845_ (.B(_02741_),
    .C(_02744_),
    .A(net16),
    .Y(_02745_));
 sg13g2_nand4_1 _07846_ (.B(_02741_),
    .C(_02720_),
    .A(_02368_),
    .Y(_02746_),
    .D(_02744_));
 sg13g2_o21ai_1 _07847_ (.B1(_02746_),
    .Y(_02747_),
    .A1(_02720_),
    .A2(_02745_));
 sg13g2_or3_1 _07848_ (.A(_02435_),
    .B(_02627_),
    .C(_02743_),
    .X(_02748_));
 sg13g2_nand3_1 _07849_ (.B(net19),
    .C(_02742_),
    .A(_02435_),
    .Y(_02749_));
 sg13g2_a21oi_1 _07850_ (.A1(_02748_),
    .A2(_02749_),
    .Y(_02750_),
    .B1(_02368_));
 sg13g2_xnor2_1 _07851_ (.Y(_02751_),
    .A(_02435_),
    .B(net19));
 sg13g2_nor3_1 _07852_ (.A(net16),
    .B(_02743_),
    .C(_02751_),
    .Y(_02752_));
 sg13g2_a21oi_1 _07853_ (.A1(_02725_),
    .A2(_02732_),
    .Y(_02753_),
    .B1(_02739_));
 sg13g2_buf_1 _07854_ (.A(_02753_),
    .X(_02754_));
 sg13g2_o21ai_1 _07855_ (.B1(net18),
    .Y(_02755_),
    .A1(_02750_),
    .A2(_02752_));
 sg13g2_inv_1 _07856_ (.Y(_02756_),
    .A(_02719_));
 sg13g2_a22oi_1 _07857_ (.Y(_02757_),
    .B1(_02435_),
    .B2(net19),
    .A2(_02367_),
    .A1(_02346_));
 sg13g2_a21oi_1 _07858_ (.A1(net16),
    .A2(_02751_),
    .Y(_02758_),
    .B1(_02757_));
 sg13g2_nand3_1 _07859_ (.B(_02756_),
    .C(_02758_),
    .A(net18),
    .Y(_02759_));
 sg13g2_nor3_1 _07860_ (.A(_02431_),
    .B(net19),
    .C(_02743_),
    .Y(_02760_));
 sg13g2_nor2_1 _07861_ (.A(_02368_),
    .B(net18),
    .Y(_02761_));
 sg13g2_a21oi_1 _07862_ (.A1(_02760_),
    .A2(_02761_),
    .Y(_02762_),
    .B1(_02166_));
 sg13g2_nand3_1 _07863_ (.B(_02759_),
    .C(_02762_),
    .A(_02755_),
    .Y(_02763_));
 sg13g2_nand3b_1 _07864_ (.B(_02435_),
    .C(_02743_),
    .Y(_02764_),
    .A_N(_02742_));
 sg13g2_nand2b_1 _07865_ (.Y(_02765_),
    .B(_02431_),
    .A_N(_02743_));
 sg13g2_nand2b_1 _07866_ (.Y(_02766_),
    .B(net18),
    .A_N(_02628_));
 sg13g2_a221oi_1 _07867_ (.B2(_02765_),
    .C1(_02766_),
    .B1(_02764_),
    .A1(_02346_),
    .Y(_02767_),
    .A2(_02367_));
 sg13g2_nor2b_1 _07868_ (.A(_02767_),
    .B_N(_02166_),
    .Y(_02768_));
 sg13g2_nand2_1 _07869_ (.Y(_02769_),
    .A(_02628_),
    .B(_02753_));
 sg13g2_or3_1 _07870_ (.A(_02368_),
    .B(_02744_),
    .C(_02769_),
    .X(_02770_));
 sg13g2_or3_1 _07871_ (.A(_02370_),
    .B(_02744_),
    .C(_02769_),
    .X(_02771_));
 sg13g2_mux2_1 _07872_ (.A0(_02770_),
    .A1(_02771_),
    .S(_02720_),
    .X(_02772_));
 sg13g2_nor3_1 _07873_ (.A(_02368_),
    .B(_02744_),
    .C(_02766_),
    .Y(_02773_));
 sg13g2_nand2_1 _07874_ (.Y(_02774_),
    .A(_02720_),
    .B(_02773_));
 sg13g2_nor2_1 _07875_ (.A(_02754_),
    .B(_02719_),
    .Y(_02775_));
 sg13g2_nor4_1 _07876_ (.A(_02370_),
    .B(_02754_),
    .C(_02743_),
    .D(_02751_),
    .Y(_02776_));
 sg13g2_a221oi_1 _07877_ (.B2(_02775_),
    .C1(_02776_),
    .B1(_02758_),
    .A1(_02740_),
    .Y(_02777_),
    .A2(_02750_));
 sg13g2_nand4_1 _07878_ (.B(_02772_),
    .C(_02774_),
    .A(_02768_),
    .Y(_02778_),
    .D(_02777_));
 sg13g2_o21ai_1 _07879_ (.B1(_02778_),
    .Y(_02779_),
    .A1(_02747_),
    .A2(_02763_));
 sg13g2_nor2b_1 _07880_ (.A(net10),
    .B_N(_02779_),
    .Y(_02780_));
 sg13g2_nand2b_2 _07881_ (.Y(_02781_),
    .B(_02780_),
    .A_N(_02648_));
 sg13g2_a221oi_1 _07882_ (.B2(_02548_),
    .C1(_02781_),
    .B1(net2),
    .A1(_02267_),
    .Y(_02782_),
    .A2(_02268_));
 sg13g2_a21o_1 _07883_ (.A2(_01949_),
    .A1(net393),
    .B1(_01944_),
    .X(_02783_));
 sg13g2_o21ai_1 _07884_ (.B1(_02783_),
    .Y(_02784_),
    .A1(net393),
    .A2(_01949_));
 sg13g2_nor2_1 _07885_ (.A(net15),
    .B(_02740_),
    .Y(_02785_));
 sg13g2_a21oi_1 _07886_ (.A1(net15),
    .A2(_02740_),
    .Y(_02786_),
    .B1(_02511_));
 sg13g2_nor3_1 _07887_ (.A(_02784_),
    .B(_02785_),
    .C(_02786_),
    .Y(_02787_));
 sg13g2_o21ai_1 _07888_ (.B1(_02784_),
    .Y(_02788_),
    .A1(_02785_),
    .A2(_02786_));
 sg13g2_nor2_1 _07889_ (.A(_02572_),
    .B(_02788_),
    .Y(_02789_));
 sg13g2_a21oi_1 _07890_ (.A1(_02572_),
    .A2(_02787_),
    .Y(_02790_),
    .B1(_02789_));
 sg13g2_xor2_1 _07891_ (.B(net15),
    .A(_02511_),
    .X(_02791_));
 sg13g2_xnor2_1 _07892_ (.Y(_02792_),
    .A(net18),
    .B(_02791_));
 sg13g2_nand2b_1 _07893_ (.Y(_02793_),
    .B(_02792_),
    .A_N(_02243_));
 sg13g2_xor2_1 _07894_ (.B(_02792_),
    .A(_02243_),
    .X(_02794_));
 sg13g2_mux2_1 _07895_ (.A0(_02793_),
    .A1(_02794_),
    .S(net17),
    .X(_02795_));
 sg13g2_o21ai_1 _07896_ (.B1(_02265_),
    .Y(_02796_),
    .A1(_02790_),
    .A2(_02795_));
 sg13g2_and2_1 _07897_ (.A(_02511_),
    .B(net15),
    .X(_02797_));
 sg13g2_mux2_1 _07898_ (.A0(_02797_),
    .A1(_02791_),
    .S(net17),
    .X(_02798_));
 sg13g2_xnor2_1 _07899_ (.Y(_02799_),
    .A(_02243_),
    .B(_02740_));
 sg13g2_nor2_1 _07900_ (.A(_02511_),
    .B(net15),
    .Y(_02800_));
 sg13g2_mux2_1 _07901_ (.A0(_02791_),
    .A1(_02800_),
    .S(net17),
    .X(_02801_));
 sg13g2_nor2_1 _07902_ (.A(_02243_),
    .B(net18),
    .Y(_02802_));
 sg13g2_and4_1 _07903_ (.A(_02243_),
    .B(net17),
    .C(net18),
    .D(_02797_),
    .X(_02803_));
 sg13g2_a221oi_1 _07904_ (.B2(_02802_),
    .C1(_02803_),
    .B1(_02801_),
    .A1(_02798_),
    .Y(_02804_),
    .A2(_02799_));
 sg13g2_nor3_1 _07905_ (.A(_02572_),
    .B(_02784_),
    .C(_02804_),
    .Y(_02805_));
 sg13g2_nand2_1 _07906_ (.Y(_02806_),
    .A(net18),
    .B(_02797_));
 sg13g2_nand2_1 _07907_ (.Y(_02807_),
    .A(_02740_),
    .B(_02791_));
 sg13g2_nand2b_1 _07908_ (.Y(_02808_),
    .B(_02243_),
    .A_N(net17));
 sg13g2_a21oi_1 _07909_ (.A1(_02806_),
    .A2(_02807_),
    .Y(_02809_),
    .B1(_02808_));
 sg13g2_o21ai_1 _07910_ (.B1(_02784_),
    .Y(_02810_),
    .A1(_02572_),
    .A2(_02809_));
 sg13g2_a21oi_1 _07911_ (.A1(_02572_),
    .A2(_02804_),
    .Y(_02811_),
    .B1(_02810_));
 sg13g2_or2_1 _07912_ (.X(_02812_),
    .B(_02811_),
    .A(_02805_));
 sg13g2_nand3b_1 _07913_ (.B(_02780_),
    .C(net7),
    .Y(_02813_),
    .A_N(_02648_));
 sg13g2_nor4_2 _07914_ (.A(net4),
    .B(_02796_),
    .C(_02812_),
    .Y(_02814_),
    .D(_02813_));
 sg13g2_buf_1 _07915_ (.A(_02814_),
    .X(_02815_));
 sg13g2_nor2_1 _07916_ (.A(_02782_),
    .B(net1),
    .Y(_02816_));
 sg13g2_nor2_2 _07917_ (.A(net10),
    .B(_02779_),
    .Y(_02817_));
 sg13g2_a221oi_1 _07918_ (.B2(_02159_),
    .C1(net4),
    .B1(_02817_),
    .A1(_01907_),
    .Y(_02818_),
    .A2(net10));
 sg13g2_a21o_1 _07919_ (.A2(_02548_),
    .A1(net4),
    .B1(_02818_),
    .X(_02819_));
 sg13g2_buf_1 _07920_ (.A(_02648_),
    .X(_02820_));
 sg13g2_mux2_1 _07921_ (.A0(_02819_),
    .A1(net457),
    .S(net6),
    .X(_02821_));
 sg13g2_and2_1 _07922_ (.A(\median_processor.median_processor.median_out [0]),
    .B(net1),
    .X(_02822_));
 sg13g2_a21o_1 _07923_ (.A2(_02821_),
    .A1(_02816_),
    .B1(_02822_),
    .X(_00064_));
 sg13g2_a221oi_1 _07924_ (.B2(_01727_),
    .C1(net2),
    .B1(_02817_),
    .A1(_01908_),
    .Y(_02823_),
    .A2(net10));
 sg13g2_nor2_1 _07925_ (.A(net6),
    .B(_02823_),
    .Y(_02824_));
 sg13g2_buf_1 _07926_ (.A(_02265_),
    .X(_02825_));
 sg13g2_nor2_1 _07927_ (.A(net428),
    .B(net9),
    .Y(_02826_));
 sg13g2_a21oi_1 _07928_ (.A1(_02055_),
    .A2(net9),
    .Y(_02827_),
    .B1(_02826_));
 sg13g2_nor2_1 _07929_ (.A(_02813_),
    .B(_02827_),
    .Y(_02828_));
 sg13g2_buf_1 _07930_ (.A(_02536_),
    .X(_02829_));
 sg13g2_nand2_1 _07931_ (.Y(_02830_),
    .A(net474),
    .B(net5));
 sg13g2_o21ai_1 _07932_ (.B1(_02830_),
    .Y(_02831_),
    .A1(_02022_),
    .A2(net5));
 sg13g2_nand2_1 _07933_ (.Y(_02832_),
    .A(net2),
    .B(_02831_));
 sg13g2_o21ai_1 _07934_ (.B1(_02832_),
    .Y(_02833_),
    .A1(_02824_),
    .A2(_02828_));
 sg13g2_nor3_1 _07935_ (.A(net468),
    .B(net7),
    .C(_02781_),
    .Y(_02834_));
 sg13g2_a221oi_1 _07936_ (.B2(_02834_),
    .C1(net1),
    .B1(_02832_),
    .A1(net458),
    .Y(_02835_),
    .A2(net6));
 sg13g2_and2_1 _07937_ (.A(\median_processor.median_processor.median_out [1]),
    .B(net1),
    .X(_02836_));
 sg13g2_a21o_1 _07938_ (.A2(_02835_),
    .A1(_02833_),
    .B1(_02836_),
    .X(_00065_));
 sg13g2_a221oi_1 _07939_ (.B2(net416),
    .C1(net2),
    .B1(_02817_),
    .A1(_02326_),
    .Y(_02837_),
    .A2(net10));
 sg13g2_nor2_1 _07940_ (.A(net6),
    .B(_02837_),
    .Y(_02838_));
 sg13g2_nor2_1 _07941_ (.A(net424),
    .B(net9),
    .Y(_02839_));
 sg13g2_a21oi_1 _07942_ (.A1(net425),
    .A2(net9),
    .Y(_02840_),
    .B1(_02839_));
 sg13g2_nor2_1 _07943_ (.A(_02813_),
    .B(_02840_),
    .Y(_02841_));
 sg13g2_nand2_1 _07944_ (.Y(_02842_),
    .A(net420),
    .B(_02536_));
 sg13g2_o21ai_1 _07945_ (.B1(_02842_),
    .Y(_02843_),
    .A1(_01979_),
    .A2(net5));
 sg13g2_nand2_1 _07946_ (.Y(_02844_),
    .A(net2),
    .B(_02843_));
 sg13g2_o21ai_1 _07947_ (.B1(_02844_),
    .Y(_02845_),
    .A1(_02838_),
    .A2(_02841_));
 sg13g2_nor3_1 _07948_ (.A(net459),
    .B(net7),
    .C(_02781_),
    .Y(_02846_));
 sg13g2_a221oi_1 _07949_ (.B2(_02846_),
    .C1(net1),
    .B1(_02844_),
    .A1(_01814_),
    .Y(_02847_),
    .A2(net6));
 sg13g2_and2_1 _07950_ (.A(\median_processor.median_processor.median_out [2]),
    .B(_02814_),
    .X(_02848_));
 sg13g2_a21o_1 _07951_ (.A2(_02847_),
    .A1(_02845_),
    .B1(_02848_),
    .X(_00066_));
 sg13g2_a221oi_1 _07952_ (.B2(net465),
    .C1(net4),
    .B1(_02817_),
    .A1(_02189_),
    .Y(_02849_),
    .A2(net10));
 sg13g2_nor2_1 _07953_ (.A(net6),
    .B(_02849_),
    .Y(_02850_));
 sg13g2_nor2_1 _07954_ (.A(net430),
    .B(net9),
    .Y(_02851_));
 sg13g2_a21oi_1 _07955_ (.A1(_01763_),
    .A2(net9),
    .Y(_02852_),
    .B1(_02851_));
 sg13g2_nor2_1 _07956_ (.A(_02813_),
    .B(_02852_),
    .Y(_02853_));
 sg13g2_nand2_1 _07957_ (.Y(_02854_),
    .A(net451),
    .B(_02536_));
 sg13g2_o21ai_1 _07958_ (.B1(_02854_),
    .Y(_02855_),
    .A1(_01977_),
    .A2(net5));
 sg13g2_nand2_1 _07959_ (.Y(_02856_),
    .A(net2),
    .B(_02855_));
 sg13g2_o21ai_1 _07960_ (.B1(_02856_),
    .Y(_02857_),
    .A1(_02850_),
    .A2(_02853_));
 sg13g2_nor3_1 _07961_ (.A(net464),
    .B(net7),
    .C(_02781_),
    .Y(_02858_));
 sg13g2_a221oi_1 _07962_ (.B2(_02858_),
    .C1(net1),
    .B1(_02856_),
    .A1(_02210_),
    .Y(_02859_),
    .A2(net6));
 sg13g2_and2_1 _07963_ (.A(\median_processor.median_processor.median_out [3]),
    .B(_02814_),
    .X(_02860_));
 sg13g2_a21o_1 _07964_ (.A2(_02859_),
    .A1(_02857_),
    .B1(_02860_),
    .X(_00067_));
 sg13g2_a221oi_1 _07965_ (.B2(_02684_),
    .C1(net4),
    .B1(_02817_),
    .A1(_02655_),
    .Y(_02861_),
    .A2(net10));
 sg13g2_nor2_1 _07966_ (.A(net6),
    .B(_02861_),
    .Y(_02862_));
 sg13g2_nor2_1 _07967_ (.A(net431),
    .B(_02265_),
    .Y(_02863_));
 sg13g2_a21oi_1 _07968_ (.A1(_01764_),
    .A2(net9),
    .Y(_02864_),
    .B1(_02863_));
 sg13g2_nor2_1 _07969_ (.A(_02813_),
    .B(_02864_),
    .Y(_02865_));
 sg13g2_nand2_1 _07970_ (.Y(_02866_),
    .A(net450),
    .B(_02536_));
 sg13g2_o21ai_1 _07971_ (.B1(_02866_),
    .Y(_02867_),
    .A1(net390),
    .A2(net5));
 sg13g2_nand2_1 _07972_ (.Y(_02868_),
    .A(net2),
    .B(_02867_));
 sg13g2_o21ai_1 _07973_ (.B1(_02868_),
    .Y(_02869_),
    .A1(_02862_),
    .A2(_02865_));
 sg13g2_nor3_1 _07974_ (.A(net456),
    .B(net7),
    .C(_02781_),
    .Y(_02870_));
 sg13g2_a221oi_1 _07975_ (.B2(_02870_),
    .C1(net1),
    .B1(_02868_),
    .A1(net387),
    .Y(_02871_),
    .A2(_02820_));
 sg13g2_and2_1 _07976_ (.A(\median_processor.median_processor.median_out [4]),
    .B(_02814_),
    .X(_02872_));
 sg13g2_a21o_1 _07977_ (.A2(_02871_),
    .A1(_02869_),
    .B1(_02872_),
    .X(_00068_));
 sg13g2_a221oi_1 _07978_ (.B2(_02687_),
    .C1(net4),
    .B1(_02817_),
    .A1(net443),
    .Y(_02873_),
    .A2(net10));
 sg13g2_nor2_1 _07979_ (.A(_02648_),
    .B(_02873_),
    .Y(_02874_));
 sg13g2_nor2_1 _07980_ (.A(net427),
    .B(_02265_),
    .Y(_02875_));
 sg13g2_a21oi_1 _07981_ (.A1(_01762_),
    .A2(net9),
    .Y(_02876_),
    .B1(_02875_));
 sg13g2_nor2_1 _07982_ (.A(_02813_),
    .B(_02876_),
    .Y(_02877_));
 sg13g2_nand2_1 _07983_ (.Y(_02878_),
    .A(net449),
    .B(_02536_));
 sg13g2_o21ai_1 _07984_ (.B1(_02878_),
    .Y(_02879_),
    .A1(net389),
    .A2(net5));
 sg13g2_nand2_1 _07985_ (.Y(_02880_),
    .A(net2),
    .B(_02879_));
 sg13g2_o21ai_1 _07986_ (.B1(_02880_),
    .Y(_02881_),
    .A1(_02874_),
    .A2(_02877_));
 sg13g2_nor3_1 _07987_ (.A(net471),
    .B(net7),
    .C(_02781_),
    .Y(_02882_));
 sg13g2_a221oi_1 _07988_ (.B2(_02882_),
    .C1(net1),
    .B1(_02880_),
    .A1(net395),
    .Y(_02883_),
    .A2(_02820_));
 sg13g2_and2_1 _07989_ (.A(\median_processor.median_processor.median_out [5]),
    .B(_02814_),
    .X(_02884_));
 sg13g2_a21o_1 _07990_ (.A2(_02883_),
    .A1(_02881_),
    .B1(_02884_),
    .X(_00069_));
 sg13g2_nand2_1 _07991_ (.Y(_02885_),
    .A(net447),
    .B(net5));
 sg13g2_o21ai_1 _07992_ (.B1(_02885_),
    .Y(_02886_),
    .A1(_01965_),
    .A2(net5));
 sg13g2_a221oi_1 _07993_ (.B2(_01710_),
    .C1(net4),
    .B1(_02817_),
    .A1(net392),
    .Y(_02887_),
    .A2(_02718_));
 sg13g2_or2_1 _07994_ (.X(_02888_),
    .B(_02887_),
    .A(_02648_));
 sg13g2_nor2_1 _07995_ (.A(net421),
    .B(_02265_),
    .Y(_02889_));
 sg13g2_a21oi_1 _07996_ (.A1(net462),
    .A2(_02825_),
    .Y(_02890_),
    .B1(_02889_));
 sg13g2_or2_1 _07997_ (.X(_02891_),
    .B(_02890_),
    .A(_02813_));
 sg13g2_a22oi_1 _07998_ (.Y(_02892_),
    .B1(_02888_),
    .B2(_02891_),
    .A2(_02886_),
    .A1(_02546_));
 sg13g2_nor2b_1 _07999_ (.A(net388),
    .B_N(_02648_),
    .Y(_02893_));
 sg13g2_nor3_1 _08000_ (.A(net470),
    .B(_02016_),
    .C(_02781_),
    .Y(_02894_));
 sg13g2_or3_1 _08001_ (.A(_02814_),
    .B(_02893_),
    .C(_02894_),
    .X(_02895_));
 sg13g2_nand2_1 _08002_ (.Y(_02896_),
    .A(\median_processor.median_processor.median_out [6]),
    .B(_02815_));
 sg13g2_o21ai_1 _08003_ (.B1(_02896_),
    .Y(_00070_),
    .A1(_02892_),
    .A2(_02895_));
 sg13g2_nand2_1 _08004_ (.Y(_02897_),
    .A(net413),
    .B(_02829_));
 sg13g2_o21ai_1 _08005_ (.B1(_02897_),
    .Y(_02898_),
    .A1(_01962_),
    .A2(_02829_));
 sg13g2_a221oi_1 _08006_ (.B2(_02131_),
    .C1(_02545_),
    .B1(_02817_),
    .A1(net222),
    .Y(_02899_),
    .A2(_02718_));
 sg13g2_or2_1 _08007_ (.X(_02900_),
    .B(_02899_),
    .A(_02648_));
 sg13g2_nor2_1 _08008_ (.A(net426),
    .B(_02265_),
    .Y(_02901_));
 sg13g2_a21oi_1 _08009_ (.A1(net391),
    .A2(_02825_),
    .Y(_02902_),
    .B1(_02901_));
 sg13g2_or2_1 _08010_ (.X(_02903_),
    .B(_02902_),
    .A(_02813_));
 sg13g2_a22oi_1 _08011_ (.Y(_02904_),
    .B1(_02900_),
    .B2(_02903_),
    .A2(_02898_),
    .A1(_02546_));
 sg13g2_and2_1 _08012_ (.A(_01847_),
    .B(_02648_),
    .X(_02905_));
 sg13g2_nor3_1 _08013_ (.A(net393),
    .B(_02016_),
    .C(_02781_),
    .Y(_02906_));
 sg13g2_or3_1 _08014_ (.A(_02814_),
    .B(_02905_),
    .C(_02906_),
    .X(_02907_));
 sg13g2_nand2_1 _08015_ (.Y(_02908_),
    .A(\median_processor.median_processor.median_out [7]),
    .B(_02815_));
 sg13g2_o21ai_1 _08016_ (.B1(_02908_),
    .Y(_00071_),
    .A1(_02904_),
    .A2(_02907_));
 sg13g2_buf_1 _08017_ (.A(\median_processor.rst ),
    .X(_02909_));
 sg13g2_buf_1 _08018_ (.A(net494),
    .X(_02910_));
 sg13g2_buf_1 _08019_ (.A(net412),
    .X(_02911_));
 sg13g2_buf_1 _08020_ (.A(data_in_p2c_1),
    .X(_02912_));
 sg13g2_nand2b_2 _08021_ (.Y(_02913_),
    .B(\median_processor.wr_enable ),
    .A_N(reg_addr_p2c_1));
 sg13g2_nor2_1 _08022_ (.A(reg_addr_p2c_3),
    .B(reg_addr_p2c_2),
    .Y(_02914_));
 sg13g2_nand2b_1 _08023_ (.Y(_02915_),
    .B(_02914_),
    .A_N(_02913_));
 sg13g2_buf_1 _08024_ (.A(_02915_),
    .X(_02916_));
 sg13g2_mux2_1 _08025_ (.A0(net493),
    .A1(net484),
    .S(net385),
    .X(_02917_));
 sg13g2_and2_1 _08026_ (.A(net386),
    .B(_02917_),
    .X(_00000_));
 sg13g2_nand3_1 _08027_ (.B(\median_processor.wr_enable ),
    .C(_02914_),
    .A(reg_addr_p2c_1),
    .Y(_02918_));
 sg13g2_buf_1 _08028_ (.A(_02918_),
    .X(_02919_));
 sg13g2_inv_2 _08029_ (.Y(_02920_),
    .A(data_in_p2c_3));
 sg13g2_nor2_1 _08030_ (.A(_02920_),
    .B(net384),
    .Y(_02921_));
 sg13g2_a21oi_1 _08031_ (.A1(net424),
    .A2(net384),
    .Y(_02922_),
    .B1(_02921_));
 sg13g2_nor2b_1 _08032_ (.A(_02922_),
    .B_N(net386),
    .Y(_00001_));
 sg13g2_buf_1 _08033_ (.A(data_in_p2c_4),
    .X(_02923_));
 sg13g2_mux2_1 _08034_ (.A0(net492),
    .A1(net430),
    .S(net384),
    .X(_02924_));
 sg13g2_and2_1 _08035_ (.A(net386),
    .B(_02924_),
    .X(_00002_));
 sg13g2_buf_1 _08036_ (.A(data_in_p2c_5),
    .X(_02925_));
 sg13g2_mux2_1 _08037_ (.A0(net491),
    .A1(net431),
    .S(net384),
    .X(_02926_));
 sg13g2_and2_1 _08038_ (.A(net386),
    .B(_02926_),
    .X(_00003_));
 sg13g2_buf_1 _08039_ (.A(data_in_p2c_6),
    .X(_02927_));
 sg13g2_mux2_1 _08040_ (.A0(net490),
    .A1(net427),
    .S(net384),
    .X(_02928_));
 sg13g2_and2_1 _08041_ (.A(net386),
    .B(_02928_),
    .X(_00004_));
 sg13g2_inv_1 _08042_ (.Y(_02929_),
    .A(net495));
 sg13g2_nor2_1 _08043_ (.A(_02929_),
    .B(net384),
    .Y(_02930_));
 sg13g2_a21oi_1 _08044_ (.A1(net421),
    .A2(_02919_),
    .Y(_02931_),
    .B1(_02930_));
 sg13g2_nor2b_1 _08045_ (.A(_02931_),
    .B_N(_02911_),
    .Y(_00005_));
 sg13g2_buf_1 _08046_ (.A(data_in_p2c_8),
    .X(_02932_));
 sg13g2_mux2_1 _08047_ (.A0(net489),
    .A1(net426),
    .S(_02919_),
    .X(_02933_));
 sg13g2_and2_1 _08048_ (.A(_02911_),
    .B(_02933_),
    .X(_00006_));
 sg13g2_nand2b_1 _08049_ (.Y(_02934_),
    .B(reg_addr_p2c_2),
    .A_N(reg_addr_p2c_3));
 sg13g2_nor2_2 _08050_ (.A(_02913_),
    .B(_02934_),
    .Y(_02935_));
 sg13g2_buf_1 _08051_ (.A(_02935_),
    .X(_02936_));
 sg13g2_nand2_1 _08052_ (.Y(_02937_),
    .A(net493),
    .B(net383));
 sg13g2_o21ai_1 _08053_ (.B1(_02937_),
    .Y(_02938_),
    .A1(_01980_),
    .A2(net383));
 sg13g2_and2_1 _08054_ (.A(net386),
    .B(_02938_),
    .X(_00007_));
 sg13g2_buf_1 _08055_ (.A(data_in_p2c_2),
    .X(_02939_));
 sg13g2_nand2_1 _08056_ (.Y(_02940_),
    .A(net488),
    .B(net383));
 sg13g2_o21ai_1 _08057_ (.B1(_02940_),
    .Y(_02941_),
    .A1(_01755_),
    .A2(net383));
 sg13g2_and2_1 _08058_ (.A(net386),
    .B(_02941_),
    .X(_00008_));
 sg13g2_mux2_1 _08059_ (.A0(_01815_),
    .A1(data_in_p2c_3),
    .S(_02935_),
    .X(_02942_));
 sg13g2_and2_1 _08060_ (.A(net386),
    .B(_02942_),
    .X(_00009_));
 sg13g2_buf_1 _08061_ (.A(net412),
    .X(_02943_));
 sg13g2_nand2_1 _08062_ (.Y(_02944_),
    .A(net492),
    .B(net383));
 sg13g2_o21ai_1 _08063_ (.B1(_02944_),
    .Y(_02945_),
    .A1(net396),
    .A2(net383));
 sg13g2_and2_1 _08064_ (.A(net382),
    .B(_02945_),
    .X(_00010_));
 sg13g2_mux2_1 _08065_ (.A0(net488),
    .A1(\median_processor.input_storage [1]),
    .S(net385),
    .X(_02946_));
 sg13g2_and2_1 _08066_ (.A(net382),
    .B(_02946_),
    .X(_00011_));
 sg13g2_nand2_1 _08067_ (.Y(_02947_),
    .A(net491),
    .B(_02935_));
 sg13g2_o21ai_1 _08068_ (.B1(_02947_),
    .Y(_02948_),
    .A1(_01872_),
    .A2(net383));
 sg13g2_and2_1 _08069_ (.A(net382),
    .B(_02948_),
    .X(_00012_));
 sg13g2_nand2_1 _08070_ (.Y(_02949_),
    .A(net490),
    .B(_02935_));
 sg13g2_o21ai_1 _08071_ (.B1(_02949_),
    .Y(_02950_),
    .A1(_01772_),
    .A2(net383));
 sg13g2_and2_1 _08072_ (.A(net382),
    .B(_02950_),
    .X(_00013_));
 sg13g2_nand2_1 _08073_ (.Y(_02951_),
    .A(net495),
    .B(_02935_));
 sg13g2_o21ai_1 _08074_ (.B1(_02951_),
    .Y(_02952_),
    .A1(_01799_),
    .A2(_02936_));
 sg13g2_and2_1 _08075_ (.A(_02943_),
    .B(_02952_),
    .X(_00014_));
 sg13g2_nand2_1 _08076_ (.Y(_02953_),
    .A(net489),
    .B(_02935_));
 sg13g2_o21ai_1 _08077_ (.B1(_02953_),
    .Y(_02954_),
    .A1(_01714_),
    .A2(_02936_));
 sg13g2_and2_1 _08078_ (.A(_02943_),
    .B(_02954_),
    .X(_00015_));
 sg13g2_nand2_2 _08079_ (.Y(_02955_),
    .A(reg_addr_p2c_1),
    .B(\median_processor.wr_enable ));
 sg13g2_nor2_2 _08080_ (.A(_02955_),
    .B(_02934_),
    .Y(_02956_));
 sg13g2_buf_1 _08081_ (.A(_02956_),
    .X(_02957_));
 sg13g2_nand2_1 _08082_ (.Y(_02958_),
    .A(net493),
    .B(net381));
 sg13g2_o21ai_1 _08083_ (.B1(_02958_),
    .Y(_02959_),
    .A1(_02159_),
    .A2(net381));
 sg13g2_and2_1 _08084_ (.A(net382),
    .B(_02959_),
    .X(_00016_));
 sg13g2_nand2_1 _08085_ (.Y(_02960_),
    .A(net488),
    .B(net381));
 sg13g2_o21ai_1 _08086_ (.B1(_02960_),
    .Y(_02961_),
    .A1(_01727_),
    .A2(net381));
 sg13g2_and2_1 _08087_ (.A(net382),
    .B(_02961_),
    .X(_00017_));
 sg13g2_nand2_1 _08088_ (.Y(_02962_),
    .A(data_in_p2c_3),
    .B(_02956_));
 sg13g2_o21ai_1 _08089_ (.B1(_02962_),
    .Y(_02963_),
    .A1(_02150_),
    .A2(net381));
 sg13g2_and2_1 _08090_ (.A(net382),
    .B(_02963_),
    .X(_00018_));
 sg13g2_nand2_1 _08091_ (.Y(_02964_),
    .A(net492),
    .B(_02956_));
 sg13g2_o21ai_1 _08092_ (.B1(_02964_),
    .Y(_02965_),
    .A1(_01731_),
    .A2(net381));
 sg13g2_and2_1 _08093_ (.A(net382),
    .B(_02965_),
    .X(_00019_));
 sg13g2_buf_1 _08094_ (.A(net412),
    .X(_02966_));
 sg13g2_nand2_1 _08095_ (.Y(_02967_),
    .A(net491),
    .B(_02956_));
 sg13g2_o21ai_1 _08096_ (.B1(_02967_),
    .Y(_02968_),
    .A1(_02684_),
    .A2(net381));
 sg13g2_and2_1 _08097_ (.A(net380),
    .B(_02968_),
    .X(_00020_));
 sg13g2_nand2_1 _08098_ (.Y(_02969_),
    .A(net490),
    .B(_02956_));
 sg13g2_o21ai_1 _08099_ (.B1(_02969_),
    .Y(_02970_),
    .A1(_02687_),
    .A2(net381));
 sg13g2_and2_1 _08100_ (.A(net380),
    .B(_02970_),
    .X(_00021_));
 sg13g2_nand2_1 _08101_ (.Y(_02971_),
    .A(net478),
    .B(net385));
 sg13g2_o21ai_1 _08102_ (.B1(_02971_),
    .Y(_02972_),
    .A1(_02920_),
    .A2(net385));
 sg13g2_and2_1 _08103_ (.A(_02966_),
    .B(_02972_),
    .X(_00022_));
 sg13g2_nand2_1 _08104_ (.Y(_02973_),
    .A(net495),
    .B(_02956_));
 sg13g2_o21ai_1 _08105_ (.B1(_02973_),
    .Y(_02974_),
    .A1(_01710_),
    .A2(_02957_));
 sg13g2_and2_1 _08106_ (.A(net380),
    .B(_02974_),
    .X(_00023_));
 sg13g2_nand2_1 _08107_ (.Y(_02975_),
    .A(net489),
    .B(_02956_));
 sg13g2_o21ai_1 _08108_ (.B1(_02975_),
    .Y(_02976_),
    .A1(_02131_),
    .A2(_02957_));
 sg13g2_and2_1 _08109_ (.A(net380),
    .B(_02976_),
    .X(_00024_));
 sg13g2_nand2b_1 _08110_ (.Y(_02977_),
    .B(reg_addr_p2c_3),
    .A_N(reg_addr_p2c_2));
 sg13g2_nor2_2 _08111_ (.A(_02913_),
    .B(_02977_),
    .Y(_02978_));
 sg13g2_buf_1 _08112_ (.A(_02978_),
    .X(_02979_));
 sg13g2_nand2_1 _08113_ (.Y(_02980_),
    .A(net493),
    .B(net379));
 sg13g2_o21ai_1 _08114_ (.B1(_02980_),
    .Y(_02981_),
    .A1(_01907_),
    .A2(net379));
 sg13g2_and2_1 _08115_ (.A(net380),
    .B(_02981_),
    .X(_00025_));
 sg13g2_nand2_1 _08116_ (.Y(_02982_),
    .A(net488),
    .B(net379));
 sg13g2_o21ai_1 _08117_ (.B1(_02982_),
    .Y(_02983_),
    .A1(_01908_),
    .A2(net379));
 sg13g2_and2_1 _08118_ (.A(net380),
    .B(_02983_),
    .X(_00026_));
 sg13g2_nand2_1 _08119_ (.Y(_02984_),
    .A(data_in_p2c_3),
    .B(_02978_));
 sg13g2_o21ai_1 _08120_ (.B1(_02984_),
    .Y(_02985_),
    .A1(_02326_),
    .A2(net379));
 sg13g2_and2_1 _08121_ (.A(net380),
    .B(_02985_),
    .X(_00027_));
 sg13g2_nand2_1 _08122_ (.Y(_02986_),
    .A(net492),
    .B(_02978_));
 sg13g2_o21ai_1 _08123_ (.B1(_02986_),
    .Y(_02987_),
    .A1(_02189_),
    .A2(net379));
 sg13g2_and2_1 _08124_ (.A(net380),
    .B(_02987_),
    .X(_00028_));
 sg13g2_nand2_1 _08125_ (.Y(_02988_),
    .A(net491),
    .B(_02978_));
 sg13g2_o21ai_1 _08126_ (.B1(_02988_),
    .Y(_02989_),
    .A1(_02655_),
    .A2(net379));
 sg13g2_and2_1 _08127_ (.A(_02966_),
    .B(_02989_),
    .X(_00029_));
 sg13g2_buf_1 _08128_ (.A(net412),
    .X(_02990_));
 sg13g2_nand2_1 _08129_ (.Y(_02991_),
    .A(net490),
    .B(_02978_));
 sg13g2_o21ai_1 _08130_ (.B1(_02991_),
    .Y(_02992_),
    .A1(_01904_),
    .A2(net379));
 sg13g2_and2_1 _08131_ (.A(net378),
    .B(_02992_),
    .X(_00030_));
 sg13g2_nand2_1 _08132_ (.Y(_02993_),
    .A(net495),
    .B(_02978_));
 sg13g2_o21ai_1 _08133_ (.B1(_02993_),
    .Y(_02994_),
    .A1(_01929_),
    .A2(_02979_));
 sg13g2_and2_1 _08134_ (.A(net378),
    .B(_02994_),
    .X(_00031_));
 sg13g2_nand2_1 _08135_ (.Y(_02995_),
    .A(net489),
    .B(_02978_));
 sg13g2_o21ai_1 _08136_ (.B1(_02995_),
    .Y(_02996_),
    .A1(_01902_),
    .A2(_02979_));
 sg13g2_and2_1 _08137_ (.A(net378),
    .B(_02996_),
    .X(_00032_));
 sg13g2_mux2_1 _08138_ (.A0(net492),
    .A1(_01752_),
    .S(net385),
    .X(_02997_));
 sg13g2_and2_1 _08139_ (.A(net378),
    .B(_02997_),
    .X(_00033_));
 sg13g2_nor2_2 _08140_ (.A(_02955_),
    .B(_02977_),
    .Y(_02998_));
 sg13g2_mux2_1 _08141_ (.A0(_01981_),
    .A1(_02912_),
    .S(_02998_),
    .X(_02999_));
 sg13g2_and2_1 _08142_ (.A(net378),
    .B(_02999_),
    .X(_00034_));
 sg13g2_buf_1 _08143_ (.A(_02998_),
    .X(_03000_));
 sg13g2_nand2_1 _08144_ (.Y(_03001_),
    .A(_02939_),
    .B(net377));
 sg13g2_o21ai_1 _08145_ (.B1(_03001_),
    .Y(_03002_),
    .A1(_02022_),
    .A2(net377));
 sg13g2_and2_1 _08146_ (.A(net378),
    .B(_03002_),
    .X(_00035_));
 sg13g2_nand2_1 _08147_ (.Y(_03003_),
    .A(data_in_p2c_3),
    .B(net377));
 sg13g2_o21ai_1 _08148_ (.B1(_03003_),
    .Y(_03004_),
    .A1(_01979_),
    .A2(net377));
 sg13g2_and2_1 _08149_ (.A(net378),
    .B(_03004_),
    .X(_00036_));
 sg13g2_nand2_1 _08150_ (.Y(_03005_),
    .A(_02923_),
    .B(net377));
 sg13g2_o21ai_1 _08151_ (.B1(_03005_),
    .Y(_03006_),
    .A1(_01977_),
    .A2(net377));
 sg13g2_and2_1 _08152_ (.A(net378),
    .B(_03006_),
    .X(_00037_));
 sg13g2_nand2_1 _08153_ (.Y(_03007_),
    .A(net491),
    .B(_02998_));
 sg13g2_o21ai_1 _08154_ (.B1(_03007_),
    .Y(_03008_),
    .A1(net390),
    .A2(net377));
 sg13g2_and2_1 _08155_ (.A(_02990_),
    .B(_03008_),
    .X(_00038_));
 sg13g2_nand2_1 _08156_ (.Y(_03009_),
    .A(_02927_),
    .B(_02998_));
 sg13g2_o21ai_1 _08157_ (.B1(_03009_),
    .Y(_03010_),
    .A1(net389),
    .A2(net377));
 sg13g2_and2_1 _08158_ (.A(_02990_),
    .B(_03010_),
    .X(_00039_));
 sg13g2_buf_1 _08159_ (.A(_02910_),
    .X(_03011_));
 sg13g2_nand2_1 _08160_ (.Y(_03012_),
    .A(data_in_p2c_7),
    .B(_02998_));
 sg13g2_o21ai_1 _08161_ (.B1(_03012_),
    .Y(_03013_),
    .A1(_01965_),
    .A2(_03000_));
 sg13g2_and2_1 _08162_ (.A(net376),
    .B(_03013_),
    .X(_00040_));
 sg13g2_nand2_1 _08163_ (.Y(_03014_),
    .A(_02932_),
    .B(_02998_));
 sg13g2_o21ai_1 _08164_ (.B1(_03014_),
    .Y(_03015_),
    .A1(net439),
    .A2(_03000_));
 sg13g2_and2_1 _08165_ (.A(net376),
    .B(_03015_),
    .X(_00041_));
 sg13g2_nand2_1 _08166_ (.Y(_03016_),
    .A(reg_addr_p2c_3),
    .B(reg_addr_p2c_2));
 sg13g2_nor2_2 _08167_ (.A(_02913_),
    .B(_03016_),
    .Y(_03017_));
 sg13g2_buf_1 _08168_ (.A(_03017_),
    .X(_03018_));
 sg13g2_nand2_1 _08169_ (.Y(_03019_),
    .A(_02912_),
    .B(net375));
 sg13g2_o21ai_1 _08170_ (.B1(_03019_),
    .Y(_03020_),
    .A1(_01876_),
    .A2(net375));
 sg13g2_and2_1 _08171_ (.A(net376),
    .B(_03020_),
    .X(_00042_));
 sg13g2_nand2_1 _08172_ (.Y(_03021_),
    .A(_02939_),
    .B(net375));
 sg13g2_o21ai_1 _08173_ (.B1(_03021_),
    .Y(_03022_),
    .A1(_01882_),
    .A2(net375));
 sg13g2_and2_1 _08174_ (.A(net376),
    .B(_03022_),
    .X(_00043_));
 sg13g2_mux2_1 _08175_ (.A0(_02925_),
    .A1(net423),
    .S(net385),
    .X(_03023_));
 sg13g2_and2_1 _08176_ (.A(net376),
    .B(_03023_),
    .X(_00044_));
 sg13g2_nand2_1 _08177_ (.Y(_03024_),
    .A(data_in_p2c_3),
    .B(_03017_));
 sg13g2_o21ai_1 _08178_ (.B1(_03024_),
    .Y(_03025_),
    .A1(_01880_),
    .A2(net375));
 sg13g2_and2_1 _08179_ (.A(net376),
    .B(_03025_),
    .X(_00045_));
 sg13g2_nand2_1 _08180_ (.Y(_03026_),
    .A(_02923_),
    .B(_03017_));
 sg13g2_o21ai_1 _08181_ (.B1(_03026_),
    .Y(_03027_),
    .A1(_02375_),
    .A2(net375));
 sg13g2_and2_1 _08182_ (.A(net376),
    .B(_03027_),
    .X(_00046_));
 sg13g2_nand2_1 _08183_ (.Y(_03028_),
    .A(_02925_),
    .B(_03017_));
 sg13g2_o21ai_1 _08184_ (.B1(_03028_),
    .Y(_03029_),
    .A1(_02099_),
    .A2(net375));
 sg13g2_and2_1 _08185_ (.A(net376),
    .B(_03029_),
    .X(_00047_));
 sg13g2_nand2_1 _08186_ (.Y(_03030_),
    .A(_02927_),
    .B(_03017_));
 sg13g2_o21ai_1 _08187_ (.B1(_03030_),
    .Y(_03031_),
    .A1(_01869_),
    .A2(net375));
 sg13g2_and2_1 _08188_ (.A(_03011_),
    .B(_03031_),
    .X(_00048_));
 sg13g2_nand2_1 _08189_ (.Y(_03032_),
    .A(data_in_p2c_7),
    .B(_03017_));
 sg13g2_o21ai_1 _08190_ (.B1(_03032_),
    .Y(_03033_),
    .A1(_01865_),
    .A2(_03018_));
 sg13g2_and2_1 _08191_ (.A(_03011_),
    .B(_03033_),
    .X(_00049_));
 sg13g2_buf_1 _08192_ (.A(_02910_),
    .X(_03034_));
 sg13g2_nand2_1 _08193_ (.Y(_03035_),
    .A(_02932_),
    .B(_03017_));
 sg13g2_o21ai_1 _08194_ (.B1(_03035_),
    .Y(_03036_),
    .A1(_01867_),
    .A2(_03018_));
 sg13g2_and2_1 _08195_ (.A(_03034_),
    .B(_03036_),
    .X(_00050_));
 sg13g2_or2_1 _08196_ (.X(_03037_),
    .B(_03016_),
    .A(_02955_));
 sg13g2_buf_1 _08197_ (.A(_03037_),
    .X(_03038_));
 sg13g2_mux2_1 _08198_ (.A0(net493),
    .A1(net457),
    .S(net373),
    .X(_03039_));
 sg13g2_and2_1 _08199_ (.A(net374),
    .B(_03039_),
    .X(_00051_));
 sg13g2_mux2_1 _08200_ (.A0(net488),
    .A1(\median_processor.input_storage [57]),
    .S(net373),
    .X(_03040_));
 sg13g2_and2_1 _08201_ (.A(net374),
    .B(_03040_),
    .X(_00052_));
 sg13g2_nand2_1 _08202_ (.Y(_03041_),
    .A(net454),
    .B(net373));
 sg13g2_o21ai_1 _08203_ (.B1(_03041_),
    .Y(_03042_),
    .A1(_02920_),
    .A2(net373));
 sg13g2_and2_1 _08204_ (.A(net374),
    .B(_03042_),
    .X(_00053_));
 sg13g2_mux2_1 _08205_ (.A0(net492),
    .A1(net453),
    .S(net373),
    .X(_03043_));
 sg13g2_and2_1 _08206_ (.A(net374),
    .B(_03043_),
    .X(_00054_));
 sg13g2_mux2_1 _08207_ (.A0(net490),
    .A1(net422),
    .S(net385),
    .X(_03044_));
 sg13g2_and2_1 _08208_ (.A(net374),
    .B(_03044_),
    .X(_00055_));
 sg13g2_mux2_1 _08209_ (.A0(net491),
    .A1(\median_processor.input_storage [60]),
    .S(net373),
    .X(_03045_));
 sg13g2_and2_1 _08210_ (.A(net374),
    .B(_03045_),
    .X(_00056_));
 sg13g2_mux2_1 _08211_ (.A0(net490),
    .A1(net455),
    .S(net373),
    .X(_03046_));
 sg13g2_and2_1 _08212_ (.A(net374),
    .B(_03046_),
    .X(_00057_));
 sg13g2_nand2_1 _08213_ (.Y(_03047_),
    .A(net388),
    .B(net373));
 sg13g2_o21ai_1 _08214_ (.B1(_03047_),
    .Y(_03048_),
    .A1(_02929_),
    .A2(_03038_));
 sg13g2_and2_1 _08215_ (.A(net374),
    .B(_03048_),
    .X(_00058_));
 sg13g2_mux2_1 _08216_ (.A0(net489),
    .A1(net473),
    .S(_03038_),
    .X(_03049_));
 sg13g2_and2_1 _08217_ (.A(_03034_),
    .B(_03049_),
    .X(_00059_));
 sg13g2_buf_1 _08218_ (.A(net494),
    .X(_03050_));
 sg13g2_buf_1 _08219_ (.A(net411),
    .X(_03051_));
 sg13g2_buf_1 _08220_ (.A(net372),
    .X(_03052_));
 sg13g2_nand2_1 _08221_ (.Y(_03053_),
    .A(net440),
    .B(net385));
 sg13g2_o21ai_1 _08222_ (.B1(_03053_),
    .Y(_03054_),
    .A1(_02929_),
    .A2(_02916_));
 sg13g2_and2_1 _08223_ (.A(net221),
    .B(_03054_),
    .X(_00060_));
 sg13g2_mux2_1 _08224_ (.A0(net489),
    .A1(net472),
    .S(_02916_),
    .X(_03055_));
 sg13g2_and2_1 _08225_ (.A(net221),
    .B(_03055_),
    .X(_00061_));
 sg13g2_mux2_1 _08226_ (.A0(net493),
    .A1(net429),
    .S(net384),
    .X(_03056_));
 sg13g2_and2_1 _08227_ (.A(_03052_),
    .B(_03056_),
    .X(_00062_));
 sg13g2_mux2_1 _08228_ (.A0(net488),
    .A1(net428),
    .S(net384),
    .X(_03057_));
 sg13g2_and2_1 _08229_ (.A(_03052_),
    .B(_03057_),
    .X(_00063_));
 sg13g2_buf_2 _08230_ (.A(aux_enable_p2c),
    .X(_03058_));
 sg13g2_buf_1 _08231_ (.A(_03058_),
    .X(_03059_));
 sg13g2_buf_1 _08232_ (.A(net410),
    .X(_03060_));
 sg13g2_and2_1 _08233_ (.A(net494),
    .B(_03060_),
    .X(_03061_));
 sg13g2_buf_1 _08234_ (.A(_03061_),
    .X(_03062_));
 sg13g2_xnor2_1 _08235_ (.Y(_03063_),
    .A(\rando_generator.lfsr_reg [27]),
    .B(\rando_generator.lfsr_reg [30]));
 sg13g2_and2_1 _08236_ (.A(net32),
    .B(_03063_),
    .X(_00072_));
 sg13g2_and2_1 _08237_ (.A(\rando_generator.lfsr_reg [9]),
    .B(net32),
    .X(_00073_));
 sg13g2_and2_1 _08238_ (.A(\rando_generator.lfsr_reg [10]),
    .B(net32),
    .X(_00074_));
 sg13g2_and2_1 _08239_ (.A(\rando_generator.lfsr_reg [11]),
    .B(net32),
    .X(_00075_));
 sg13g2_and2_1 _08240_ (.A(\rando_generator.lfsr_reg [12]),
    .B(net32),
    .X(_00076_));
 sg13g2_and2_1 _08241_ (.A(\rando_generator.lfsr_reg [13]),
    .B(net32),
    .X(_00077_));
 sg13g2_and2_1 _08242_ (.A(\rando_generator.lfsr_reg [14]),
    .B(net32),
    .X(_00078_));
 sg13g2_and2_1 _08243_ (.A(\rando_generator.lfsr_reg [15]),
    .B(net32),
    .X(_00079_));
 sg13g2_and2_1 _08244_ (.A(\rando_generator.lfsr_reg [16]),
    .B(_03062_),
    .X(_00080_));
 sg13g2_and2_1 _08245_ (.A(\rando_generator.lfsr_reg [17]),
    .B(_03062_),
    .X(_00081_));
 sg13g2_buf_1 _08246_ (.A(_03061_),
    .X(_03064_));
 sg13g2_and2_1 _08247_ (.A(\rando_generator.lfsr_reg [18]),
    .B(net31),
    .X(_00082_));
 sg13g2_and2_1 _08248_ (.A(lfsr_out_c2p),
    .B(net31),
    .X(_00083_));
 sg13g2_and2_1 _08249_ (.A(\rando_generator.lfsr_reg [19]),
    .B(net31),
    .X(_00084_));
 sg13g2_and2_1 _08250_ (.A(\rando_generator.lfsr_reg [20]),
    .B(net31),
    .X(_00085_));
 sg13g2_and2_1 _08251_ (.A(\rando_generator.lfsr_reg [21]),
    .B(net31),
    .X(_00086_));
 sg13g2_and2_1 _08252_ (.A(\rando_generator.lfsr_reg [22]),
    .B(net31),
    .X(_00087_));
 sg13g2_and2_1 _08253_ (.A(\rando_generator.lfsr_reg [23]),
    .B(net31),
    .X(_00088_));
 sg13g2_and2_1 _08254_ (.A(\rando_generator.lfsr_reg [24]),
    .B(net31),
    .X(_00089_));
 sg13g2_and2_1 _08255_ (.A(\rando_generator.lfsr_reg [25]),
    .B(_03064_),
    .X(_00090_));
 sg13g2_and2_1 _08256_ (.A(\rando_generator.lfsr_reg [26]),
    .B(_03064_),
    .X(_00091_));
 sg13g2_buf_1 _08257_ (.A(_03061_),
    .X(_03065_));
 sg13g2_and2_1 _08258_ (.A(\rando_generator.lfsr_reg [27]),
    .B(net30),
    .X(_00092_));
 sg13g2_and2_1 _08259_ (.A(\rando_generator.lfsr_reg [28]),
    .B(net30),
    .X(_00093_));
 sg13g2_and2_1 _08260_ (.A(\rando_generator.lfsr_reg [1]),
    .B(net30),
    .X(_00094_));
 sg13g2_and2_1 _08261_ (.A(\rando_generator.lfsr_reg [29]),
    .B(net30),
    .X(_00095_));
 sg13g2_and2_1 _08262_ (.A(\rando_generator.lfsr_reg [2]),
    .B(net30),
    .X(_00096_));
 sg13g2_and2_1 _08263_ (.A(\rando_generator.lfsr_reg [3]),
    .B(net30),
    .X(_00097_));
 sg13g2_and2_1 _08264_ (.A(\rando_generator.lfsr_reg [4]),
    .B(net30),
    .X(_00098_));
 sg13g2_and2_1 _08265_ (.A(\rando_generator.lfsr_reg [5]),
    .B(net30),
    .X(_00099_));
 sg13g2_and2_1 _08266_ (.A(\rando_generator.lfsr_reg [6]),
    .B(_03065_),
    .X(_00100_));
 sg13g2_and2_1 _08267_ (.A(\rando_generator.lfsr_reg [7]),
    .B(_03065_),
    .X(_00101_));
 sg13g2_and2_1 _08268_ (.A(\rando_generator.lfsr_reg [8]),
    .B(_03061_),
    .X(_00102_));
 sg13g2_buf_1 _08269_ (.A(net371),
    .X(_03066_));
 sg13g2_mux2_1 _08270_ (.A0(\shift_storage.storage [0]),
    .A1(\shift_storage.shreg_in ),
    .S(_03066_),
    .X(_03067_));
 sg13g2_and2_1 _08271_ (.A(net221),
    .B(_03067_),
    .X(_00103_));
 sg13g2_mux2_1 _08272_ (.A0(\shift_storage.storage [1000]),
    .A1(\shift_storage.storage [999]),
    .S(net220),
    .X(_03068_));
 sg13g2_and2_1 _08273_ (.A(net221),
    .B(_03068_),
    .X(_00104_));
 sg13g2_mux2_1 _08274_ (.A0(\shift_storage.storage [1001]),
    .A1(\shift_storage.storage [1000]),
    .S(net220),
    .X(_03069_));
 sg13g2_and2_1 _08275_ (.A(net221),
    .B(_03069_),
    .X(_00105_));
 sg13g2_mux2_1 _08276_ (.A0(\shift_storage.storage [1002]),
    .A1(\shift_storage.storage [1001]),
    .S(net220),
    .X(_03070_));
 sg13g2_and2_1 _08277_ (.A(net221),
    .B(_03070_),
    .X(_00106_));
 sg13g2_mux2_1 _08278_ (.A0(\shift_storage.storage [1003]),
    .A1(\shift_storage.storage [1002]),
    .S(net220),
    .X(_03071_));
 sg13g2_and2_1 _08279_ (.A(net221),
    .B(_03071_),
    .X(_00107_));
 sg13g2_mux2_1 _08280_ (.A0(\shift_storage.storage [1004]),
    .A1(\shift_storage.storage [1003]),
    .S(net220),
    .X(_03072_));
 sg13g2_and2_1 _08281_ (.A(net221),
    .B(_03072_),
    .X(_00108_));
 sg13g2_buf_1 _08282_ (.A(net372),
    .X(_03073_));
 sg13g2_mux2_1 _08283_ (.A0(\shift_storage.storage [1005]),
    .A1(\shift_storage.storage [1004]),
    .S(net220),
    .X(_03074_));
 sg13g2_and2_1 _08284_ (.A(net219),
    .B(_03074_),
    .X(_00109_));
 sg13g2_mux2_1 _08285_ (.A0(\shift_storage.storage [1006]),
    .A1(\shift_storage.storage [1005]),
    .S(net220),
    .X(_03075_));
 sg13g2_and2_1 _08286_ (.A(net219),
    .B(_03075_),
    .X(_00110_));
 sg13g2_mux2_1 _08287_ (.A0(\shift_storage.storage [1007]),
    .A1(\shift_storage.storage [1006]),
    .S(_03066_),
    .X(_03076_));
 sg13g2_and2_1 _08288_ (.A(_03073_),
    .B(_03076_),
    .X(_00111_));
 sg13g2_mux2_1 _08289_ (.A0(\shift_storage.storage [1008]),
    .A1(\shift_storage.storage [1007]),
    .S(net220),
    .X(_03077_));
 sg13g2_and2_1 _08290_ (.A(_03073_),
    .B(_03077_),
    .X(_00112_));
 sg13g2_buf_1 _08291_ (.A(net371),
    .X(_03078_));
 sg13g2_mux2_1 _08292_ (.A0(\shift_storage.storage [1009]),
    .A1(\shift_storage.storage [1008]),
    .S(net218),
    .X(_03079_));
 sg13g2_and2_1 _08293_ (.A(net219),
    .B(_03079_),
    .X(_00113_));
 sg13g2_mux2_1 _08294_ (.A0(\shift_storage.storage [100]),
    .A1(\shift_storage.storage [99]),
    .S(net218),
    .X(_03080_));
 sg13g2_and2_1 _08295_ (.A(net219),
    .B(_03080_),
    .X(_00114_));
 sg13g2_mux2_1 _08296_ (.A0(\shift_storage.storage [1010]),
    .A1(\shift_storage.storage [1009]),
    .S(net218),
    .X(_03081_));
 sg13g2_and2_1 _08297_ (.A(net219),
    .B(_03081_),
    .X(_00115_));
 sg13g2_mux2_1 _08298_ (.A0(\shift_storage.storage [1011]),
    .A1(\shift_storage.storage [1010]),
    .S(net218),
    .X(_03082_));
 sg13g2_and2_1 _08299_ (.A(net219),
    .B(_03082_),
    .X(_00116_));
 sg13g2_mux2_1 _08300_ (.A0(\shift_storage.storage [1012]),
    .A1(\shift_storage.storage [1011]),
    .S(_03078_),
    .X(_03083_));
 sg13g2_and2_1 _08301_ (.A(net219),
    .B(_03083_),
    .X(_00117_));
 sg13g2_mux2_1 _08302_ (.A0(\shift_storage.storage [1013]),
    .A1(\shift_storage.storage [1012]),
    .S(_03078_),
    .X(_03084_));
 sg13g2_and2_1 _08303_ (.A(net219),
    .B(_03084_),
    .X(_00118_));
 sg13g2_buf_1 _08304_ (.A(net372),
    .X(_03085_));
 sg13g2_mux2_1 _08305_ (.A0(\shift_storage.storage [1014]),
    .A1(\shift_storage.storage [1013]),
    .S(net218),
    .X(_03086_));
 sg13g2_and2_1 _08306_ (.A(net217),
    .B(_03086_),
    .X(_00119_));
 sg13g2_mux2_1 _08307_ (.A0(\shift_storage.storage [1015]),
    .A1(\shift_storage.storage [1014]),
    .S(net218),
    .X(_03087_));
 sg13g2_and2_1 _08308_ (.A(net217),
    .B(_03087_),
    .X(_00120_));
 sg13g2_mux2_1 _08309_ (.A0(\shift_storage.storage [1016]),
    .A1(\shift_storage.storage [1015]),
    .S(net218),
    .X(_03088_));
 sg13g2_and2_1 _08310_ (.A(net217),
    .B(_03088_),
    .X(_00121_));
 sg13g2_mux2_1 _08311_ (.A0(\shift_storage.storage [1017]),
    .A1(\shift_storage.storage [1016]),
    .S(net218),
    .X(_03089_));
 sg13g2_and2_1 _08312_ (.A(_03085_),
    .B(_03089_),
    .X(_00122_));
 sg13g2_buf_1 _08313_ (.A(net371),
    .X(_03090_));
 sg13g2_mux2_1 _08314_ (.A0(\shift_storage.storage [1018]),
    .A1(\shift_storage.storage [1017]),
    .S(net216),
    .X(_03091_));
 sg13g2_and2_1 _08315_ (.A(net217),
    .B(_03091_),
    .X(_00123_));
 sg13g2_mux2_1 _08316_ (.A0(\shift_storage.storage [1019]),
    .A1(\shift_storage.storage [1018]),
    .S(net216),
    .X(_03092_));
 sg13g2_and2_1 _08317_ (.A(net217),
    .B(_03092_),
    .X(_00124_));
 sg13g2_mux2_1 _08318_ (.A0(\shift_storage.storage [101]),
    .A1(\shift_storage.storage [100]),
    .S(_03090_),
    .X(_03093_));
 sg13g2_and2_1 _08319_ (.A(_03085_),
    .B(_03093_),
    .X(_00125_));
 sg13g2_mux2_1 _08320_ (.A0(\shift_storage.storage [1020]),
    .A1(\shift_storage.storage [1019]),
    .S(net216),
    .X(_03094_));
 sg13g2_and2_1 _08321_ (.A(net217),
    .B(_03094_),
    .X(_00126_));
 sg13g2_mux2_1 _08322_ (.A0(\shift_storage.storage [1021]),
    .A1(\shift_storage.storage [1020]),
    .S(net216),
    .X(_03095_));
 sg13g2_and2_1 _08323_ (.A(net217),
    .B(_03095_),
    .X(_00127_));
 sg13g2_mux2_1 _08324_ (.A0(\shift_storage.storage [1022]),
    .A1(\shift_storage.storage [1021]),
    .S(net216),
    .X(_03096_));
 sg13g2_and2_1 _08325_ (.A(net217),
    .B(_03096_),
    .X(_00128_));
 sg13g2_buf_1 _08326_ (.A(net372),
    .X(_03097_));
 sg13g2_mux2_1 _08327_ (.A0(\shift_storage.storage [1023]),
    .A1(\shift_storage.storage [1022]),
    .S(net216),
    .X(_03098_));
 sg13g2_and2_1 _08328_ (.A(net215),
    .B(_03098_),
    .X(_00129_));
 sg13g2_mux2_1 _08329_ (.A0(\shift_storage.storage [1024]),
    .A1(\shift_storage.storage [1023]),
    .S(net216),
    .X(_03099_));
 sg13g2_and2_1 _08330_ (.A(net215),
    .B(_03099_),
    .X(_00130_));
 sg13g2_mux2_1 _08331_ (.A0(\shift_storage.storage [1025]),
    .A1(\shift_storage.storage [1024]),
    .S(net216),
    .X(_03100_));
 sg13g2_and2_1 _08332_ (.A(net215),
    .B(_03100_),
    .X(_00131_));
 sg13g2_mux2_1 _08333_ (.A0(\shift_storage.storage [1026]),
    .A1(\shift_storage.storage [1025]),
    .S(_03090_),
    .X(_03101_));
 sg13g2_and2_1 _08334_ (.A(net215),
    .B(_03101_),
    .X(_00132_));
 sg13g2_buf_1 _08335_ (.A(net371),
    .X(_03102_));
 sg13g2_mux2_1 _08336_ (.A0(\shift_storage.storage [1027]),
    .A1(\shift_storage.storage [1026]),
    .S(net214),
    .X(_03103_));
 sg13g2_and2_1 _08337_ (.A(_03097_),
    .B(_03103_),
    .X(_00133_));
 sg13g2_mux2_1 _08338_ (.A0(\shift_storage.storage [1028]),
    .A1(\shift_storage.storage [1027]),
    .S(net214),
    .X(_03104_));
 sg13g2_and2_1 _08339_ (.A(net215),
    .B(_03104_),
    .X(_00134_));
 sg13g2_mux2_1 _08340_ (.A0(\shift_storage.storage [1029]),
    .A1(\shift_storage.storage [1028]),
    .S(net214),
    .X(_03105_));
 sg13g2_and2_1 _08341_ (.A(net215),
    .B(_03105_),
    .X(_00135_));
 sg13g2_mux2_1 _08342_ (.A0(\shift_storage.storage [102]),
    .A1(\shift_storage.storage [101]),
    .S(net214),
    .X(_03106_));
 sg13g2_and2_1 _08343_ (.A(_03097_),
    .B(_03106_),
    .X(_00136_));
 sg13g2_mux2_1 _08344_ (.A0(\shift_storage.storage [1030]),
    .A1(\shift_storage.storage [1029]),
    .S(net214),
    .X(_03107_));
 sg13g2_and2_1 _08345_ (.A(net215),
    .B(_03107_),
    .X(_00137_));
 sg13g2_mux2_1 _08346_ (.A0(\shift_storage.storage [1031]),
    .A1(\shift_storage.storage [1030]),
    .S(net214),
    .X(_03108_));
 sg13g2_and2_1 _08347_ (.A(net215),
    .B(_03108_),
    .X(_00138_));
 sg13g2_buf_1 _08348_ (.A(net372),
    .X(_03109_));
 sg13g2_mux2_1 _08349_ (.A0(\shift_storage.storage [1032]),
    .A1(\shift_storage.storage [1031]),
    .S(net214),
    .X(_03110_));
 sg13g2_and2_1 _08350_ (.A(net213),
    .B(_03110_),
    .X(_00139_));
 sg13g2_mux2_1 _08351_ (.A0(\shift_storage.storage [1033]),
    .A1(\shift_storage.storage [1032]),
    .S(net214),
    .X(_03111_));
 sg13g2_and2_1 _08352_ (.A(net213),
    .B(_03111_),
    .X(_00140_));
 sg13g2_mux2_1 _08353_ (.A0(\shift_storage.storage [1034]),
    .A1(\shift_storage.storage [1033]),
    .S(_03102_),
    .X(_03112_));
 sg13g2_and2_1 _08354_ (.A(net213),
    .B(_03112_),
    .X(_00141_));
 sg13g2_mux2_1 _08355_ (.A0(\shift_storage.storage [1035]),
    .A1(\shift_storage.storage [1034]),
    .S(_03102_),
    .X(_03113_));
 sg13g2_and2_1 _08356_ (.A(net213),
    .B(_03113_),
    .X(_00142_));
 sg13g2_buf_1 _08357_ (.A(net371),
    .X(_03114_));
 sg13g2_mux2_1 _08358_ (.A0(\shift_storage.storage [1036]),
    .A1(\shift_storage.storage [1035]),
    .S(net212),
    .X(_03115_));
 sg13g2_and2_1 _08359_ (.A(net213),
    .B(_03115_),
    .X(_00143_));
 sg13g2_mux2_1 _08360_ (.A0(\shift_storage.storage [1037]),
    .A1(\shift_storage.storage [1036]),
    .S(net212),
    .X(_03116_));
 sg13g2_and2_1 _08361_ (.A(net213),
    .B(_03116_),
    .X(_00144_));
 sg13g2_mux2_1 _08362_ (.A0(\shift_storage.storage [1038]),
    .A1(\shift_storage.storage [1037]),
    .S(net212),
    .X(_03117_));
 sg13g2_and2_1 _08363_ (.A(net213),
    .B(_03117_),
    .X(_00145_));
 sg13g2_mux2_1 _08364_ (.A0(\shift_storage.storage [1039]),
    .A1(\shift_storage.storage [1038]),
    .S(net212),
    .X(_03118_));
 sg13g2_and2_1 _08365_ (.A(_03109_),
    .B(_03118_),
    .X(_00146_));
 sg13g2_mux2_1 _08366_ (.A0(\shift_storage.storage [103]),
    .A1(\shift_storage.storage [102]),
    .S(net212),
    .X(_03119_));
 sg13g2_and2_1 _08367_ (.A(net213),
    .B(_03119_),
    .X(_00147_));
 sg13g2_mux2_1 _08368_ (.A0(\shift_storage.storage [1040]),
    .A1(\shift_storage.storage [1039]),
    .S(net212),
    .X(_03120_));
 sg13g2_and2_1 _08369_ (.A(_03109_),
    .B(_03120_),
    .X(_00148_));
 sg13g2_buf_1 _08370_ (.A(net372),
    .X(_03121_));
 sg13g2_mux2_1 _08371_ (.A0(\shift_storage.storage [1041]),
    .A1(\shift_storage.storage [1040]),
    .S(net212),
    .X(_03122_));
 sg13g2_and2_1 _08372_ (.A(net211),
    .B(_03122_),
    .X(_00149_));
 sg13g2_mux2_1 _08373_ (.A0(\shift_storage.storage [1042]),
    .A1(\shift_storage.storage [1041]),
    .S(net212),
    .X(_03123_));
 sg13g2_and2_1 _08374_ (.A(net211),
    .B(_03123_),
    .X(_00150_));
 sg13g2_mux2_1 _08375_ (.A0(\shift_storage.storage [1043]),
    .A1(\shift_storage.storage [1042]),
    .S(_03114_),
    .X(_03124_));
 sg13g2_and2_1 _08376_ (.A(net211),
    .B(_03124_),
    .X(_00151_));
 sg13g2_mux2_1 _08377_ (.A0(\shift_storage.storage [1044]),
    .A1(\shift_storage.storage [1043]),
    .S(_03114_),
    .X(_03125_));
 sg13g2_and2_1 _08378_ (.A(net211),
    .B(_03125_),
    .X(_00152_));
 sg13g2_buf_1 _08379_ (.A(net371),
    .X(_03126_));
 sg13g2_mux2_1 _08380_ (.A0(\shift_storage.storage [1045]),
    .A1(\shift_storage.storage [1044]),
    .S(net210),
    .X(_03127_));
 sg13g2_and2_1 _08381_ (.A(net211),
    .B(_03127_),
    .X(_00153_));
 sg13g2_mux2_1 _08382_ (.A0(\shift_storage.storage [1046]),
    .A1(\shift_storage.storage [1045]),
    .S(net210),
    .X(_03128_));
 sg13g2_and2_1 _08383_ (.A(net211),
    .B(_03128_),
    .X(_00154_));
 sg13g2_mux2_1 _08384_ (.A0(\shift_storage.storage [1047]),
    .A1(\shift_storage.storage [1046]),
    .S(net210),
    .X(_03129_));
 sg13g2_and2_1 _08385_ (.A(net211),
    .B(_03129_),
    .X(_00155_));
 sg13g2_mux2_1 _08386_ (.A0(\shift_storage.storage [1048]),
    .A1(\shift_storage.storage [1047]),
    .S(net210),
    .X(_03130_));
 sg13g2_and2_1 _08387_ (.A(_03121_),
    .B(_03130_),
    .X(_00156_));
 sg13g2_mux2_1 _08388_ (.A0(\shift_storage.storage [1049]),
    .A1(\shift_storage.storage [1048]),
    .S(net210),
    .X(_03131_));
 sg13g2_and2_1 _08389_ (.A(_03121_),
    .B(_03131_),
    .X(_00157_));
 sg13g2_mux2_1 _08390_ (.A0(\shift_storage.storage [104]),
    .A1(\shift_storage.storage [103]),
    .S(_03126_),
    .X(_03132_));
 sg13g2_and2_1 _08391_ (.A(net211),
    .B(_03132_),
    .X(_00158_));
 sg13g2_buf_1 _08392_ (.A(net372),
    .X(_03133_));
 sg13g2_mux2_1 _08393_ (.A0(\shift_storage.storage [1050]),
    .A1(\shift_storage.storage [1049]),
    .S(net210),
    .X(_03134_));
 sg13g2_and2_1 _08394_ (.A(net209),
    .B(_03134_),
    .X(_00159_));
 sg13g2_mux2_1 _08395_ (.A0(\shift_storage.storage [1051]),
    .A1(\shift_storage.storage [1050]),
    .S(net210),
    .X(_03135_));
 sg13g2_and2_1 _08396_ (.A(net209),
    .B(_03135_),
    .X(_00160_));
 sg13g2_mux2_1 _08397_ (.A0(\shift_storage.storage [1052]),
    .A1(\shift_storage.storage [1051]),
    .S(net210),
    .X(_03136_));
 sg13g2_and2_1 _08398_ (.A(net209),
    .B(_03136_),
    .X(_00161_));
 sg13g2_mux2_1 _08399_ (.A0(\shift_storage.storage [1053]),
    .A1(\shift_storage.storage [1052]),
    .S(_03126_),
    .X(_03137_));
 sg13g2_and2_1 _08400_ (.A(_03133_),
    .B(_03137_),
    .X(_00162_));
 sg13g2_buf_1 _08401_ (.A(net371),
    .X(_03138_));
 sg13g2_mux2_1 _08402_ (.A0(\shift_storage.storage [1054]),
    .A1(\shift_storage.storage [1053]),
    .S(net208),
    .X(_03139_));
 sg13g2_and2_1 _08403_ (.A(_03133_),
    .B(_03139_),
    .X(_00163_));
 sg13g2_mux2_1 _08404_ (.A0(\shift_storage.storage [1055]),
    .A1(\shift_storage.storage [1054]),
    .S(net208),
    .X(_03140_));
 sg13g2_and2_1 _08405_ (.A(net209),
    .B(_03140_),
    .X(_00164_));
 sg13g2_mux2_1 _08406_ (.A0(\shift_storage.storage [1056]),
    .A1(\shift_storage.storage [1055]),
    .S(net208),
    .X(_03141_));
 sg13g2_and2_1 _08407_ (.A(net209),
    .B(_03141_),
    .X(_00165_));
 sg13g2_mux2_1 _08408_ (.A0(\shift_storage.storage [1057]),
    .A1(\shift_storage.storage [1056]),
    .S(net208),
    .X(_03142_));
 sg13g2_and2_1 _08409_ (.A(net209),
    .B(_03142_),
    .X(_00166_));
 sg13g2_mux2_1 _08410_ (.A0(\shift_storage.storage [1058]),
    .A1(\shift_storage.storage [1057]),
    .S(_03138_),
    .X(_03143_));
 sg13g2_and2_1 _08411_ (.A(net209),
    .B(_03143_),
    .X(_00167_));
 sg13g2_mux2_1 _08412_ (.A0(\shift_storage.storage [1059]),
    .A1(\shift_storage.storage [1058]),
    .S(_03138_),
    .X(_03144_));
 sg13g2_and2_1 _08413_ (.A(net209),
    .B(_03144_),
    .X(_00168_));
 sg13g2_buf_1 _08414_ (.A(net372),
    .X(_03145_));
 sg13g2_mux2_1 _08415_ (.A0(\shift_storage.storage [105]),
    .A1(\shift_storage.storage [104]),
    .S(net208),
    .X(_03146_));
 sg13g2_and2_1 _08416_ (.A(net207),
    .B(_03146_),
    .X(_00169_));
 sg13g2_mux2_1 _08417_ (.A0(\shift_storage.storage [1060]),
    .A1(\shift_storage.storage [1059]),
    .S(net208),
    .X(_03147_));
 sg13g2_and2_1 _08418_ (.A(net207),
    .B(_03147_),
    .X(_00170_));
 sg13g2_mux2_1 _08419_ (.A0(\shift_storage.storage [1061]),
    .A1(\shift_storage.storage [1060]),
    .S(net208),
    .X(_03148_));
 sg13g2_and2_1 _08420_ (.A(net207),
    .B(_03148_),
    .X(_00171_));
 sg13g2_mux2_1 _08421_ (.A0(\shift_storage.storage [1062]),
    .A1(\shift_storage.storage [1061]),
    .S(net208),
    .X(_03149_));
 sg13g2_and2_1 _08422_ (.A(net207),
    .B(_03149_),
    .X(_00172_));
 sg13g2_buf_1 _08423_ (.A(net371),
    .X(_03150_));
 sg13g2_mux2_1 _08424_ (.A0(\shift_storage.storage [1063]),
    .A1(\shift_storage.storage [1062]),
    .S(net206),
    .X(_03151_));
 sg13g2_and2_1 _08425_ (.A(net207),
    .B(_03151_),
    .X(_00173_));
 sg13g2_mux2_1 _08426_ (.A0(\shift_storage.storage [1064]),
    .A1(\shift_storage.storage [1063]),
    .S(net206),
    .X(_03152_));
 sg13g2_and2_1 _08427_ (.A(net207),
    .B(_03152_),
    .X(_00174_));
 sg13g2_mux2_1 _08428_ (.A0(\shift_storage.storage [1065]),
    .A1(\shift_storage.storage [1064]),
    .S(net206),
    .X(_03153_));
 sg13g2_and2_1 _08429_ (.A(net207),
    .B(_03153_),
    .X(_00175_));
 sg13g2_mux2_1 _08430_ (.A0(\shift_storage.storage [1066]),
    .A1(\shift_storage.storage [1065]),
    .S(_03150_),
    .X(_03154_));
 sg13g2_and2_1 _08431_ (.A(net207),
    .B(_03154_),
    .X(_00176_));
 sg13g2_mux2_1 _08432_ (.A0(\shift_storage.storage [1067]),
    .A1(\shift_storage.storage [1066]),
    .S(_03150_),
    .X(_03155_));
 sg13g2_and2_1 _08433_ (.A(_03145_),
    .B(_03155_),
    .X(_00177_));
 sg13g2_mux2_1 _08434_ (.A0(\shift_storage.storage [1068]),
    .A1(\shift_storage.storage [1067]),
    .S(net206),
    .X(_03156_));
 sg13g2_and2_1 _08435_ (.A(_03145_),
    .B(_03156_),
    .X(_00178_));
 sg13g2_buf_1 _08436_ (.A(_03051_),
    .X(_03157_));
 sg13g2_mux2_1 _08437_ (.A0(\shift_storage.storage [1069]),
    .A1(\shift_storage.storage [1068]),
    .S(net206),
    .X(_03158_));
 sg13g2_and2_1 _08438_ (.A(net205),
    .B(_03158_),
    .X(_00179_));
 sg13g2_mux2_1 _08439_ (.A0(\shift_storage.storage [106]),
    .A1(\shift_storage.storage [105]),
    .S(net206),
    .X(_03159_));
 sg13g2_and2_1 _08440_ (.A(net205),
    .B(_03159_),
    .X(_00180_));
 sg13g2_mux2_1 _08441_ (.A0(\shift_storage.storage [1070]),
    .A1(\shift_storage.storage [1069]),
    .S(net206),
    .X(_03160_));
 sg13g2_and2_1 _08442_ (.A(net205),
    .B(_03160_),
    .X(_00181_));
 sg13g2_mux2_1 _08443_ (.A0(\shift_storage.storage [1071]),
    .A1(\shift_storage.storage [1070]),
    .S(net206),
    .X(_03161_));
 sg13g2_and2_1 _08444_ (.A(net205),
    .B(_03161_),
    .X(_00182_));
 sg13g2_buf_1 _08445_ (.A(_03060_),
    .X(_03162_));
 sg13g2_mux2_1 _08446_ (.A0(\shift_storage.storage [1072]),
    .A1(\shift_storage.storage [1071]),
    .S(net204),
    .X(_03163_));
 sg13g2_and2_1 _08447_ (.A(net205),
    .B(_03163_),
    .X(_00183_));
 sg13g2_mux2_1 _08448_ (.A0(\shift_storage.storage [1073]),
    .A1(\shift_storage.storage [1072]),
    .S(net204),
    .X(_03164_));
 sg13g2_and2_1 _08449_ (.A(net205),
    .B(_03164_),
    .X(_00184_));
 sg13g2_mux2_1 _08450_ (.A0(\shift_storage.storage [1074]),
    .A1(\shift_storage.storage [1073]),
    .S(net204),
    .X(_03165_));
 sg13g2_and2_1 _08451_ (.A(_03157_),
    .B(_03165_),
    .X(_00185_));
 sg13g2_mux2_1 _08452_ (.A0(\shift_storage.storage [1075]),
    .A1(\shift_storage.storage [1074]),
    .S(_03162_),
    .X(_03166_));
 sg13g2_and2_1 _08453_ (.A(_03157_),
    .B(_03166_),
    .X(_00186_));
 sg13g2_mux2_1 _08454_ (.A0(\shift_storage.storage [1076]),
    .A1(\shift_storage.storage [1075]),
    .S(net204),
    .X(_03167_));
 sg13g2_and2_1 _08455_ (.A(net205),
    .B(_03167_),
    .X(_00187_));
 sg13g2_mux2_1 _08456_ (.A0(\shift_storage.storage [1077]),
    .A1(\shift_storage.storage [1076]),
    .S(net204),
    .X(_03168_));
 sg13g2_and2_1 _08457_ (.A(net205),
    .B(_03168_),
    .X(_00188_));
 sg13g2_buf_1 _08458_ (.A(_03051_),
    .X(_03169_));
 sg13g2_mux2_1 _08459_ (.A0(\shift_storage.storage [1078]),
    .A1(\shift_storage.storage [1077]),
    .S(net204),
    .X(_03170_));
 sg13g2_and2_1 _08460_ (.A(net203),
    .B(_03170_),
    .X(_00189_));
 sg13g2_mux2_1 _08461_ (.A0(\shift_storage.storage [1079]),
    .A1(\shift_storage.storage [1078]),
    .S(net204),
    .X(_03171_));
 sg13g2_and2_1 _08462_ (.A(net203),
    .B(_03171_),
    .X(_00190_));
 sg13g2_mux2_1 _08463_ (.A0(\shift_storage.storage [107]),
    .A1(\shift_storage.storage [106]),
    .S(net204),
    .X(_03172_));
 sg13g2_and2_1 _08464_ (.A(net203),
    .B(_03172_),
    .X(_00191_));
 sg13g2_mux2_1 _08465_ (.A0(\shift_storage.storage [1080]),
    .A1(\shift_storage.storage [1079]),
    .S(_03162_),
    .X(_03173_));
 sg13g2_and2_1 _08466_ (.A(_03169_),
    .B(_03173_),
    .X(_00192_));
 sg13g2_buf_1 _08467_ (.A(net410),
    .X(_03174_));
 sg13g2_buf_1 _08468_ (.A(net370),
    .X(_03175_));
 sg13g2_mux2_1 _08469_ (.A0(\shift_storage.storage [1081]),
    .A1(\shift_storage.storage [1080]),
    .S(net202),
    .X(_03176_));
 sg13g2_and2_1 _08470_ (.A(_03169_),
    .B(_03176_),
    .X(_00193_));
 sg13g2_mux2_1 _08471_ (.A0(\shift_storage.storage [1082]),
    .A1(\shift_storage.storage [1081]),
    .S(net202),
    .X(_03177_));
 sg13g2_and2_1 _08472_ (.A(net203),
    .B(_03177_),
    .X(_00194_));
 sg13g2_mux2_1 _08473_ (.A0(\shift_storage.storage [1083]),
    .A1(\shift_storage.storage [1082]),
    .S(net202),
    .X(_03178_));
 sg13g2_and2_1 _08474_ (.A(net203),
    .B(_03178_),
    .X(_00195_));
 sg13g2_mux2_1 _08475_ (.A0(\shift_storage.storage [1084]),
    .A1(\shift_storage.storage [1083]),
    .S(net202),
    .X(_03179_));
 sg13g2_and2_1 _08476_ (.A(net203),
    .B(_03179_),
    .X(_00196_));
 sg13g2_mux2_1 _08477_ (.A0(\shift_storage.storage [1085]),
    .A1(\shift_storage.storage [1084]),
    .S(_03175_),
    .X(_03180_));
 sg13g2_and2_1 _08478_ (.A(net203),
    .B(_03180_),
    .X(_00197_));
 sg13g2_mux2_1 _08479_ (.A0(\shift_storage.storage [1086]),
    .A1(\shift_storage.storage [1085]),
    .S(_03175_),
    .X(_03181_));
 sg13g2_and2_1 _08480_ (.A(net203),
    .B(_03181_),
    .X(_00198_));
 sg13g2_buf_1 _08481_ (.A(net411),
    .X(_03182_));
 sg13g2_buf_1 _08482_ (.A(net369),
    .X(_03183_));
 sg13g2_mux2_1 _08483_ (.A0(\shift_storage.storage [1087]),
    .A1(\shift_storage.storage [1086]),
    .S(net202),
    .X(_03184_));
 sg13g2_and2_1 _08484_ (.A(net201),
    .B(_03184_),
    .X(_00199_));
 sg13g2_mux2_1 _08485_ (.A0(\shift_storage.storage [1088]),
    .A1(\shift_storage.storage [1087]),
    .S(net202),
    .X(_03185_));
 sg13g2_and2_1 _08486_ (.A(net201),
    .B(_03185_),
    .X(_00200_));
 sg13g2_mux2_1 _08487_ (.A0(\shift_storage.storage [1089]),
    .A1(\shift_storage.storage [1088]),
    .S(net202),
    .X(_03186_));
 sg13g2_and2_1 _08488_ (.A(net201),
    .B(_03186_),
    .X(_00201_));
 sg13g2_mux2_1 _08489_ (.A0(\shift_storage.storage [108]),
    .A1(\shift_storage.storage [107]),
    .S(net202),
    .X(_03187_));
 sg13g2_and2_1 _08490_ (.A(_03183_),
    .B(_03187_),
    .X(_00202_));
 sg13g2_buf_1 _08491_ (.A(net370),
    .X(_03188_));
 sg13g2_mux2_1 _08492_ (.A0(\shift_storage.storage [1090]),
    .A1(\shift_storage.storage [1089]),
    .S(net200),
    .X(_03189_));
 sg13g2_and2_1 _08493_ (.A(_03183_),
    .B(_03189_),
    .X(_00203_));
 sg13g2_mux2_1 _08494_ (.A0(\shift_storage.storage [1091]),
    .A1(\shift_storage.storage [1090]),
    .S(net200),
    .X(_03190_));
 sg13g2_and2_1 _08495_ (.A(net201),
    .B(_03190_),
    .X(_00204_));
 sg13g2_mux2_1 _08496_ (.A0(\shift_storage.storage [1092]),
    .A1(\shift_storage.storage [1091]),
    .S(net200),
    .X(_03191_));
 sg13g2_and2_1 _08497_ (.A(net201),
    .B(_03191_),
    .X(_00205_));
 sg13g2_mux2_1 _08498_ (.A0(\shift_storage.storage [1093]),
    .A1(\shift_storage.storage [1092]),
    .S(net200),
    .X(_03192_));
 sg13g2_and2_1 _08499_ (.A(net201),
    .B(_03192_),
    .X(_00206_));
 sg13g2_mux2_1 _08500_ (.A0(\shift_storage.storage [1094]),
    .A1(\shift_storage.storage [1093]),
    .S(net200),
    .X(_03193_));
 sg13g2_and2_1 _08501_ (.A(net201),
    .B(_03193_),
    .X(_00207_));
 sg13g2_mux2_1 _08502_ (.A0(\shift_storage.storage [1095]),
    .A1(\shift_storage.storage [1094]),
    .S(net200),
    .X(_03194_));
 sg13g2_and2_1 _08503_ (.A(net201),
    .B(_03194_),
    .X(_00208_));
 sg13g2_buf_1 _08504_ (.A(net369),
    .X(_03195_));
 sg13g2_mux2_1 _08505_ (.A0(\shift_storage.storage [1096]),
    .A1(\shift_storage.storage [1095]),
    .S(net200),
    .X(_03196_));
 sg13g2_and2_1 _08506_ (.A(net199),
    .B(_03196_),
    .X(_00209_));
 sg13g2_mux2_1 _08507_ (.A0(\shift_storage.storage [1097]),
    .A1(\shift_storage.storage [1096]),
    .S(net200),
    .X(_03197_));
 sg13g2_and2_1 _08508_ (.A(net199),
    .B(_03197_),
    .X(_00210_));
 sg13g2_mux2_1 _08509_ (.A0(\shift_storage.storage [1098]),
    .A1(\shift_storage.storage [1097]),
    .S(_03188_),
    .X(_03198_));
 sg13g2_and2_1 _08510_ (.A(net199),
    .B(_03198_),
    .X(_00211_));
 sg13g2_mux2_1 _08511_ (.A0(\shift_storage.storage [1099]),
    .A1(\shift_storage.storage [1098]),
    .S(_03188_),
    .X(_03199_));
 sg13g2_and2_1 _08512_ (.A(net199),
    .B(_03199_),
    .X(_00212_));
 sg13g2_buf_1 _08513_ (.A(net370),
    .X(_03200_));
 sg13g2_mux2_1 _08514_ (.A0(\shift_storage.storage [109]),
    .A1(\shift_storage.storage [108]),
    .S(net198),
    .X(_03201_));
 sg13g2_and2_1 _08515_ (.A(net199),
    .B(_03201_),
    .X(_00213_));
 sg13g2_mux2_1 _08516_ (.A0(\shift_storage.storage [10]),
    .A1(\shift_storage.storage [9]),
    .S(net198),
    .X(_03202_));
 sg13g2_and2_1 _08517_ (.A(net199),
    .B(_03202_),
    .X(_00214_));
 sg13g2_mux2_1 _08518_ (.A0(\shift_storage.storage [1100]),
    .A1(\shift_storage.storage [1099]),
    .S(net198),
    .X(_03203_));
 sg13g2_and2_1 _08519_ (.A(net199),
    .B(_03203_),
    .X(_00215_));
 sg13g2_mux2_1 _08520_ (.A0(\shift_storage.storage [1101]),
    .A1(\shift_storage.storage [1100]),
    .S(net198),
    .X(_03204_));
 sg13g2_and2_1 _08521_ (.A(net199),
    .B(_03204_),
    .X(_00216_));
 sg13g2_mux2_1 _08522_ (.A0(\shift_storage.storage [1102]),
    .A1(\shift_storage.storage [1101]),
    .S(net198),
    .X(_03205_));
 sg13g2_and2_1 _08523_ (.A(_03195_),
    .B(_03205_),
    .X(_00217_));
 sg13g2_mux2_1 _08524_ (.A0(\shift_storage.storage [1103]),
    .A1(\shift_storage.storage [1102]),
    .S(net198),
    .X(_03206_));
 sg13g2_and2_1 _08525_ (.A(_03195_),
    .B(_03206_),
    .X(_00218_));
 sg13g2_buf_1 _08526_ (.A(net369),
    .X(_03207_));
 sg13g2_mux2_1 _08527_ (.A0(\shift_storage.storage [1104]),
    .A1(\shift_storage.storage [1103]),
    .S(net198),
    .X(_03208_));
 sg13g2_and2_1 _08528_ (.A(net197),
    .B(_03208_),
    .X(_00219_));
 sg13g2_mux2_1 _08529_ (.A0(\shift_storage.storage [1105]),
    .A1(\shift_storage.storage [1104]),
    .S(net198),
    .X(_03209_));
 sg13g2_and2_1 _08530_ (.A(net197),
    .B(_03209_),
    .X(_00220_));
 sg13g2_mux2_1 _08531_ (.A0(\shift_storage.storage [1106]),
    .A1(\shift_storage.storage [1105]),
    .S(_03200_),
    .X(_03210_));
 sg13g2_and2_1 _08532_ (.A(net197),
    .B(_03210_),
    .X(_00221_));
 sg13g2_mux2_1 _08533_ (.A0(\shift_storage.storage [1107]),
    .A1(\shift_storage.storage [1106]),
    .S(_03200_),
    .X(_03211_));
 sg13g2_and2_1 _08534_ (.A(net197),
    .B(_03211_),
    .X(_00222_));
 sg13g2_buf_1 _08535_ (.A(_03174_),
    .X(_03212_));
 sg13g2_mux2_1 _08536_ (.A0(\shift_storage.storage [1108]),
    .A1(\shift_storage.storage [1107]),
    .S(net196),
    .X(_03213_));
 sg13g2_and2_1 _08537_ (.A(net197),
    .B(_03213_),
    .X(_00223_));
 sg13g2_mux2_1 _08538_ (.A0(\shift_storage.storage [1109]),
    .A1(\shift_storage.storage [1108]),
    .S(net196),
    .X(_03214_));
 sg13g2_and2_1 _08539_ (.A(_03207_),
    .B(_03214_),
    .X(_00224_));
 sg13g2_mux2_1 _08540_ (.A0(\shift_storage.storage [110]),
    .A1(\shift_storage.storage [109]),
    .S(net196),
    .X(_03215_));
 sg13g2_and2_1 _08541_ (.A(net197),
    .B(_03215_),
    .X(_00225_));
 sg13g2_mux2_1 _08542_ (.A0(\shift_storage.storage [1110]),
    .A1(\shift_storage.storage [1109]),
    .S(net196),
    .X(_03216_));
 sg13g2_and2_1 _08543_ (.A(_03207_),
    .B(_03216_),
    .X(_00226_));
 sg13g2_mux2_1 _08544_ (.A0(\shift_storage.storage [1111]),
    .A1(\shift_storage.storage [1110]),
    .S(net196),
    .X(_03217_));
 sg13g2_and2_1 _08545_ (.A(net197),
    .B(_03217_),
    .X(_00227_));
 sg13g2_mux2_1 _08546_ (.A0(\shift_storage.storage [1112]),
    .A1(\shift_storage.storage [1111]),
    .S(net196),
    .X(_03218_));
 sg13g2_and2_1 _08547_ (.A(net197),
    .B(_03218_),
    .X(_00228_));
 sg13g2_buf_1 _08548_ (.A(net369),
    .X(_03219_));
 sg13g2_mux2_1 _08549_ (.A0(\shift_storage.storage [1113]),
    .A1(\shift_storage.storage [1112]),
    .S(_03212_),
    .X(_03220_));
 sg13g2_and2_1 _08550_ (.A(net195),
    .B(_03220_),
    .X(_00229_));
 sg13g2_mux2_1 _08551_ (.A0(\shift_storage.storage [1114]),
    .A1(\shift_storage.storage [1113]),
    .S(_03212_),
    .X(_03221_));
 sg13g2_and2_1 _08552_ (.A(net195),
    .B(_03221_),
    .X(_00230_));
 sg13g2_mux2_1 _08553_ (.A0(\shift_storage.storage [1115]),
    .A1(\shift_storage.storage [1114]),
    .S(net196),
    .X(_03222_));
 sg13g2_and2_1 _08554_ (.A(net195),
    .B(_03222_),
    .X(_00231_));
 sg13g2_mux2_1 _08555_ (.A0(\shift_storage.storage [1116]),
    .A1(\shift_storage.storage [1115]),
    .S(net196),
    .X(_03223_));
 sg13g2_and2_1 _08556_ (.A(net195),
    .B(_03223_),
    .X(_00232_));
 sg13g2_buf_1 _08557_ (.A(net370),
    .X(_03224_));
 sg13g2_mux2_1 _08558_ (.A0(\shift_storage.storage [1117]),
    .A1(\shift_storage.storage [1116]),
    .S(net194),
    .X(_03225_));
 sg13g2_and2_1 _08559_ (.A(net195),
    .B(_03225_),
    .X(_00233_));
 sg13g2_mux2_1 _08560_ (.A0(\shift_storage.storage [1118]),
    .A1(\shift_storage.storage [1117]),
    .S(net194),
    .X(_03226_));
 sg13g2_and2_1 _08561_ (.A(net195),
    .B(_03226_),
    .X(_00234_));
 sg13g2_mux2_1 _08562_ (.A0(\shift_storage.storage [1119]),
    .A1(\shift_storage.storage [1118]),
    .S(net194),
    .X(_03227_));
 sg13g2_and2_1 _08563_ (.A(net195),
    .B(_03227_),
    .X(_00235_));
 sg13g2_mux2_1 _08564_ (.A0(\shift_storage.storage [111]),
    .A1(\shift_storage.storage [110]),
    .S(net194),
    .X(_03228_));
 sg13g2_and2_1 _08565_ (.A(net195),
    .B(_03228_),
    .X(_00236_));
 sg13g2_mux2_1 _08566_ (.A0(\shift_storage.storage [1120]),
    .A1(\shift_storage.storage [1119]),
    .S(_03224_),
    .X(_03229_));
 sg13g2_and2_1 _08567_ (.A(_03219_),
    .B(_03229_),
    .X(_00237_));
 sg13g2_mux2_1 _08568_ (.A0(\shift_storage.storage [1121]),
    .A1(\shift_storage.storage [1120]),
    .S(_03224_),
    .X(_03230_));
 sg13g2_and2_1 _08569_ (.A(_03219_),
    .B(_03230_),
    .X(_00238_));
 sg13g2_buf_1 _08570_ (.A(net369),
    .X(_03231_));
 sg13g2_mux2_1 _08571_ (.A0(\shift_storage.storage [1122]),
    .A1(\shift_storage.storage [1121]),
    .S(net194),
    .X(_03232_));
 sg13g2_and2_1 _08572_ (.A(net193),
    .B(_03232_),
    .X(_00239_));
 sg13g2_mux2_1 _08573_ (.A0(\shift_storage.storage [1123]),
    .A1(\shift_storage.storage [1122]),
    .S(net194),
    .X(_03233_));
 sg13g2_and2_1 _08574_ (.A(net193),
    .B(_03233_),
    .X(_00240_));
 sg13g2_mux2_1 _08575_ (.A0(\shift_storage.storage [1124]),
    .A1(\shift_storage.storage [1123]),
    .S(net194),
    .X(_03234_));
 sg13g2_and2_1 _08576_ (.A(_03231_),
    .B(_03234_),
    .X(_00241_));
 sg13g2_mux2_1 _08577_ (.A0(\shift_storage.storage [1125]),
    .A1(\shift_storage.storage [1124]),
    .S(net194),
    .X(_03235_));
 sg13g2_and2_1 _08578_ (.A(_03231_),
    .B(_03235_),
    .X(_00242_));
 sg13g2_buf_1 _08579_ (.A(net370),
    .X(_03236_));
 sg13g2_mux2_1 _08580_ (.A0(\shift_storage.storage [1126]),
    .A1(\shift_storage.storage [1125]),
    .S(net192),
    .X(_03237_));
 sg13g2_and2_1 _08581_ (.A(net193),
    .B(_03237_),
    .X(_00243_));
 sg13g2_mux2_1 _08582_ (.A0(\shift_storage.storage [1127]),
    .A1(\shift_storage.storage [1126]),
    .S(net192),
    .X(_03238_));
 sg13g2_and2_1 _08583_ (.A(net193),
    .B(_03238_),
    .X(_00244_));
 sg13g2_mux2_1 _08584_ (.A0(\shift_storage.storage [1128]),
    .A1(\shift_storage.storage [1127]),
    .S(net192),
    .X(_03239_));
 sg13g2_and2_1 _08585_ (.A(net193),
    .B(_03239_),
    .X(_00245_));
 sg13g2_mux2_1 _08586_ (.A0(\shift_storage.storage [1129]),
    .A1(\shift_storage.storage [1128]),
    .S(net192),
    .X(_03240_));
 sg13g2_and2_1 _08587_ (.A(net193),
    .B(_03240_),
    .X(_00246_));
 sg13g2_mux2_1 _08588_ (.A0(\shift_storage.storage [112]),
    .A1(\shift_storage.storage [111]),
    .S(net192),
    .X(_03241_));
 sg13g2_and2_1 _08589_ (.A(net193),
    .B(_03241_),
    .X(_00247_));
 sg13g2_mux2_1 _08590_ (.A0(\shift_storage.storage [1130]),
    .A1(\shift_storage.storage [1129]),
    .S(net192),
    .X(_03242_));
 sg13g2_and2_1 _08591_ (.A(net193),
    .B(_03242_),
    .X(_00248_));
 sg13g2_buf_1 _08592_ (.A(_03182_),
    .X(_03243_));
 sg13g2_mux2_1 _08593_ (.A0(\shift_storage.storage [1131]),
    .A1(\shift_storage.storage [1130]),
    .S(net192),
    .X(_03244_));
 sg13g2_and2_1 _08594_ (.A(net191),
    .B(_03244_),
    .X(_00249_));
 sg13g2_mux2_1 _08595_ (.A0(\shift_storage.storage [1132]),
    .A1(\shift_storage.storage [1131]),
    .S(net192),
    .X(_03245_));
 sg13g2_and2_1 _08596_ (.A(net191),
    .B(_03245_),
    .X(_00250_));
 sg13g2_mux2_1 _08597_ (.A0(\shift_storage.storage [1133]),
    .A1(\shift_storage.storage [1132]),
    .S(_03236_),
    .X(_03246_));
 sg13g2_and2_1 _08598_ (.A(net191),
    .B(_03246_),
    .X(_00251_));
 sg13g2_mux2_1 _08599_ (.A0(\shift_storage.storage [1134]),
    .A1(\shift_storage.storage [1133]),
    .S(_03236_),
    .X(_03247_));
 sg13g2_and2_1 _08600_ (.A(net191),
    .B(_03247_),
    .X(_00252_));
 sg13g2_buf_1 _08601_ (.A(_03174_),
    .X(_03248_));
 sg13g2_mux2_1 _08602_ (.A0(\shift_storage.storage [1135]),
    .A1(\shift_storage.storage [1134]),
    .S(net190),
    .X(_03249_));
 sg13g2_and2_1 _08603_ (.A(_03243_),
    .B(_03249_),
    .X(_00253_));
 sg13g2_mux2_1 _08604_ (.A0(\shift_storage.storage [1136]),
    .A1(\shift_storage.storage [1135]),
    .S(net190),
    .X(_03250_));
 sg13g2_and2_1 _08605_ (.A(net191),
    .B(_03250_),
    .X(_00254_));
 sg13g2_mux2_1 _08606_ (.A0(\shift_storage.storage [1137]),
    .A1(\shift_storage.storage [1136]),
    .S(net190),
    .X(_03251_));
 sg13g2_and2_1 _08607_ (.A(net191),
    .B(_03251_),
    .X(_00255_));
 sg13g2_mux2_1 _08608_ (.A0(\shift_storage.storage [1138]),
    .A1(\shift_storage.storage [1137]),
    .S(_03248_),
    .X(_03252_));
 sg13g2_and2_1 _08609_ (.A(net191),
    .B(_03252_),
    .X(_00256_));
 sg13g2_mux2_1 _08610_ (.A0(\shift_storage.storage [1139]),
    .A1(\shift_storage.storage [1138]),
    .S(net190),
    .X(_03253_));
 sg13g2_and2_1 _08611_ (.A(net191),
    .B(_03253_),
    .X(_00257_));
 sg13g2_mux2_1 _08612_ (.A0(\shift_storage.storage [113]),
    .A1(\shift_storage.storage [112]),
    .S(_03248_),
    .X(_03254_));
 sg13g2_and2_1 _08613_ (.A(_03243_),
    .B(_03254_),
    .X(_00258_));
 sg13g2_buf_1 _08614_ (.A(_03182_),
    .X(_03255_));
 sg13g2_mux2_1 _08615_ (.A0(\shift_storage.storage [1140]),
    .A1(\shift_storage.storage [1139]),
    .S(net190),
    .X(_03256_));
 sg13g2_and2_1 _08616_ (.A(net189),
    .B(_03256_),
    .X(_00259_));
 sg13g2_mux2_1 _08617_ (.A0(\shift_storage.storage [1141]),
    .A1(\shift_storage.storage [1140]),
    .S(net190),
    .X(_03257_));
 sg13g2_and2_1 _08618_ (.A(net189),
    .B(_03257_),
    .X(_00260_));
 sg13g2_mux2_1 _08619_ (.A0(\shift_storage.storage [1142]),
    .A1(\shift_storage.storage [1141]),
    .S(net190),
    .X(_03258_));
 sg13g2_and2_1 _08620_ (.A(net189),
    .B(_03258_),
    .X(_00261_));
 sg13g2_mux2_1 _08621_ (.A0(\shift_storage.storage [1143]),
    .A1(\shift_storage.storage [1142]),
    .S(net190),
    .X(_03259_));
 sg13g2_and2_1 _08622_ (.A(net189),
    .B(_03259_),
    .X(_00262_));
 sg13g2_buf_1 _08623_ (.A(net370),
    .X(_03260_));
 sg13g2_mux2_1 _08624_ (.A0(\shift_storage.storage [1144]),
    .A1(\shift_storage.storage [1143]),
    .S(net188),
    .X(_03261_));
 sg13g2_and2_1 _08625_ (.A(net189),
    .B(_03261_),
    .X(_00263_));
 sg13g2_mux2_1 _08626_ (.A0(\shift_storage.storage [1145]),
    .A1(\shift_storage.storage [1144]),
    .S(net188),
    .X(_03262_));
 sg13g2_and2_1 _08627_ (.A(net189),
    .B(_03262_),
    .X(_00264_));
 sg13g2_mux2_1 _08628_ (.A0(\shift_storage.storage [1146]),
    .A1(\shift_storage.storage [1145]),
    .S(net188),
    .X(_03263_));
 sg13g2_and2_1 _08629_ (.A(net189),
    .B(_03263_),
    .X(_00265_));
 sg13g2_mux2_1 _08630_ (.A0(\shift_storage.storage [1147]),
    .A1(\shift_storage.storage [1146]),
    .S(net188),
    .X(_03264_));
 sg13g2_and2_1 _08631_ (.A(net189),
    .B(_03264_),
    .X(_00266_));
 sg13g2_mux2_1 _08632_ (.A0(\shift_storage.storage [1148]),
    .A1(\shift_storage.storage [1147]),
    .S(net188),
    .X(_03265_));
 sg13g2_and2_1 _08633_ (.A(_03255_),
    .B(_03265_),
    .X(_00267_));
 sg13g2_mux2_1 _08634_ (.A0(\shift_storage.storage [1149]),
    .A1(\shift_storage.storage [1148]),
    .S(net188),
    .X(_03266_));
 sg13g2_and2_1 _08635_ (.A(_03255_),
    .B(_03266_),
    .X(_00268_));
 sg13g2_buf_1 _08636_ (.A(net369),
    .X(_03267_));
 sg13g2_mux2_1 _08637_ (.A0(\shift_storage.storage [114]),
    .A1(\shift_storage.storage [113]),
    .S(_03260_),
    .X(_03268_));
 sg13g2_and2_1 _08638_ (.A(net187),
    .B(_03268_),
    .X(_00269_));
 sg13g2_mux2_1 _08639_ (.A0(\shift_storage.storage [1150]),
    .A1(\shift_storage.storage [1149]),
    .S(_03260_),
    .X(_03269_));
 sg13g2_and2_1 _08640_ (.A(net187),
    .B(_03269_),
    .X(_00270_));
 sg13g2_mux2_1 _08641_ (.A0(\shift_storage.storage [1151]),
    .A1(\shift_storage.storage [1150]),
    .S(net188),
    .X(_03270_));
 sg13g2_and2_1 _08642_ (.A(net187),
    .B(_03270_),
    .X(_00271_));
 sg13g2_mux2_1 _08643_ (.A0(\shift_storage.storage [1152]),
    .A1(\shift_storage.storage [1151]),
    .S(net188),
    .X(_03271_));
 sg13g2_and2_1 _08644_ (.A(net187),
    .B(_03271_),
    .X(_00272_));
 sg13g2_buf_1 _08645_ (.A(net370),
    .X(_03272_));
 sg13g2_mux2_1 _08646_ (.A0(\shift_storage.storage [1153]),
    .A1(\shift_storage.storage [1152]),
    .S(net186),
    .X(_03273_));
 sg13g2_and2_1 _08647_ (.A(net187),
    .B(_03273_),
    .X(_00273_));
 sg13g2_mux2_1 _08648_ (.A0(\shift_storage.storage [1154]),
    .A1(\shift_storage.storage [1153]),
    .S(net186),
    .X(_03274_));
 sg13g2_and2_1 _08649_ (.A(net187),
    .B(_03274_),
    .X(_00274_));
 sg13g2_mux2_1 _08650_ (.A0(\shift_storage.storage [1155]),
    .A1(\shift_storage.storage [1154]),
    .S(net186),
    .X(_03275_));
 sg13g2_and2_1 _08651_ (.A(net187),
    .B(_03275_),
    .X(_00275_));
 sg13g2_mux2_1 _08652_ (.A0(\shift_storage.storage [1156]),
    .A1(\shift_storage.storage [1155]),
    .S(net186),
    .X(_03276_));
 sg13g2_and2_1 _08653_ (.A(net187),
    .B(_03276_),
    .X(_00276_));
 sg13g2_mux2_1 _08654_ (.A0(\shift_storage.storage [1157]),
    .A1(\shift_storage.storage [1156]),
    .S(net186),
    .X(_03277_));
 sg13g2_and2_1 _08655_ (.A(_03267_),
    .B(_03277_),
    .X(_00277_));
 sg13g2_mux2_1 _08656_ (.A0(\shift_storage.storage [1158]),
    .A1(\shift_storage.storage [1157]),
    .S(net186),
    .X(_03278_));
 sg13g2_and2_1 _08657_ (.A(_03267_),
    .B(_03278_),
    .X(_00278_));
 sg13g2_buf_1 _08658_ (.A(net369),
    .X(_03279_));
 sg13g2_mux2_1 _08659_ (.A0(\shift_storage.storage [1159]),
    .A1(\shift_storage.storage [1158]),
    .S(net186),
    .X(_03280_));
 sg13g2_and2_1 _08660_ (.A(net185),
    .B(_03280_),
    .X(_00279_));
 sg13g2_mux2_1 _08661_ (.A0(\shift_storage.storage [115]),
    .A1(\shift_storage.storage [114]),
    .S(net186),
    .X(_03281_));
 sg13g2_and2_1 _08662_ (.A(net185),
    .B(_03281_),
    .X(_00280_));
 sg13g2_mux2_1 _08663_ (.A0(\shift_storage.storage [1160]),
    .A1(\shift_storage.storage [1159]),
    .S(_03272_),
    .X(_03282_));
 sg13g2_and2_1 _08664_ (.A(net185),
    .B(_03282_),
    .X(_00281_));
 sg13g2_mux2_1 _08665_ (.A0(\shift_storage.storage [1161]),
    .A1(\shift_storage.storage [1160]),
    .S(_03272_),
    .X(_03283_));
 sg13g2_and2_1 _08666_ (.A(net185),
    .B(_03283_),
    .X(_00282_));
 sg13g2_buf_1 _08667_ (.A(net370),
    .X(_03284_));
 sg13g2_mux2_1 _08668_ (.A0(\shift_storage.storage [1162]),
    .A1(\shift_storage.storage [1161]),
    .S(net184),
    .X(_03285_));
 sg13g2_and2_1 _08669_ (.A(net185),
    .B(_03285_),
    .X(_00283_));
 sg13g2_mux2_1 _08670_ (.A0(\shift_storage.storage [1163]),
    .A1(\shift_storage.storage [1162]),
    .S(net184),
    .X(_03286_));
 sg13g2_and2_1 _08671_ (.A(net185),
    .B(_03286_),
    .X(_00284_));
 sg13g2_mux2_1 _08672_ (.A0(\shift_storage.storage [1164]),
    .A1(\shift_storage.storage [1163]),
    .S(net184),
    .X(_03287_));
 sg13g2_and2_1 _08673_ (.A(net185),
    .B(_03287_),
    .X(_00285_));
 sg13g2_mux2_1 _08674_ (.A0(\shift_storage.storage [1165]),
    .A1(\shift_storage.storage [1164]),
    .S(net184),
    .X(_03288_));
 sg13g2_and2_1 _08675_ (.A(net185),
    .B(_03288_),
    .X(_00286_));
 sg13g2_mux2_1 _08676_ (.A0(\shift_storage.storage [1166]),
    .A1(\shift_storage.storage [1165]),
    .S(net184),
    .X(_03289_));
 sg13g2_and2_1 _08677_ (.A(_03279_),
    .B(_03289_),
    .X(_00287_));
 sg13g2_mux2_1 _08678_ (.A0(\shift_storage.storage [1167]),
    .A1(\shift_storage.storage [1166]),
    .S(net184),
    .X(_03290_));
 sg13g2_and2_1 _08679_ (.A(_03279_),
    .B(_03290_),
    .X(_00288_));
 sg13g2_buf_1 _08680_ (.A(net369),
    .X(_03291_));
 sg13g2_mux2_1 _08681_ (.A0(\shift_storage.storage [1168]),
    .A1(\shift_storage.storage [1167]),
    .S(net184),
    .X(_03292_));
 sg13g2_and2_1 _08682_ (.A(net183),
    .B(_03292_),
    .X(_00289_));
 sg13g2_mux2_1 _08683_ (.A0(\shift_storage.storage [1169]),
    .A1(\shift_storage.storage [1168]),
    .S(net184),
    .X(_03293_));
 sg13g2_and2_1 _08684_ (.A(net183),
    .B(_03293_),
    .X(_00290_));
 sg13g2_mux2_1 _08685_ (.A0(\shift_storage.storage [116]),
    .A1(\shift_storage.storage [115]),
    .S(_03284_),
    .X(_03294_));
 sg13g2_and2_1 _08686_ (.A(net183),
    .B(_03294_),
    .X(_00291_));
 sg13g2_mux2_1 _08687_ (.A0(\shift_storage.storage [1170]),
    .A1(\shift_storage.storage [1169]),
    .S(_03284_),
    .X(_03295_));
 sg13g2_and2_1 _08688_ (.A(net183),
    .B(_03295_),
    .X(_00292_));
 sg13g2_buf_1 _08689_ (.A(net410),
    .X(_03296_));
 sg13g2_buf_1 _08690_ (.A(net368),
    .X(_03297_));
 sg13g2_mux2_1 _08691_ (.A0(\shift_storage.storage [1171]),
    .A1(\shift_storage.storage [1170]),
    .S(net182),
    .X(_03298_));
 sg13g2_and2_1 _08692_ (.A(_03291_),
    .B(_03298_),
    .X(_00293_));
 sg13g2_mux2_1 _08693_ (.A0(\shift_storage.storage [1172]),
    .A1(\shift_storage.storage [1171]),
    .S(net182),
    .X(_03299_));
 sg13g2_and2_1 _08694_ (.A(_03291_),
    .B(_03299_),
    .X(_00294_));
 sg13g2_mux2_1 _08695_ (.A0(\shift_storage.storage [1173]),
    .A1(\shift_storage.storage [1172]),
    .S(_03297_),
    .X(_03300_));
 sg13g2_and2_1 _08696_ (.A(net183),
    .B(_03300_),
    .X(_00295_));
 sg13g2_mux2_1 _08697_ (.A0(\shift_storage.storage [1174]),
    .A1(\shift_storage.storage [1173]),
    .S(net182),
    .X(_03301_));
 sg13g2_and2_1 _08698_ (.A(net183),
    .B(_03301_),
    .X(_00296_));
 sg13g2_mux2_1 _08699_ (.A0(\shift_storage.storage [1175]),
    .A1(\shift_storage.storage [1174]),
    .S(net182),
    .X(_03302_));
 sg13g2_and2_1 _08700_ (.A(net183),
    .B(_03302_),
    .X(_00297_));
 sg13g2_mux2_1 _08701_ (.A0(\shift_storage.storage [1176]),
    .A1(\shift_storage.storage [1175]),
    .S(net182),
    .X(_03303_));
 sg13g2_and2_1 _08702_ (.A(net183),
    .B(_03303_),
    .X(_00298_));
 sg13g2_buf_1 _08703_ (.A(net411),
    .X(_03304_));
 sg13g2_buf_1 _08704_ (.A(net367),
    .X(_03305_));
 sg13g2_mux2_1 _08705_ (.A0(\shift_storage.storage [1177]),
    .A1(\shift_storage.storage [1176]),
    .S(net182),
    .X(_03306_));
 sg13g2_and2_1 _08706_ (.A(net181),
    .B(_03306_),
    .X(_00299_));
 sg13g2_mux2_1 _08707_ (.A0(\shift_storage.storage [1178]),
    .A1(\shift_storage.storage [1177]),
    .S(net182),
    .X(_03307_));
 sg13g2_and2_1 _08708_ (.A(net181),
    .B(_03307_),
    .X(_00300_));
 sg13g2_mux2_1 _08709_ (.A0(\shift_storage.storage [1179]),
    .A1(\shift_storage.storage [1178]),
    .S(net182),
    .X(_03308_));
 sg13g2_and2_1 _08710_ (.A(net181),
    .B(_03308_),
    .X(_00301_));
 sg13g2_mux2_1 _08711_ (.A0(\shift_storage.storage [117]),
    .A1(\shift_storage.storage [116]),
    .S(_03297_),
    .X(_03309_));
 sg13g2_and2_1 _08712_ (.A(net181),
    .B(_03309_),
    .X(_00302_));
 sg13g2_buf_1 _08713_ (.A(net368),
    .X(_03310_));
 sg13g2_mux2_1 _08714_ (.A0(\shift_storage.storage [1180]),
    .A1(\shift_storage.storage [1179]),
    .S(net180),
    .X(_03311_));
 sg13g2_and2_1 _08715_ (.A(net181),
    .B(_03311_),
    .X(_00303_));
 sg13g2_mux2_1 _08716_ (.A0(\shift_storage.storage [1181]),
    .A1(\shift_storage.storage [1180]),
    .S(net180),
    .X(_03312_));
 sg13g2_and2_1 _08717_ (.A(net181),
    .B(_03312_),
    .X(_00304_));
 sg13g2_mux2_1 _08718_ (.A0(\shift_storage.storage [1182]),
    .A1(\shift_storage.storage [1181]),
    .S(net180),
    .X(_03313_));
 sg13g2_and2_1 _08719_ (.A(net181),
    .B(_03313_),
    .X(_00305_));
 sg13g2_mux2_1 _08720_ (.A0(\shift_storage.storage [1183]),
    .A1(\shift_storage.storage [1182]),
    .S(net180),
    .X(_03314_));
 sg13g2_and2_1 _08721_ (.A(net181),
    .B(_03314_),
    .X(_00306_));
 sg13g2_mux2_1 _08722_ (.A0(\shift_storage.storage [1184]),
    .A1(\shift_storage.storage [1183]),
    .S(net180),
    .X(_03315_));
 sg13g2_and2_1 _08723_ (.A(_03305_),
    .B(_03315_),
    .X(_00307_));
 sg13g2_mux2_1 _08724_ (.A0(\shift_storage.storage [1185]),
    .A1(\shift_storage.storage [1184]),
    .S(net180),
    .X(_03316_));
 sg13g2_and2_1 _08725_ (.A(_03305_),
    .B(_03316_),
    .X(_00308_));
 sg13g2_buf_1 _08726_ (.A(net367),
    .X(_03317_));
 sg13g2_mux2_1 _08727_ (.A0(\shift_storage.storage [1186]),
    .A1(\shift_storage.storage [1185]),
    .S(net180),
    .X(_03318_));
 sg13g2_and2_1 _08728_ (.A(net179),
    .B(_03318_),
    .X(_00309_));
 sg13g2_mux2_1 _08729_ (.A0(\shift_storage.storage [1187]),
    .A1(\shift_storage.storage [1186]),
    .S(net180),
    .X(_03319_));
 sg13g2_and2_1 _08730_ (.A(net179),
    .B(_03319_),
    .X(_00310_));
 sg13g2_mux2_1 _08731_ (.A0(\shift_storage.storage [1188]),
    .A1(\shift_storage.storage [1187]),
    .S(_03310_),
    .X(_03320_));
 sg13g2_and2_1 _08732_ (.A(net179),
    .B(_03320_),
    .X(_00311_));
 sg13g2_mux2_1 _08733_ (.A0(\shift_storage.storage [1189]),
    .A1(\shift_storage.storage [1188]),
    .S(_03310_),
    .X(_03321_));
 sg13g2_and2_1 _08734_ (.A(net179),
    .B(_03321_),
    .X(_00312_));
 sg13g2_buf_1 _08735_ (.A(net368),
    .X(_03322_));
 sg13g2_mux2_1 _08736_ (.A0(\shift_storage.storage [118]),
    .A1(\shift_storage.storage [117]),
    .S(net178),
    .X(_03323_));
 sg13g2_and2_1 _08737_ (.A(net179),
    .B(_03323_),
    .X(_00313_));
 sg13g2_mux2_1 _08738_ (.A0(\shift_storage.storage [1190]),
    .A1(\shift_storage.storage [1189]),
    .S(net178),
    .X(_03324_));
 sg13g2_and2_1 _08739_ (.A(net179),
    .B(_03324_),
    .X(_00314_));
 sg13g2_mux2_1 _08740_ (.A0(\shift_storage.storage [1191]),
    .A1(\shift_storage.storage [1190]),
    .S(net178),
    .X(_03325_));
 sg13g2_and2_1 _08741_ (.A(net179),
    .B(_03325_),
    .X(_00315_));
 sg13g2_mux2_1 _08742_ (.A0(\shift_storage.storage [1192]),
    .A1(\shift_storage.storage [1191]),
    .S(net178),
    .X(_03326_));
 sg13g2_and2_1 _08743_ (.A(net179),
    .B(_03326_),
    .X(_00316_));
 sg13g2_mux2_1 _08744_ (.A0(\shift_storage.storage [1193]),
    .A1(\shift_storage.storage [1192]),
    .S(net178),
    .X(_03327_));
 sg13g2_and2_1 _08745_ (.A(_03317_),
    .B(_03327_),
    .X(_00317_));
 sg13g2_mux2_1 _08746_ (.A0(\shift_storage.storage [1194]),
    .A1(\shift_storage.storage [1193]),
    .S(net178),
    .X(_03328_));
 sg13g2_and2_1 _08747_ (.A(_03317_),
    .B(_03328_),
    .X(_00318_));
 sg13g2_buf_1 _08748_ (.A(_03304_),
    .X(_03329_));
 sg13g2_mux2_1 _08749_ (.A0(\shift_storage.storage [1195]),
    .A1(\shift_storage.storage [1194]),
    .S(net178),
    .X(_03330_));
 sg13g2_and2_1 _08750_ (.A(net177),
    .B(_03330_),
    .X(_00319_));
 sg13g2_mux2_1 _08751_ (.A0(\shift_storage.storage [1196]),
    .A1(\shift_storage.storage [1195]),
    .S(net178),
    .X(_03331_));
 sg13g2_and2_1 _08752_ (.A(net177),
    .B(_03331_),
    .X(_00320_));
 sg13g2_mux2_1 _08753_ (.A0(\shift_storage.storage [1197]),
    .A1(\shift_storage.storage [1196]),
    .S(_03322_),
    .X(_03332_));
 sg13g2_and2_1 _08754_ (.A(net177),
    .B(_03332_),
    .X(_00321_));
 sg13g2_mux2_1 _08755_ (.A0(\shift_storage.storage [1198]),
    .A1(\shift_storage.storage [1197]),
    .S(_03322_),
    .X(_03333_));
 sg13g2_and2_1 _08756_ (.A(net177),
    .B(_03333_),
    .X(_00322_));
 sg13g2_buf_1 _08757_ (.A(_03296_),
    .X(_03334_));
 sg13g2_mux2_1 _08758_ (.A0(\shift_storage.storage [1199]),
    .A1(\shift_storage.storage [1198]),
    .S(net176),
    .X(_03335_));
 sg13g2_and2_1 _08759_ (.A(net177),
    .B(_03335_),
    .X(_00323_));
 sg13g2_mux2_1 _08760_ (.A0(\shift_storage.storage [119]),
    .A1(\shift_storage.storage [118]),
    .S(net176),
    .X(_03336_));
 sg13g2_and2_1 _08761_ (.A(net177),
    .B(_03336_),
    .X(_00324_));
 sg13g2_mux2_1 _08762_ (.A0(\shift_storage.storage [11]),
    .A1(\shift_storage.storage [10]),
    .S(net176),
    .X(_03337_));
 sg13g2_and2_1 _08763_ (.A(net177),
    .B(_03337_),
    .X(_00325_));
 sg13g2_mux2_1 _08764_ (.A0(\shift_storage.storage [1200]),
    .A1(\shift_storage.storage [1199]),
    .S(net176),
    .X(_03338_));
 sg13g2_and2_1 _08765_ (.A(net177),
    .B(_03338_),
    .X(_00326_));
 sg13g2_mux2_1 _08766_ (.A0(\shift_storage.storage [1201]),
    .A1(\shift_storage.storage [1200]),
    .S(net176),
    .X(_03339_));
 sg13g2_and2_1 _08767_ (.A(_03329_),
    .B(_03339_),
    .X(_00327_));
 sg13g2_mux2_1 _08768_ (.A0(\shift_storage.storage [1202]),
    .A1(\shift_storage.storage [1201]),
    .S(net176),
    .X(_03340_));
 sg13g2_and2_1 _08769_ (.A(_03329_),
    .B(_03340_),
    .X(_00328_));
 sg13g2_buf_1 _08770_ (.A(_03304_),
    .X(_03341_));
 sg13g2_mux2_1 _08771_ (.A0(\shift_storage.storage [1203]),
    .A1(\shift_storage.storage [1202]),
    .S(net176),
    .X(_03342_));
 sg13g2_and2_1 _08772_ (.A(net175),
    .B(_03342_),
    .X(_00329_));
 sg13g2_mux2_1 _08773_ (.A0(\shift_storage.storage [1204]),
    .A1(\shift_storage.storage [1203]),
    .S(_03334_),
    .X(_03343_));
 sg13g2_and2_1 _08774_ (.A(_03341_),
    .B(_03343_),
    .X(_00330_));
 sg13g2_mux2_1 _08775_ (.A0(\shift_storage.storage [1205]),
    .A1(\shift_storage.storage [1204]),
    .S(_03334_),
    .X(_03344_));
 sg13g2_and2_1 _08776_ (.A(_03341_),
    .B(_03344_),
    .X(_00331_));
 sg13g2_mux2_1 _08777_ (.A0(\shift_storage.storage [1206]),
    .A1(\shift_storage.storage [1205]),
    .S(net176),
    .X(_03345_));
 sg13g2_and2_1 _08778_ (.A(net175),
    .B(_03345_),
    .X(_00332_));
 sg13g2_buf_1 _08779_ (.A(_03296_),
    .X(_03346_));
 sg13g2_mux2_1 _08780_ (.A0(\shift_storage.storage [1207]),
    .A1(\shift_storage.storage [1206]),
    .S(net174),
    .X(_03347_));
 sg13g2_and2_1 _08781_ (.A(net175),
    .B(_03347_),
    .X(_00333_));
 sg13g2_mux2_1 _08782_ (.A0(\shift_storage.storage [1208]),
    .A1(\shift_storage.storage [1207]),
    .S(net174),
    .X(_03348_));
 sg13g2_and2_1 _08783_ (.A(net175),
    .B(_03348_),
    .X(_00334_));
 sg13g2_mux2_1 _08784_ (.A0(\shift_storage.storage [1209]),
    .A1(\shift_storage.storage [1208]),
    .S(net174),
    .X(_03349_));
 sg13g2_and2_1 _08785_ (.A(net175),
    .B(_03349_),
    .X(_00335_));
 sg13g2_mux2_1 _08786_ (.A0(\shift_storage.storage [120]),
    .A1(\shift_storage.storage [119]),
    .S(_03346_),
    .X(_03350_));
 sg13g2_and2_1 _08787_ (.A(net175),
    .B(_03350_),
    .X(_00336_));
 sg13g2_mux2_1 _08788_ (.A0(\shift_storage.storage [1210]),
    .A1(\shift_storage.storage [1209]),
    .S(_03346_),
    .X(_03351_));
 sg13g2_and2_1 _08789_ (.A(net175),
    .B(_03351_),
    .X(_00337_));
 sg13g2_mux2_1 _08790_ (.A0(\shift_storage.storage [1211]),
    .A1(\shift_storage.storage [1210]),
    .S(net174),
    .X(_03352_));
 sg13g2_and2_1 _08791_ (.A(net175),
    .B(_03352_),
    .X(_00338_));
 sg13g2_buf_1 _08792_ (.A(net367),
    .X(_03353_));
 sg13g2_mux2_1 _08793_ (.A0(\shift_storage.storage [1212]),
    .A1(\shift_storage.storage [1211]),
    .S(net174),
    .X(_03354_));
 sg13g2_and2_1 _08794_ (.A(net173),
    .B(_03354_),
    .X(_00339_));
 sg13g2_mux2_1 _08795_ (.A0(\shift_storage.storage [1213]),
    .A1(\shift_storage.storage [1212]),
    .S(net174),
    .X(_03355_));
 sg13g2_and2_1 _08796_ (.A(net173),
    .B(_03355_),
    .X(_00340_));
 sg13g2_mux2_1 _08797_ (.A0(\shift_storage.storage [1214]),
    .A1(\shift_storage.storage [1213]),
    .S(net174),
    .X(_03356_));
 sg13g2_and2_1 _08798_ (.A(net173),
    .B(_03356_),
    .X(_00341_));
 sg13g2_mux2_1 _08799_ (.A0(\shift_storage.storage [1215]),
    .A1(\shift_storage.storage [1214]),
    .S(net174),
    .X(_03357_));
 sg13g2_and2_1 _08800_ (.A(net173),
    .B(_03357_),
    .X(_00342_));
 sg13g2_buf_1 _08801_ (.A(net368),
    .X(_03358_));
 sg13g2_mux2_1 _08802_ (.A0(\shift_storage.storage [1216]),
    .A1(\shift_storage.storage [1215]),
    .S(net172),
    .X(_03359_));
 sg13g2_and2_1 _08803_ (.A(net173),
    .B(_03359_),
    .X(_00343_));
 sg13g2_mux2_1 _08804_ (.A0(\shift_storage.storage [1217]),
    .A1(\shift_storage.storage [1216]),
    .S(net172),
    .X(_03360_));
 sg13g2_and2_1 _08805_ (.A(net173),
    .B(_03360_),
    .X(_00344_));
 sg13g2_mux2_1 _08806_ (.A0(\shift_storage.storage [1218]),
    .A1(\shift_storage.storage [1217]),
    .S(_03358_),
    .X(_03361_));
 sg13g2_and2_1 _08807_ (.A(net173),
    .B(_03361_),
    .X(_00345_));
 sg13g2_mux2_1 _08808_ (.A0(\shift_storage.storage [1219]),
    .A1(\shift_storage.storage [1218]),
    .S(net172),
    .X(_03362_));
 sg13g2_and2_1 _08809_ (.A(_03353_),
    .B(_03362_),
    .X(_00346_));
 sg13g2_mux2_1 _08810_ (.A0(\shift_storage.storage [121]),
    .A1(\shift_storage.storage [120]),
    .S(_03358_),
    .X(_03363_));
 sg13g2_and2_1 _08811_ (.A(net173),
    .B(_03363_),
    .X(_00347_));
 sg13g2_mux2_1 _08812_ (.A0(\shift_storage.storage [1220]),
    .A1(\shift_storage.storage [1219]),
    .S(net172),
    .X(_03364_));
 sg13g2_and2_1 _08813_ (.A(_03353_),
    .B(_03364_),
    .X(_00348_));
 sg13g2_buf_1 _08814_ (.A(net367),
    .X(_03365_));
 sg13g2_mux2_1 _08815_ (.A0(\shift_storage.storage [1221]),
    .A1(\shift_storage.storage [1220]),
    .S(net172),
    .X(_03366_));
 sg13g2_and2_1 _08816_ (.A(net171),
    .B(_03366_),
    .X(_00349_));
 sg13g2_mux2_1 _08817_ (.A0(\shift_storage.storage [1222]),
    .A1(\shift_storage.storage [1221]),
    .S(net172),
    .X(_03367_));
 sg13g2_and2_1 _08818_ (.A(net171),
    .B(_03367_),
    .X(_00350_));
 sg13g2_mux2_1 _08819_ (.A0(\shift_storage.storage [1223]),
    .A1(\shift_storage.storage [1222]),
    .S(net172),
    .X(_03368_));
 sg13g2_and2_1 _08820_ (.A(_03365_),
    .B(_03368_),
    .X(_00351_));
 sg13g2_mux2_1 _08821_ (.A0(\shift_storage.storage [1224]),
    .A1(\shift_storage.storage [1223]),
    .S(net172),
    .X(_03369_));
 sg13g2_and2_1 _08822_ (.A(net171),
    .B(_03369_),
    .X(_00352_));
 sg13g2_buf_1 _08823_ (.A(net368),
    .X(_03370_));
 sg13g2_mux2_1 _08824_ (.A0(\shift_storage.storage [1225]),
    .A1(\shift_storage.storage [1224]),
    .S(net170),
    .X(_03371_));
 sg13g2_and2_1 _08825_ (.A(net171),
    .B(_03371_),
    .X(_00353_));
 sg13g2_mux2_1 _08826_ (.A0(\shift_storage.storage [1226]),
    .A1(\shift_storage.storage [1225]),
    .S(net170),
    .X(_03372_));
 sg13g2_and2_1 _08827_ (.A(net171),
    .B(_03372_),
    .X(_00354_));
 sg13g2_mux2_1 _08828_ (.A0(\shift_storage.storage [1227]),
    .A1(\shift_storage.storage [1226]),
    .S(net170),
    .X(_03373_));
 sg13g2_and2_1 _08829_ (.A(net171),
    .B(_03373_),
    .X(_00355_));
 sg13g2_mux2_1 _08830_ (.A0(\shift_storage.storage [1228]),
    .A1(\shift_storage.storage [1227]),
    .S(_03370_),
    .X(_03374_));
 sg13g2_and2_1 _08831_ (.A(net171),
    .B(_03374_),
    .X(_00356_));
 sg13g2_mux2_1 _08832_ (.A0(\shift_storage.storage [1229]),
    .A1(\shift_storage.storage [1228]),
    .S(net170),
    .X(_03375_));
 sg13g2_and2_1 _08833_ (.A(net171),
    .B(_03375_),
    .X(_00357_));
 sg13g2_mux2_1 _08834_ (.A0(\shift_storage.storage [122]),
    .A1(\shift_storage.storage [121]),
    .S(_03370_),
    .X(_03376_));
 sg13g2_and2_1 _08835_ (.A(_03365_),
    .B(_03376_),
    .X(_00358_));
 sg13g2_buf_1 _08836_ (.A(net367),
    .X(_03377_));
 sg13g2_mux2_1 _08837_ (.A0(\shift_storage.storage [1230]),
    .A1(\shift_storage.storage [1229]),
    .S(net170),
    .X(_03378_));
 sg13g2_and2_1 _08838_ (.A(net169),
    .B(_03378_),
    .X(_00359_));
 sg13g2_mux2_1 _08839_ (.A0(\shift_storage.storage [1231]),
    .A1(\shift_storage.storage [1230]),
    .S(net170),
    .X(_03379_));
 sg13g2_and2_1 _08840_ (.A(net169),
    .B(_03379_),
    .X(_00360_));
 sg13g2_mux2_1 _08841_ (.A0(\shift_storage.storage [1232]),
    .A1(\shift_storage.storage [1231]),
    .S(net170),
    .X(_03380_));
 sg13g2_and2_1 _08842_ (.A(net169),
    .B(_03380_),
    .X(_00361_));
 sg13g2_mux2_1 _08843_ (.A0(\shift_storage.storage [1233]),
    .A1(\shift_storage.storage [1232]),
    .S(net170),
    .X(_03381_));
 sg13g2_and2_1 _08844_ (.A(_03377_),
    .B(_03381_),
    .X(_00362_));
 sg13g2_buf_1 _08845_ (.A(net368),
    .X(_03382_));
 sg13g2_mux2_1 _08846_ (.A0(\shift_storage.storage [1234]),
    .A1(\shift_storage.storage [1233]),
    .S(_03382_),
    .X(_03383_));
 sg13g2_and2_1 _08847_ (.A(_03377_),
    .B(_03383_),
    .X(_00363_));
 sg13g2_mux2_1 _08848_ (.A0(\shift_storage.storage [1235]),
    .A1(\shift_storage.storage [1234]),
    .S(net168),
    .X(_03384_));
 sg13g2_and2_1 _08849_ (.A(net169),
    .B(_03384_),
    .X(_00364_));
 sg13g2_mux2_1 _08850_ (.A0(\shift_storage.storage [1236]),
    .A1(\shift_storage.storage [1235]),
    .S(net168),
    .X(_03385_));
 sg13g2_and2_1 _08851_ (.A(net169),
    .B(_03385_),
    .X(_00365_));
 sg13g2_mux2_1 _08852_ (.A0(\shift_storage.storage [1237]),
    .A1(\shift_storage.storage [1236]),
    .S(net168),
    .X(_03386_));
 sg13g2_and2_1 _08853_ (.A(net169),
    .B(_03386_),
    .X(_00366_));
 sg13g2_mux2_1 _08854_ (.A0(\shift_storage.storage [1238]),
    .A1(\shift_storage.storage [1237]),
    .S(net168),
    .X(_03387_));
 sg13g2_and2_1 _08855_ (.A(net169),
    .B(_03387_),
    .X(_00367_));
 sg13g2_mux2_1 _08856_ (.A0(\shift_storage.storage [1239]),
    .A1(\shift_storage.storage [1238]),
    .S(net168),
    .X(_03388_));
 sg13g2_and2_1 _08857_ (.A(net169),
    .B(_03388_),
    .X(_00368_));
 sg13g2_buf_1 _08858_ (.A(net367),
    .X(_03389_));
 sg13g2_mux2_1 _08859_ (.A0(\shift_storage.storage [123]),
    .A1(\shift_storage.storage [122]),
    .S(_03382_),
    .X(_03390_));
 sg13g2_and2_1 _08860_ (.A(net167),
    .B(_03390_),
    .X(_00369_));
 sg13g2_mux2_1 _08861_ (.A0(\shift_storage.storage [1240]),
    .A1(\shift_storage.storage [1239]),
    .S(net168),
    .X(_03391_));
 sg13g2_and2_1 _08862_ (.A(net167),
    .B(_03391_),
    .X(_00370_));
 sg13g2_mux2_1 _08863_ (.A0(\shift_storage.storage [1241]),
    .A1(\shift_storage.storage [1240]),
    .S(net168),
    .X(_03392_));
 sg13g2_and2_1 _08864_ (.A(net167),
    .B(_03392_),
    .X(_00371_));
 sg13g2_mux2_1 _08865_ (.A0(\shift_storage.storage [1242]),
    .A1(\shift_storage.storage [1241]),
    .S(net168),
    .X(_03393_));
 sg13g2_and2_1 _08866_ (.A(net167),
    .B(_03393_),
    .X(_00372_));
 sg13g2_buf_1 _08867_ (.A(net368),
    .X(_03394_));
 sg13g2_mux2_1 _08868_ (.A0(\shift_storage.storage [1243]),
    .A1(\shift_storage.storage [1242]),
    .S(net166),
    .X(_03395_));
 sg13g2_and2_1 _08869_ (.A(_03389_),
    .B(_03395_),
    .X(_00373_));
 sg13g2_mux2_1 _08870_ (.A0(\shift_storage.storage [1244]),
    .A1(\shift_storage.storage [1243]),
    .S(_03394_),
    .X(_03396_));
 sg13g2_and2_1 _08871_ (.A(_03389_),
    .B(_03396_),
    .X(_00374_));
 sg13g2_mux2_1 _08872_ (.A0(\shift_storage.storage [1245]),
    .A1(\shift_storage.storage [1244]),
    .S(net166),
    .X(_03397_));
 sg13g2_and2_1 _08873_ (.A(net167),
    .B(_03397_),
    .X(_00375_));
 sg13g2_mux2_1 _08874_ (.A0(\shift_storage.storage [1246]),
    .A1(\shift_storage.storage [1245]),
    .S(net166),
    .X(_03398_));
 sg13g2_and2_1 _08875_ (.A(net167),
    .B(_03398_),
    .X(_00376_));
 sg13g2_mux2_1 _08876_ (.A0(\shift_storage.storage [1247]),
    .A1(\shift_storage.storage [1246]),
    .S(net166),
    .X(_03399_));
 sg13g2_and2_1 _08877_ (.A(net167),
    .B(_03399_),
    .X(_00377_));
 sg13g2_mux2_1 _08878_ (.A0(\shift_storage.storage [1248]),
    .A1(\shift_storage.storage [1247]),
    .S(net166),
    .X(_03400_));
 sg13g2_and2_1 _08879_ (.A(net167),
    .B(_03400_),
    .X(_00378_));
 sg13g2_buf_1 _08880_ (.A(net367),
    .X(_03401_));
 sg13g2_mux2_1 _08881_ (.A0(\shift_storage.storage [1249]),
    .A1(\shift_storage.storage [1248]),
    .S(net166),
    .X(_03402_));
 sg13g2_and2_1 _08882_ (.A(net165),
    .B(_03402_),
    .X(_00379_));
 sg13g2_mux2_1 _08883_ (.A0(\shift_storage.storage [124]),
    .A1(\shift_storage.storage [123]),
    .S(_03394_),
    .X(_03403_));
 sg13g2_and2_1 _08884_ (.A(net165),
    .B(_03403_),
    .X(_00380_));
 sg13g2_mux2_1 _08885_ (.A0(\shift_storage.storage [1250]),
    .A1(\shift_storage.storage [1249]),
    .S(net166),
    .X(_03404_));
 sg13g2_and2_1 _08886_ (.A(net165),
    .B(_03404_),
    .X(_00381_));
 sg13g2_mux2_1 _08887_ (.A0(\shift_storage.storage [1251]),
    .A1(\shift_storage.storage [1250]),
    .S(net166),
    .X(_03405_));
 sg13g2_and2_1 _08888_ (.A(net165),
    .B(_03405_),
    .X(_00382_));
 sg13g2_buf_1 _08889_ (.A(net368),
    .X(_03406_));
 sg13g2_mux2_1 _08890_ (.A0(\shift_storage.storage [1252]),
    .A1(\shift_storage.storage [1251]),
    .S(net164),
    .X(_03407_));
 sg13g2_and2_1 _08891_ (.A(net165),
    .B(_03407_),
    .X(_00383_));
 sg13g2_mux2_1 _08892_ (.A0(\shift_storage.storage [1253]),
    .A1(\shift_storage.storage [1252]),
    .S(net164),
    .X(_03408_));
 sg13g2_and2_1 _08893_ (.A(net165),
    .B(_03408_),
    .X(_00384_));
 sg13g2_mux2_1 _08894_ (.A0(\shift_storage.storage [1254]),
    .A1(\shift_storage.storage [1253]),
    .S(net164),
    .X(_03409_));
 sg13g2_and2_1 _08895_ (.A(net165),
    .B(_03409_),
    .X(_00385_));
 sg13g2_mux2_1 _08896_ (.A0(\shift_storage.storage [1255]),
    .A1(\shift_storage.storage [1254]),
    .S(net164),
    .X(_03410_));
 sg13g2_and2_1 _08897_ (.A(net165),
    .B(_03410_),
    .X(_00386_));
 sg13g2_mux2_1 _08898_ (.A0(\shift_storage.storage [1256]),
    .A1(\shift_storage.storage [1255]),
    .S(net164),
    .X(_03411_));
 sg13g2_and2_1 _08899_ (.A(_03401_),
    .B(_03411_),
    .X(_00387_));
 sg13g2_mux2_1 _08900_ (.A0(\shift_storage.storage [1257]),
    .A1(\shift_storage.storage [1256]),
    .S(net164),
    .X(_03412_));
 sg13g2_and2_1 _08901_ (.A(_03401_),
    .B(_03412_),
    .X(_00388_));
 sg13g2_buf_1 _08902_ (.A(net367),
    .X(_03413_));
 sg13g2_mux2_1 _08903_ (.A0(\shift_storage.storage [1258]),
    .A1(\shift_storage.storage [1257]),
    .S(net164),
    .X(_03414_));
 sg13g2_and2_1 _08904_ (.A(net163),
    .B(_03414_),
    .X(_00389_));
 sg13g2_mux2_1 _08905_ (.A0(\shift_storage.storage [1259]),
    .A1(\shift_storage.storage [1258]),
    .S(net164),
    .X(_03415_));
 sg13g2_and2_1 _08906_ (.A(net163),
    .B(_03415_),
    .X(_00390_));
 sg13g2_mux2_1 _08907_ (.A0(\shift_storage.storage [125]),
    .A1(\shift_storage.storage [124]),
    .S(_03406_),
    .X(_03416_));
 sg13g2_and2_1 _08908_ (.A(net163),
    .B(_03416_),
    .X(_00391_));
 sg13g2_mux2_1 _08909_ (.A0(\shift_storage.storage [1260]),
    .A1(\shift_storage.storage [1259]),
    .S(_03406_),
    .X(_03417_));
 sg13g2_and2_1 _08910_ (.A(net163),
    .B(_03417_),
    .X(_00392_));
 sg13g2_buf_1 _08911_ (.A(net410),
    .X(_03418_));
 sg13g2_buf_1 _08912_ (.A(net366),
    .X(_03419_));
 sg13g2_mux2_1 _08913_ (.A0(\shift_storage.storage [1261]),
    .A1(\shift_storage.storage [1260]),
    .S(net162),
    .X(_03420_));
 sg13g2_and2_1 _08914_ (.A(net163),
    .B(_03420_),
    .X(_00393_));
 sg13g2_mux2_1 _08915_ (.A0(\shift_storage.storage [1262]),
    .A1(\shift_storage.storage [1261]),
    .S(net162),
    .X(_03421_));
 sg13g2_and2_1 _08916_ (.A(net163),
    .B(_03421_),
    .X(_00394_));
 sg13g2_mux2_1 _08917_ (.A0(\shift_storage.storage [1263]),
    .A1(\shift_storage.storage [1262]),
    .S(net162),
    .X(_03422_));
 sg13g2_and2_1 _08918_ (.A(net163),
    .B(_03422_),
    .X(_00395_));
 sg13g2_mux2_1 _08919_ (.A0(\shift_storage.storage [1264]),
    .A1(\shift_storage.storage [1263]),
    .S(net162),
    .X(_03423_));
 sg13g2_and2_1 _08920_ (.A(net163),
    .B(_03423_),
    .X(_00396_));
 sg13g2_mux2_1 _08921_ (.A0(\shift_storage.storage [1265]),
    .A1(\shift_storage.storage [1264]),
    .S(net162),
    .X(_03424_));
 sg13g2_and2_1 _08922_ (.A(_03413_),
    .B(_03424_),
    .X(_00397_));
 sg13g2_mux2_1 _08923_ (.A0(\shift_storage.storage [1266]),
    .A1(\shift_storage.storage [1265]),
    .S(net162),
    .X(_03425_));
 sg13g2_and2_1 _08924_ (.A(_03413_),
    .B(_03425_),
    .X(_00398_));
 sg13g2_buf_1 _08925_ (.A(net411),
    .X(_03426_));
 sg13g2_buf_1 _08926_ (.A(net365),
    .X(_03427_));
 sg13g2_mux2_1 _08927_ (.A0(\shift_storage.storage [1267]),
    .A1(\shift_storage.storage [1266]),
    .S(net162),
    .X(_03428_));
 sg13g2_and2_1 _08928_ (.A(net161),
    .B(_03428_),
    .X(_00399_));
 sg13g2_mux2_1 _08929_ (.A0(\shift_storage.storage [1268]),
    .A1(\shift_storage.storage [1267]),
    .S(net162),
    .X(_03429_));
 sg13g2_and2_1 _08930_ (.A(net161),
    .B(_03429_),
    .X(_00400_));
 sg13g2_mux2_1 _08931_ (.A0(\shift_storage.storage [1269]),
    .A1(\shift_storage.storage [1268]),
    .S(_03419_),
    .X(_03430_));
 sg13g2_and2_1 _08932_ (.A(net161),
    .B(_03430_),
    .X(_00401_));
 sg13g2_mux2_1 _08933_ (.A0(\shift_storage.storage [126]),
    .A1(\shift_storage.storage [125]),
    .S(_03419_),
    .X(_03431_));
 sg13g2_and2_1 _08934_ (.A(net161),
    .B(_03431_),
    .X(_00402_));
 sg13g2_buf_1 _08935_ (.A(net366),
    .X(_03432_));
 sg13g2_mux2_1 _08936_ (.A0(\shift_storage.storage [1270]),
    .A1(\shift_storage.storage [1269]),
    .S(net160),
    .X(_03433_));
 sg13g2_and2_1 _08937_ (.A(net161),
    .B(_03433_),
    .X(_00403_));
 sg13g2_mux2_1 _08938_ (.A0(\shift_storage.storage [1271]),
    .A1(\shift_storage.storage [1270]),
    .S(net160),
    .X(_03434_));
 sg13g2_and2_1 _08939_ (.A(net161),
    .B(_03434_),
    .X(_00404_));
 sg13g2_mux2_1 _08940_ (.A0(\shift_storage.storage [1272]),
    .A1(\shift_storage.storage [1271]),
    .S(net160),
    .X(_03435_));
 sg13g2_and2_1 _08941_ (.A(net161),
    .B(_03435_),
    .X(_00405_));
 sg13g2_mux2_1 _08942_ (.A0(\shift_storage.storage [1273]),
    .A1(\shift_storage.storage [1272]),
    .S(net160),
    .X(_03436_));
 sg13g2_and2_1 _08943_ (.A(net161),
    .B(_03436_),
    .X(_00406_));
 sg13g2_mux2_1 _08944_ (.A0(\shift_storage.storage [1274]),
    .A1(\shift_storage.storage [1273]),
    .S(net160),
    .X(_03437_));
 sg13g2_and2_1 _08945_ (.A(_03427_),
    .B(_03437_),
    .X(_00407_));
 sg13g2_mux2_1 _08946_ (.A0(\shift_storage.storage [1275]),
    .A1(\shift_storage.storage [1274]),
    .S(net160),
    .X(_03438_));
 sg13g2_and2_1 _08947_ (.A(_03427_),
    .B(_03438_),
    .X(_00408_));
 sg13g2_buf_1 _08948_ (.A(net365),
    .X(_03439_));
 sg13g2_mux2_1 _08949_ (.A0(\shift_storage.storage [1276]),
    .A1(\shift_storage.storage [1275]),
    .S(_03432_),
    .X(_03440_));
 sg13g2_and2_1 _08950_ (.A(net159),
    .B(_03440_),
    .X(_00409_));
 sg13g2_mux2_1 _08951_ (.A0(\shift_storage.storage [1277]),
    .A1(\shift_storage.storage [1276]),
    .S(_03432_),
    .X(_03441_));
 sg13g2_and2_1 _08952_ (.A(net159),
    .B(_03441_),
    .X(_00410_));
 sg13g2_mux2_1 _08953_ (.A0(\shift_storage.storage [1278]),
    .A1(\shift_storage.storage [1277]),
    .S(net160),
    .X(_03442_));
 sg13g2_and2_1 _08954_ (.A(_03439_),
    .B(_03442_),
    .X(_00411_));
 sg13g2_mux2_1 _08955_ (.A0(\shift_storage.storage [1279]),
    .A1(\shift_storage.storage [1278]),
    .S(net160),
    .X(_03443_));
 sg13g2_and2_1 _08956_ (.A(_03439_),
    .B(_03443_),
    .X(_00412_));
 sg13g2_buf_1 _08957_ (.A(net366),
    .X(_03444_));
 sg13g2_mux2_1 _08958_ (.A0(\shift_storage.storage [127]),
    .A1(\shift_storage.storage [126]),
    .S(net158),
    .X(_03445_));
 sg13g2_and2_1 _08959_ (.A(net159),
    .B(_03445_),
    .X(_00413_));
 sg13g2_mux2_1 _08960_ (.A0(\shift_storage.storage [1280]),
    .A1(\shift_storage.storage [1279]),
    .S(net158),
    .X(_03446_));
 sg13g2_and2_1 _08961_ (.A(net159),
    .B(_03446_),
    .X(_00414_));
 sg13g2_mux2_1 _08962_ (.A0(\shift_storage.storage [1281]),
    .A1(\shift_storage.storage [1280]),
    .S(net158),
    .X(_03447_));
 sg13g2_and2_1 _08963_ (.A(net159),
    .B(_03447_),
    .X(_00415_));
 sg13g2_mux2_1 _08964_ (.A0(\shift_storage.storage [1282]),
    .A1(\shift_storage.storage [1281]),
    .S(net158),
    .X(_03448_));
 sg13g2_and2_1 _08965_ (.A(net159),
    .B(_03448_),
    .X(_00416_));
 sg13g2_mux2_1 _08966_ (.A0(\shift_storage.storage [1283]),
    .A1(\shift_storage.storage [1282]),
    .S(_03444_),
    .X(_03449_));
 sg13g2_and2_1 _08967_ (.A(net159),
    .B(_03449_),
    .X(_00417_));
 sg13g2_mux2_1 _08968_ (.A0(\shift_storage.storage [1284]),
    .A1(\shift_storage.storage [1283]),
    .S(_03444_),
    .X(_03450_));
 sg13g2_and2_1 _08969_ (.A(net159),
    .B(_03450_),
    .X(_00418_));
 sg13g2_buf_1 _08970_ (.A(net365),
    .X(_03451_));
 sg13g2_mux2_1 _08971_ (.A0(\shift_storage.storage [1285]),
    .A1(\shift_storage.storage [1284]),
    .S(net158),
    .X(_03452_));
 sg13g2_and2_1 _08972_ (.A(net157),
    .B(_03452_),
    .X(_00419_));
 sg13g2_mux2_1 _08973_ (.A0(\shift_storage.storage [1286]),
    .A1(\shift_storage.storage [1285]),
    .S(net158),
    .X(_03453_));
 sg13g2_and2_1 _08974_ (.A(net157),
    .B(_03453_),
    .X(_00420_));
 sg13g2_mux2_1 _08975_ (.A0(\shift_storage.storage [1287]),
    .A1(\shift_storage.storage [1286]),
    .S(net158),
    .X(_03454_));
 sg13g2_and2_1 _08976_ (.A(net157),
    .B(_03454_),
    .X(_00421_));
 sg13g2_mux2_1 _08977_ (.A0(\shift_storage.storage [1288]),
    .A1(\shift_storage.storage [1287]),
    .S(net158),
    .X(_03455_));
 sg13g2_and2_1 _08978_ (.A(net157),
    .B(_03455_),
    .X(_00422_));
 sg13g2_buf_1 _08979_ (.A(net366),
    .X(_03456_));
 sg13g2_mux2_1 _08980_ (.A0(\shift_storage.storage [1289]),
    .A1(\shift_storage.storage [1288]),
    .S(net156),
    .X(_03457_));
 sg13g2_and2_1 _08981_ (.A(net157),
    .B(_03457_),
    .X(_00423_));
 sg13g2_mux2_1 _08982_ (.A0(\shift_storage.storage [128]),
    .A1(\shift_storage.storage [127]),
    .S(net156),
    .X(_03458_));
 sg13g2_and2_1 _08983_ (.A(net157),
    .B(_03458_),
    .X(_00424_));
 sg13g2_mux2_1 _08984_ (.A0(\shift_storage.storage [1290]),
    .A1(\shift_storage.storage [1289]),
    .S(net156),
    .X(_03459_));
 sg13g2_and2_1 _08985_ (.A(net157),
    .B(_03459_),
    .X(_00425_));
 sg13g2_mux2_1 _08986_ (.A0(\shift_storage.storage [1291]),
    .A1(\shift_storage.storage [1290]),
    .S(net156),
    .X(_03460_));
 sg13g2_and2_1 _08987_ (.A(net157),
    .B(_03460_),
    .X(_00426_));
 sg13g2_mux2_1 _08988_ (.A0(\shift_storage.storage [1292]),
    .A1(\shift_storage.storage [1291]),
    .S(net156),
    .X(_03461_));
 sg13g2_and2_1 _08989_ (.A(_03451_),
    .B(_03461_),
    .X(_00427_));
 sg13g2_mux2_1 _08990_ (.A0(\shift_storage.storage [1293]),
    .A1(\shift_storage.storage [1292]),
    .S(net156),
    .X(_03462_));
 sg13g2_and2_1 _08991_ (.A(_03451_),
    .B(_03462_),
    .X(_00428_));
 sg13g2_buf_1 _08992_ (.A(net365),
    .X(_03463_));
 sg13g2_mux2_1 _08993_ (.A0(\shift_storage.storage [1294]),
    .A1(\shift_storage.storage [1293]),
    .S(net156),
    .X(_03464_));
 sg13g2_and2_1 _08994_ (.A(net155),
    .B(_03464_),
    .X(_00429_));
 sg13g2_mux2_1 _08995_ (.A0(\shift_storage.storage [1295]),
    .A1(\shift_storage.storage [1294]),
    .S(net156),
    .X(_03465_));
 sg13g2_and2_1 _08996_ (.A(net155),
    .B(_03465_),
    .X(_00430_));
 sg13g2_mux2_1 _08997_ (.A0(\shift_storage.storage [1296]),
    .A1(\shift_storage.storage [1295]),
    .S(_03456_),
    .X(_03466_));
 sg13g2_and2_1 _08998_ (.A(_03463_),
    .B(_03466_),
    .X(_00431_));
 sg13g2_mux2_1 _08999_ (.A0(\shift_storage.storage [1297]),
    .A1(\shift_storage.storage [1296]),
    .S(_03456_),
    .X(_03467_));
 sg13g2_and2_1 _09000_ (.A(net155),
    .B(_03467_),
    .X(_00432_));
 sg13g2_buf_1 _09001_ (.A(net366),
    .X(_03468_));
 sg13g2_mux2_1 _09002_ (.A0(\shift_storage.storage [1298]),
    .A1(\shift_storage.storage [1297]),
    .S(net154),
    .X(_03469_));
 sg13g2_and2_1 _09003_ (.A(net155),
    .B(_03469_),
    .X(_00433_));
 sg13g2_mux2_1 _09004_ (.A0(\shift_storage.storage [1299]),
    .A1(\shift_storage.storage [1298]),
    .S(net154),
    .X(_03470_));
 sg13g2_and2_1 _09005_ (.A(net155),
    .B(_03470_),
    .X(_00434_));
 sg13g2_mux2_1 _09006_ (.A0(\shift_storage.storage [129]),
    .A1(\shift_storage.storage [128]),
    .S(net154),
    .X(_03471_));
 sg13g2_and2_1 _09007_ (.A(_03463_),
    .B(_03471_),
    .X(_00435_));
 sg13g2_mux2_1 _09008_ (.A0(\shift_storage.storage [12]),
    .A1(\shift_storage.storage [11]),
    .S(net154),
    .X(_03472_));
 sg13g2_and2_1 _09009_ (.A(net155),
    .B(_03472_),
    .X(_00436_));
 sg13g2_mux2_1 _09010_ (.A0(\shift_storage.storage [1300]),
    .A1(\shift_storage.storage [1299]),
    .S(net154),
    .X(_03473_));
 sg13g2_and2_1 _09011_ (.A(net155),
    .B(_03473_),
    .X(_00437_));
 sg13g2_mux2_1 _09012_ (.A0(\shift_storage.storage [1301]),
    .A1(\shift_storage.storage [1300]),
    .S(net154),
    .X(_03474_));
 sg13g2_and2_1 _09013_ (.A(net155),
    .B(_03474_),
    .X(_00438_));
 sg13g2_buf_1 _09014_ (.A(net365),
    .X(_03475_));
 sg13g2_mux2_1 _09015_ (.A0(\shift_storage.storage [1302]),
    .A1(\shift_storage.storage [1301]),
    .S(net154),
    .X(_03476_));
 sg13g2_and2_1 _09016_ (.A(net153),
    .B(_03476_),
    .X(_00439_));
 sg13g2_mux2_1 _09017_ (.A0(\shift_storage.storage [1303]),
    .A1(\shift_storage.storage [1302]),
    .S(net154),
    .X(_03477_));
 sg13g2_and2_1 _09018_ (.A(net153),
    .B(_03477_),
    .X(_00440_));
 sg13g2_mux2_1 _09019_ (.A0(\shift_storage.storage [1304]),
    .A1(\shift_storage.storage [1303]),
    .S(_03468_),
    .X(_03478_));
 sg13g2_and2_1 _09020_ (.A(net153),
    .B(_03478_),
    .X(_00441_));
 sg13g2_mux2_1 _09021_ (.A0(\shift_storage.storage [1305]),
    .A1(\shift_storage.storage [1304]),
    .S(_03468_),
    .X(_03479_));
 sg13g2_and2_1 _09022_ (.A(net153),
    .B(_03479_),
    .X(_00442_));
 sg13g2_buf_1 _09023_ (.A(net366),
    .X(_03480_));
 sg13g2_mux2_1 _09024_ (.A0(\shift_storage.storage [1306]),
    .A1(\shift_storage.storage [1305]),
    .S(net152),
    .X(_03481_));
 sg13g2_and2_1 _09025_ (.A(net153),
    .B(_03481_),
    .X(_00443_));
 sg13g2_mux2_1 _09026_ (.A0(\shift_storage.storage [1307]),
    .A1(\shift_storage.storage [1306]),
    .S(net152),
    .X(_03482_));
 sg13g2_and2_1 _09027_ (.A(net153),
    .B(_03482_),
    .X(_00444_));
 sg13g2_mux2_1 _09028_ (.A0(\shift_storage.storage [1308]),
    .A1(\shift_storage.storage [1307]),
    .S(net152),
    .X(_03483_));
 sg13g2_and2_1 _09029_ (.A(net153),
    .B(_03483_),
    .X(_00445_));
 sg13g2_mux2_1 _09030_ (.A0(\shift_storage.storage [1309]),
    .A1(\shift_storage.storage [1308]),
    .S(_03480_),
    .X(_03484_));
 sg13g2_and2_1 _09031_ (.A(net153),
    .B(_03484_),
    .X(_00446_));
 sg13g2_mux2_1 _09032_ (.A0(\shift_storage.storage [130]),
    .A1(\shift_storage.storage [129]),
    .S(_03480_),
    .X(_03485_));
 sg13g2_and2_1 _09033_ (.A(_03475_),
    .B(_03485_),
    .X(_00447_));
 sg13g2_mux2_1 _09034_ (.A0(\shift_storage.storage [1310]),
    .A1(\shift_storage.storage [1309]),
    .S(net152),
    .X(_03486_));
 sg13g2_and2_1 _09035_ (.A(_03475_),
    .B(_03486_),
    .X(_00448_));
 sg13g2_buf_1 _09036_ (.A(net365),
    .X(_03487_));
 sg13g2_mux2_1 _09037_ (.A0(\shift_storage.storage [1311]),
    .A1(\shift_storage.storage [1310]),
    .S(net152),
    .X(_03488_));
 sg13g2_and2_1 _09038_ (.A(net151),
    .B(_03488_),
    .X(_00449_));
 sg13g2_mux2_1 _09039_ (.A0(\shift_storage.storage [1312]),
    .A1(\shift_storage.storage [1311]),
    .S(net152),
    .X(_03489_));
 sg13g2_and2_1 _09040_ (.A(net151),
    .B(_03489_),
    .X(_00450_));
 sg13g2_mux2_1 _09041_ (.A0(\shift_storage.storage [1313]),
    .A1(\shift_storage.storage [1312]),
    .S(net152),
    .X(_03490_));
 sg13g2_and2_1 _09042_ (.A(net151),
    .B(_03490_),
    .X(_00451_));
 sg13g2_mux2_1 _09043_ (.A0(\shift_storage.storage [1314]),
    .A1(\shift_storage.storage [1313]),
    .S(net152),
    .X(_03491_));
 sg13g2_and2_1 _09044_ (.A(net151),
    .B(_03491_),
    .X(_00452_));
 sg13g2_buf_1 _09045_ (.A(net366),
    .X(_03492_));
 sg13g2_mux2_1 _09046_ (.A0(\shift_storage.storage [1315]),
    .A1(\shift_storage.storage [1314]),
    .S(net150),
    .X(_03493_));
 sg13g2_and2_1 _09047_ (.A(net151),
    .B(_03493_),
    .X(_00453_));
 sg13g2_mux2_1 _09048_ (.A0(\shift_storage.storage [1316]),
    .A1(\shift_storage.storage [1315]),
    .S(net150),
    .X(_03494_));
 sg13g2_and2_1 _09049_ (.A(net151),
    .B(_03494_),
    .X(_00454_));
 sg13g2_mux2_1 _09050_ (.A0(\shift_storage.storage [1317]),
    .A1(\shift_storage.storage [1316]),
    .S(net150),
    .X(_03495_));
 sg13g2_and2_1 _09051_ (.A(net151),
    .B(_03495_),
    .X(_00455_));
 sg13g2_mux2_1 _09052_ (.A0(\shift_storage.storage [1318]),
    .A1(\shift_storage.storage [1317]),
    .S(net150),
    .X(_03496_));
 sg13g2_and2_1 _09053_ (.A(net151),
    .B(_03496_),
    .X(_00456_));
 sg13g2_mux2_1 _09054_ (.A0(\shift_storage.storage [1319]),
    .A1(\shift_storage.storage [1318]),
    .S(net150),
    .X(_03497_));
 sg13g2_and2_1 _09055_ (.A(_03487_),
    .B(_03497_),
    .X(_00457_));
 sg13g2_mux2_1 _09056_ (.A0(\shift_storage.storage [131]),
    .A1(\shift_storage.storage [130]),
    .S(net150),
    .X(_03498_));
 sg13g2_and2_1 _09057_ (.A(_03487_),
    .B(_03498_),
    .X(_00458_));
 sg13g2_buf_1 _09058_ (.A(net365),
    .X(_03499_));
 sg13g2_mux2_1 _09059_ (.A0(\shift_storage.storage [1320]),
    .A1(\shift_storage.storage [1319]),
    .S(net150),
    .X(_03500_));
 sg13g2_and2_1 _09060_ (.A(net149),
    .B(_03500_),
    .X(_00459_));
 sg13g2_mux2_1 _09061_ (.A0(\shift_storage.storage [1321]),
    .A1(\shift_storage.storage [1320]),
    .S(net150),
    .X(_03501_));
 sg13g2_and2_1 _09062_ (.A(net149),
    .B(_03501_),
    .X(_00460_));
 sg13g2_mux2_1 _09063_ (.A0(\shift_storage.storage [1322]),
    .A1(\shift_storage.storage [1321]),
    .S(_03492_),
    .X(_03502_));
 sg13g2_and2_1 _09064_ (.A(net149),
    .B(_03502_),
    .X(_00461_));
 sg13g2_mux2_1 _09065_ (.A0(\shift_storage.storage [1323]),
    .A1(\shift_storage.storage [1322]),
    .S(_03492_),
    .X(_03503_));
 sg13g2_and2_1 _09066_ (.A(net149),
    .B(_03503_),
    .X(_00462_));
 sg13g2_buf_1 _09067_ (.A(net366),
    .X(_03504_));
 sg13g2_mux2_1 _09068_ (.A0(\shift_storage.storage [1324]),
    .A1(\shift_storage.storage [1323]),
    .S(net148),
    .X(_03505_));
 sg13g2_and2_1 _09069_ (.A(net149),
    .B(_03505_),
    .X(_00463_));
 sg13g2_mux2_1 _09070_ (.A0(\shift_storage.storage [1325]),
    .A1(\shift_storage.storage [1324]),
    .S(net148),
    .X(_03506_));
 sg13g2_and2_1 _09071_ (.A(net149),
    .B(_03506_),
    .X(_00464_));
 sg13g2_mux2_1 _09072_ (.A0(\shift_storage.storage [1326]),
    .A1(\shift_storage.storage [1325]),
    .S(net148),
    .X(_03507_));
 sg13g2_and2_1 _09073_ (.A(_03499_),
    .B(_03507_),
    .X(_00465_));
 sg13g2_mux2_1 _09074_ (.A0(\shift_storage.storage [1327]),
    .A1(\shift_storage.storage [1326]),
    .S(net148),
    .X(_03508_));
 sg13g2_and2_1 _09075_ (.A(_03499_),
    .B(_03508_),
    .X(_00466_));
 sg13g2_mux2_1 _09076_ (.A0(\shift_storage.storage [1328]),
    .A1(\shift_storage.storage [1327]),
    .S(net148),
    .X(_03509_));
 sg13g2_and2_1 _09077_ (.A(net149),
    .B(_03509_),
    .X(_00467_));
 sg13g2_mux2_1 _09078_ (.A0(\shift_storage.storage [1329]),
    .A1(\shift_storage.storage [1328]),
    .S(net148),
    .X(_03510_));
 sg13g2_and2_1 _09079_ (.A(net149),
    .B(_03510_),
    .X(_00468_));
 sg13g2_buf_1 _09080_ (.A(net365),
    .X(_03511_));
 sg13g2_mux2_1 _09081_ (.A0(\shift_storage.storage [132]),
    .A1(\shift_storage.storage [131]),
    .S(net148),
    .X(_03512_));
 sg13g2_and2_1 _09082_ (.A(net147),
    .B(_03512_),
    .X(_00469_));
 sg13g2_mux2_1 _09083_ (.A0(\shift_storage.storage [1330]),
    .A1(\shift_storage.storage [1329]),
    .S(net148),
    .X(_03513_));
 sg13g2_and2_1 _09084_ (.A(net147),
    .B(_03513_),
    .X(_00470_));
 sg13g2_mux2_1 _09085_ (.A0(\shift_storage.storage [1331]),
    .A1(\shift_storage.storage [1330]),
    .S(_03504_),
    .X(_03514_));
 sg13g2_and2_1 _09086_ (.A(net147),
    .B(_03514_),
    .X(_00471_));
 sg13g2_mux2_1 _09087_ (.A0(\shift_storage.storage [1332]),
    .A1(\shift_storage.storage [1331]),
    .S(_03504_),
    .X(_03515_));
 sg13g2_and2_1 _09088_ (.A(net147),
    .B(_03515_),
    .X(_00472_));
 sg13g2_buf_1 _09089_ (.A(_03418_),
    .X(_03516_));
 sg13g2_mux2_1 _09090_ (.A0(\shift_storage.storage [1333]),
    .A1(\shift_storage.storage [1332]),
    .S(net146),
    .X(_03517_));
 sg13g2_and2_1 _09091_ (.A(net147),
    .B(_03517_),
    .X(_00473_));
 sg13g2_mux2_1 _09092_ (.A0(\shift_storage.storage [1334]),
    .A1(\shift_storage.storage [1333]),
    .S(net146),
    .X(_03518_));
 sg13g2_and2_1 _09093_ (.A(net147),
    .B(_03518_),
    .X(_00474_));
 sg13g2_mux2_1 _09094_ (.A0(\shift_storage.storage [1335]),
    .A1(\shift_storage.storage [1334]),
    .S(net146),
    .X(_03519_));
 sg13g2_and2_1 _09095_ (.A(net147),
    .B(_03519_),
    .X(_00475_));
 sg13g2_mux2_1 _09096_ (.A0(\shift_storage.storage [1336]),
    .A1(\shift_storage.storage [1335]),
    .S(net146),
    .X(_03520_));
 sg13g2_and2_1 _09097_ (.A(net147),
    .B(_03520_),
    .X(_00476_));
 sg13g2_mux2_1 _09098_ (.A0(\shift_storage.storage [1337]),
    .A1(\shift_storage.storage [1336]),
    .S(net146),
    .X(_03521_));
 sg13g2_and2_1 _09099_ (.A(_03511_),
    .B(_03521_),
    .X(_00477_));
 sg13g2_mux2_1 _09100_ (.A0(\shift_storage.storage [1338]),
    .A1(\shift_storage.storage [1337]),
    .S(net146),
    .X(_03522_));
 sg13g2_and2_1 _09101_ (.A(_03511_),
    .B(_03522_),
    .X(_00478_));
 sg13g2_buf_1 _09102_ (.A(_03426_),
    .X(_03523_));
 sg13g2_mux2_1 _09103_ (.A0(\shift_storage.storage [1339]),
    .A1(\shift_storage.storage [1338]),
    .S(net146),
    .X(_03524_));
 sg13g2_and2_1 _09104_ (.A(net145),
    .B(_03524_),
    .X(_00479_));
 sg13g2_mux2_1 _09105_ (.A0(\shift_storage.storage [133]),
    .A1(\shift_storage.storage [132]),
    .S(net146),
    .X(_03525_));
 sg13g2_and2_1 _09106_ (.A(net145),
    .B(_03525_),
    .X(_00480_));
 sg13g2_mux2_1 _09107_ (.A0(\shift_storage.storage [1340]),
    .A1(\shift_storage.storage [1339]),
    .S(_03516_),
    .X(_03526_));
 sg13g2_and2_1 _09108_ (.A(net145),
    .B(_03526_),
    .X(_00481_));
 sg13g2_mux2_1 _09109_ (.A0(\shift_storage.storage [1341]),
    .A1(\shift_storage.storage [1340]),
    .S(_03516_),
    .X(_03527_));
 sg13g2_and2_1 _09110_ (.A(net145),
    .B(_03527_),
    .X(_00482_));
 sg13g2_buf_1 _09111_ (.A(_03418_),
    .X(_03528_));
 sg13g2_mux2_1 _09112_ (.A0(\shift_storage.storage [1342]),
    .A1(\shift_storage.storage [1341]),
    .S(net144),
    .X(_03529_));
 sg13g2_and2_1 _09113_ (.A(net145),
    .B(_03529_),
    .X(_00483_));
 sg13g2_mux2_1 _09114_ (.A0(\shift_storage.storage [1343]),
    .A1(\shift_storage.storage [1342]),
    .S(net144),
    .X(_03530_));
 sg13g2_and2_1 _09115_ (.A(_03523_),
    .B(_03530_),
    .X(_00484_));
 sg13g2_mux2_1 _09116_ (.A0(\shift_storage.storage [1344]),
    .A1(\shift_storage.storage [1343]),
    .S(_03528_),
    .X(_03531_));
 sg13g2_and2_1 _09117_ (.A(_03523_),
    .B(_03531_),
    .X(_00485_));
 sg13g2_mux2_1 _09118_ (.A0(\shift_storage.storage [1345]),
    .A1(\shift_storage.storage [1344]),
    .S(_03528_),
    .X(_03532_));
 sg13g2_and2_1 _09119_ (.A(net145),
    .B(_03532_),
    .X(_00486_));
 sg13g2_mux2_1 _09120_ (.A0(\shift_storage.storage [1346]),
    .A1(\shift_storage.storage [1345]),
    .S(net144),
    .X(_03533_));
 sg13g2_and2_1 _09121_ (.A(net145),
    .B(_03533_),
    .X(_00487_));
 sg13g2_mux2_1 _09122_ (.A0(\shift_storage.storage [1347]),
    .A1(\shift_storage.storage [1346]),
    .S(net144),
    .X(_03534_));
 sg13g2_and2_1 _09123_ (.A(net145),
    .B(_03534_),
    .X(_00488_));
 sg13g2_buf_1 _09124_ (.A(_03426_),
    .X(_03535_));
 sg13g2_mux2_1 _09125_ (.A0(\shift_storage.storage [1348]),
    .A1(\shift_storage.storage [1347]),
    .S(net144),
    .X(_03536_));
 sg13g2_and2_1 _09126_ (.A(net143),
    .B(_03536_),
    .X(_00489_));
 sg13g2_mux2_1 _09127_ (.A0(\shift_storage.storage [1349]),
    .A1(\shift_storage.storage [1348]),
    .S(net144),
    .X(_03537_));
 sg13g2_and2_1 _09128_ (.A(net143),
    .B(_03537_),
    .X(_00490_));
 sg13g2_mux2_1 _09129_ (.A0(\shift_storage.storage [134]),
    .A1(\shift_storage.storage [133]),
    .S(net144),
    .X(_03538_));
 sg13g2_and2_1 _09130_ (.A(net143),
    .B(_03538_),
    .X(_00491_));
 sg13g2_mux2_1 _09131_ (.A0(\shift_storage.storage [1350]),
    .A1(\shift_storage.storage [1349]),
    .S(net144),
    .X(_03539_));
 sg13g2_and2_1 _09132_ (.A(net143),
    .B(_03539_),
    .X(_00492_));
 sg13g2_buf_1 _09133_ (.A(net410),
    .X(_03540_));
 sg13g2_buf_1 _09134_ (.A(net364),
    .X(_03541_));
 sg13g2_mux2_1 _09135_ (.A0(\shift_storage.storage [1351]),
    .A1(\shift_storage.storage [1350]),
    .S(net142),
    .X(_03542_));
 sg13g2_and2_1 _09136_ (.A(net143),
    .B(_03542_),
    .X(_00493_));
 sg13g2_mux2_1 _09137_ (.A0(\shift_storage.storage [1352]),
    .A1(\shift_storage.storage [1351]),
    .S(net142),
    .X(_03543_));
 sg13g2_and2_1 _09138_ (.A(net143),
    .B(_03543_),
    .X(_00494_));
 sg13g2_mux2_1 _09139_ (.A0(\shift_storage.storage [1353]),
    .A1(\shift_storage.storage [1352]),
    .S(net142),
    .X(_03544_));
 sg13g2_and2_1 _09140_ (.A(net143),
    .B(_03544_),
    .X(_00495_));
 sg13g2_mux2_1 _09141_ (.A0(\shift_storage.storage [1354]),
    .A1(\shift_storage.storage [1353]),
    .S(net142),
    .X(_03545_));
 sg13g2_and2_1 _09142_ (.A(net143),
    .B(_03545_),
    .X(_00496_));
 sg13g2_mux2_1 _09143_ (.A0(\shift_storage.storage [1355]),
    .A1(\shift_storage.storage [1354]),
    .S(_03541_),
    .X(_03546_));
 sg13g2_and2_1 _09144_ (.A(_03535_),
    .B(_03546_),
    .X(_00497_));
 sg13g2_mux2_1 _09145_ (.A0(\shift_storage.storage [1356]),
    .A1(\shift_storage.storage [1355]),
    .S(_03541_),
    .X(_03547_));
 sg13g2_and2_1 _09146_ (.A(_03535_),
    .B(_03547_),
    .X(_00498_));
 sg13g2_buf_1 _09147_ (.A(net411),
    .X(_03548_));
 sg13g2_buf_1 _09148_ (.A(net363),
    .X(_03549_));
 sg13g2_mux2_1 _09149_ (.A0(\shift_storage.storage [1357]),
    .A1(\shift_storage.storage [1356]),
    .S(net142),
    .X(_03550_));
 sg13g2_and2_1 _09150_ (.A(net141),
    .B(_03550_),
    .X(_00499_));
 sg13g2_mux2_1 _09151_ (.A0(\shift_storage.storage [1358]),
    .A1(\shift_storage.storage [1357]),
    .S(net142),
    .X(_03551_));
 sg13g2_and2_1 _09152_ (.A(net141),
    .B(_03551_),
    .X(_00500_));
 sg13g2_mux2_1 _09153_ (.A0(\shift_storage.storage [1359]),
    .A1(\shift_storage.storage [1358]),
    .S(net142),
    .X(_03552_));
 sg13g2_and2_1 _09154_ (.A(net141),
    .B(_03552_),
    .X(_00501_));
 sg13g2_mux2_1 _09155_ (.A0(\shift_storage.storage [135]),
    .A1(\shift_storage.storage [134]),
    .S(net142),
    .X(_03553_));
 sg13g2_and2_1 _09156_ (.A(net141),
    .B(_03553_),
    .X(_00502_));
 sg13g2_buf_1 _09157_ (.A(net364),
    .X(_03554_));
 sg13g2_mux2_1 _09158_ (.A0(\shift_storage.storage [1360]),
    .A1(\shift_storage.storage [1359]),
    .S(net140),
    .X(_03555_));
 sg13g2_and2_1 _09159_ (.A(_03549_),
    .B(_03555_),
    .X(_00503_));
 sg13g2_mux2_1 _09160_ (.A0(\shift_storage.storage [1361]),
    .A1(\shift_storage.storage [1360]),
    .S(net140),
    .X(_03556_));
 sg13g2_and2_1 _09161_ (.A(_03549_),
    .B(_03556_),
    .X(_00504_));
 sg13g2_mux2_1 _09162_ (.A0(\shift_storage.storage [1362]),
    .A1(\shift_storage.storage [1361]),
    .S(net140),
    .X(_03557_));
 sg13g2_and2_1 _09163_ (.A(net141),
    .B(_03557_),
    .X(_00505_));
 sg13g2_mux2_1 _09164_ (.A0(\shift_storage.storage [1363]),
    .A1(\shift_storage.storage [1362]),
    .S(net140),
    .X(_03558_));
 sg13g2_and2_1 _09165_ (.A(net141),
    .B(_03558_),
    .X(_00506_));
 sg13g2_mux2_1 _09166_ (.A0(\shift_storage.storage [1364]),
    .A1(\shift_storage.storage [1363]),
    .S(_03554_),
    .X(_03559_));
 sg13g2_and2_1 _09167_ (.A(net141),
    .B(_03559_),
    .X(_00507_));
 sg13g2_mux2_1 _09168_ (.A0(\shift_storage.storage [1365]),
    .A1(\shift_storage.storage [1364]),
    .S(_03554_),
    .X(_03560_));
 sg13g2_and2_1 _09169_ (.A(net141),
    .B(_03560_),
    .X(_00508_));
 sg13g2_buf_1 _09170_ (.A(net363),
    .X(_03561_));
 sg13g2_mux2_1 _09171_ (.A0(\shift_storage.storage [1366]),
    .A1(\shift_storage.storage [1365]),
    .S(net140),
    .X(_03562_));
 sg13g2_and2_1 _09172_ (.A(net139),
    .B(_03562_),
    .X(_00509_));
 sg13g2_mux2_1 _09173_ (.A0(\shift_storage.storage [1367]),
    .A1(\shift_storage.storage [1366]),
    .S(net140),
    .X(_03563_));
 sg13g2_and2_1 _09174_ (.A(net139),
    .B(_03563_),
    .X(_00510_));
 sg13g2_mux2_1 _09175_ (.A0(\shift_storage.storage [1368]),
    .A1(\shift_storage.storage [1367]),
    .S(net140),
    .X(_03564_));
 sg13g2_and2_1 _09176_ (.A(net139),
    .B(_03564_),
    .X(_00511_));
 sg13g2_mux2_1 _09177_ (.A0(\shift_storage.storage [1369]),
    .A1(\shift_storage.storage [1368]),
    .S(net140),
    .X(_03565_));
 sg13g2_and2_1 _09178_ (.A(net139),
    .B(_03565_),
    .X(_00512_));
 sg13g2_buf_1 _09179_ (.A(net364),
    .X(_03566_));
 sg13g2_mux2_1 _09180_ (.A0(\shift_storage.storage [136]),
    .A1(\shift_storage.storage [135]),
    .S(net138),
    .X(_03567_));
 sg13g2_and2_1 _09181_ (.A(_03561_),
    .B(_03567_),
    .X(_00513_));
 sg13g2_mux2_1 _09182_ (.A0(\shift_storage.storage [1370]),
    .A1(\shift_storage.storage [1369]),
    .S(net138),
    .X(_03568_));
 sg13g2_and2_1 _09183_ (.A(net139),
    .B(_03568_),
    .X(_00514_));
 sg13g2_mux2_1 _09184_ (.A0(\shift_storage.storage [1371]),
    .A1(\shift_storage.storage [1370]),
    .S(net138),
    .X(_03569_));
 sg13g2_and2_1 _09185_ (.A(net139),
    .B(_03569_),
    .X(_00515_));
 sg13g2_mux2_1 _09186_ (.A0(\shift_storage.storage [1372]),
    .A1(\shift_storage.storage [1371]),
    .S(net138),
    .X(_03570_));
 sg13g2_and2_1 _09187_ (.A(net139),
    .B(_03570_),
    .X(_00516_));
 sg13g2_mux2_1 _09188_ (.A0(\shift_storage.storage [1373]),
    .A1(\shift_storage.storage [1372]),
    .S(net138),
    .X(_03571_));
 sg13g2_and2_1 _09189_ (.A(net139),
    .B(_03571_),
    .X(_00517_));
 sg13g2_mux2_1 _09190_ (.A0(\shift_storage.storage [1374]),
    .A1(\shift_storage.storage [1373]),
    .S(net138),
    .X(_03572_));
 sg13g2_and2_1 _09191_ (.A(_03561_),
    .B(_03572_),
    .X(_00518_));
 sg13g2_buf_1 _09192_ (.A(net363),
    .X(_03573_));
 sg13g2_mux2_1 _09193_ (.A0(\shift_storage.storage [1375]),
    .A1(\shift_storage.storage [1374]),
    .S(net138),
    .X(_03574_));
 sg13g2_and2_1 _09194_ (.A(net137),
    .B(_03574_),
    .X(_00519_));
 sg13g2_mux2_1 _09195_ (.A0(\shift_storage.storage [1376]),
    .A1(\shift_storage.storage [1375]),
    .S(net138),
    .X(_03575_));
 sg13g2_and2_1 _09196_ (.A(net137),
    .B(_03575_),
    .X(_00520_));
 sg13g2_mux2_1 _09197_ (.A0(\shift_storage.storage [1377]),
    .A1(\shift_storage.storage [1376]),
    .S(_03566_),
    .X(_03576_));
 sg13g2_and2_1 _09198_ (.A(net137),
    .B(_03576_),
    .X(_00521_));
 sg13g2_mux2_1 _09199_ (.A0(\shift_storage.storage [1378]),
    .A1(\shift_storage.storage [1377]),
    .S(_03566_),
    .X(_03577_));
 sg13g2_and2_1 _09200_ (.A(net137),
    .B(_03577_),
    .X(_00522_));
 sg13g2_buf_1 _09201_ (.A(net364),
    .X(_03578_));
 sg13g2_mux2_1 _09202_ (.A0(\shift_storage.storage [1379]),
    .A1(\shift_storage.storage [1378]),
    .S(net136),
    .X(_03579_));
 sg13g2_and2_1 _09203_ (.A(net137),
    .B(_03579_),
    .X(_00523_));
 sg13g2_mux2_1 _09204_ (.A0(\shift_storage.storage [137]),
    .A1(\shift_storage.storage [136]),
    .S(net136),
    .X(_03580_));
 sg13g2_and2_1 _09205_ (.A(net137),
    .B(_03580_),
    .X(_00524_));
 sg13g2_mux2_1 _09206_ (.A0(\shift_storage.storage [1380]),
    .A1(\shift_storage.storage [1379]),
    .S(net136),
    .X(_03581_));
 sg13g2_and2_1 _09207_ (.A(net137),
    .B(_03581_),
    .X(_00525_));
 sg13g2_mux2_1 _09208_ (.A0(\shift_storage.storage [1381]),
    .A1(\shift_storage.storage [1380]),
    .S(net136),
    .X(_03582_));
 sg13g2_and2_1 _09209_ (.A(net137),
    .B(_03582_),
    .X(_00526_));
 sg13g2_mux2_1 _09210_ (.A0(\shift_storage.storage [1382]),
    .A1(\shift_storage.storage [1381]),
    .S(net136),
    .X(_03583_));
 sg13g2_and2_1 _09211_ (.A(_03573_),
    .B(_03583_),
    .X(_00527_));
 sg13g2_mux2_1 _09212_ (.A0(\shift_storage.storage [1383]),
    .A1(\shift_storage.storage [1382]),
    .S(net136),
    .X(_03584_));
 sg13g2_and2_1 _09213_ (.A(_03573_),
    .B(_03584_),
    .X(_00528_));
 sg13g2_buf_1 _09214_ (.A(_03548_),
    .X(_03585_));
 sg13g2_mux2_1 _09215_ (.A0(\shift_storage.storage [1384]),
    .A1(\shift_storage.storage [1383]),
    .S(net136),
    .X(_03586_));
 sg13g2_and2_1 _09216_ (.A(net135),
    .B(_03586_),
    .X(_00529_));
 sg13g2_mux2_1 _09217_ (.A0(\shift_storage.storage [1385]),
    .A1(\shift_storage.storage [1384]),
    .S(net136),
    .X(_03587_));
 sg13g2_and2_1 _09218_ (.A(net135),
    .B(_03587_),
    .X(_00530_));
 sg13g2_mux2_1 _09219_ (.A0(\shift_storage.storage [1386]),
    .A1(\shift_storage.storage [1385]),
    .S(_03578_),
    .X(_03588_));
 sg13g2_and2_1 _09220_ (.A(net135),
    .B(_03588_),
    .X(_00531_));
 sg13g2_mux2_1 _09221_ (.A0(\shift_storage.storage [1387]),
    .A1(\shift_storage.storage [1386]),
    .S(_03578_),
    .X(_03589_));
 sg13g2_and2_1 _09222_ (.A(net135),
    .B(_03589_),
    .X(_00532_));
 sg13g2_buf_1 _09223_ (.A(_03540_),
    .X(_03590_));
 sg13g2_mux2_1 _09224_ (.A0(\shift_storage.storage [1388]),
    .A1(\shift_storage.storage [1387]),
    .S(net134),
    .X(_03591_));
 sg13g2_and2_1 _09225_ (.A(net135),
    .B(_03591_),
    .X(_00533_));
 sg13g2_mux2_1 _09226_ (.A0(\shift_storage.storage [1389]),
    .A1(\shift_storage.storage [1388]),
    .S(net134),
    .X(_03592_));
 sg13g2_and2_1 _09227_ (.A(net135),
    .B(_03592_),
    .X(_00534_));
 sg13g2_mux2_1 _09228_ (.A0(\shift_storage.storage [138]),
    .A1(\shift_storage.storage [137]),
    .S(net134),
    .X(_03593_));
 sg13g2_and2_1 _09229_ (.A(net135),
    .B(_03593_),
    .X(_00535_));
 sg13g2_mux2_1 _09230_ (.A0(\shift_storage.storage [1390]),
    .A1(\shift_storage.storage [1389]),
    .S(net134),
    .X(_03594_));
 sg13g2_and2_1 _09231_ (.A(net135),
    .B(_03594_),
    .X(_00536_));
 sg13g2_mux2_1 _09232_ (.A0(\shift_storage.storage [1391]),
    .A1(\shift_storage.storage [1390]),
    .S(net134),
    .X(_03595_));
 sg13g2_and2_1 _09233_ (.A(_03585_),
    .B(_03595_),
    .X(_00537_));
 sg13g2_mux2_1 _09234_ (.A0(\shift_storage.storage [1392]),
    .A1(\shift_storage.storage [1391]),
    .S(net134),
    .X(_03596_));
 sg13g2_and2_1 _09235_ (.A(_03585_),
    .B(_03596_),
    .X(_00538_));
 sg13g2_buf_1 _09236_ (.A(_03548_),
    .X(_03597_));
 sg13g2_mux2_1 _09237_ (.A0(\shift_storage.storage [1393]),
    .A1(\shift_storage.storage [1392]),
    .S(net134),
    .X(_03598_));
 sg13g2_and2_1 _09238_ (.A(net133),
    .B(_03598_),
    .X(_00539_));
 sg13g2_mux2_1 _09239_ (.A0(\shift_storage.storage [1394]),
    .A1(\shift_storage.storage [1393]),
    .S(net134),
    .X(_03599_));
 sg13g2_and2_1 _09240_ (.A(net133),
    .B(_03599_),
    .X(_00540_));
 sg13g2_mux2_1 _09241_ (.A0(\shift_storage.storage [1395]),
    .A1(\shift_storage.storage [1394]),
    .S(_03590_),
    .X(_03600_));
 sg13g2_and2_1 _09242_ (.A(net133),
    .B(_03600_),
    .X(_00541_));
 sg13g2_mux2_1 _09243_ (.A0(\shift_storage.storage [1396]),
    .A1(\shift_storage.storage [1395]),
    .S(_03590_),
    .X(_03601_));
 sg13g2_and2_1 _09244_ (.A(net133),
    .B(_03601_),
    .X(_00542_));
 sg13g2_buf_1 _09245_ (.A(_03540_),
    .X(_03602_));
 sg13g2_mux2_1 _09246_ (.A0(\shift_storage.storage [1397]),
    .A1(\shift_storage.storage [1396]),
    .S(net132),
    .X(_03603_));
 sg13g2_and2_1 _09247_ (.A(net133),
    .B(_03603_),
    .X(_00543_));
 sg13g2_mux2_1 _09248_ (.A0(\shift_storage.storage [1398]),
    .A1(\shift_storage.storage [1397]),
    .S(net132),
    .X(_03604_));
 sg13g2_and2_1 _09249_ (.A(_03597_),
    .B(_03604_),
    .X(_00544_));
 sg13g2_mux2_1 _09250_ (.A0(\shift_storage.storage [1399]),
    .A1(\shift_storage.storage [1398]),
    .S(net132),
    .X(_03605_));
 sg13g2_and2_1 _09251_ (.A(net133),
    .B(_03605_),
    .X(_00545_));
 sg13g2_mux2_1 _09252_ (.A0(\shift_storage.storage [139]),
    .A1(\shift_storage.storage [138]),
    .S(net132),
    .X(_03606_));
 sg13g2_and2_1 _09253_ (.A(net133),
    .B(_03606_),
    .X(_00546_));
 sg13g2_mux2_1 _09254_ (.A0(\shift_storage.storage [13]),
    .A1(\shift_storage.storage [12]),
    .S(net132),
    .X(_03607_));
 sg13g2_and2_1 _09255_ (.A(_03597_),
    .B(_03607_),
    .X(_00547_));
 sg13g2_mux2_1 _09256_ (.A0(\shift_storage.storage [1400]),
    .A1(\shift_storage.storage [1399]),
    .S(net132),
    .X(_03608_));
 sg13g2_and2_1 _09257_ (.A(net133),
    .B(_03608_),
    .X(_00548_));
 sg13g2_buf_1 _09258_ (.A(net363),
    .X(_03609_));
 sg13g2_mux2_1 _09259_ (.A0(\shift_storage.storage [1401]),
    .A1(\shift_storage.storage [1400]),
    .S(net132),
    .X(_03610_));
 sg13g2_and2_1 _09260_ (.A(net131),
    .B(_03610_),
    .X(_00549_));
 sg13g2_mux2_1 _09261_ (.A0(\shift_storage.storage [1402]),
    .A1(\shift_storage.storage [1401]),
    .S(net132),
    .X(_03611_));
 sg13g2_and2_1 _09262_ (.A(net131),
    .B(_03611_),
    .X(_00550_));
 sg13g2_mux2_1 _09263_ (.A0(\shift_storage.storage [1403]),
    .A1(\shift_storage.storage [1402]),
    .S(_03602_),
    .X(_03612_));
 sg13g2_and2_1 _09264_ (.A(net131),
    .B(_03612_),
    .X(_00551_));
 sg13g2_mux2_1 _09265_ (.A0(\shift_storage.storage [1404]),
    .A1(\shift_storage.storage [1403]),
    .S(_03602_),
    .X(_03613_));
 sg13g2_and2_1 _09266_ (.A(net131),
    .B(_03613_),
    .X(_00552_));
 sg13g2_buf_1 _09267_ (.A(net364),
    .X(_03614_));
 sg13g2_mux2_1 _09268_ (.A0(\shift_storage.storage [1405]),
    .A1(\shift_storage.storage [1404]),
    .S(net130),
    .X(_03615_));
 sg13g2_and2_1 _09269_ (.A(net131),
    .B(_03615_),
    .X(_00553_));
 sg13g2_mux2_1 _09270_ (.A0(\shift_storage.storage [1406]),
    .A1(\shift_storage.storage [1405]),
    .S(net130),
    .X(_03616_));
 sg13g2_and2_1 _09271_ (.A(_03609_),
    .B(_03616_),
    .X(_00554_));
 sg13g2_mux2_1 _09272_ (.A0(\shift_storage.storage [1407]),
    .A1(\shift_storage.storage [1406]),
    .S(_03614_),
    .X(_03617_));
 sg13g2_and2_1 _09273_ (.A(_03609_),
    .B(_03617_),
    .X(_00555_));
 sg13g2_mux2_1 _09274_ (.A0(\shift_storage.storage [1408]),
    .A1(\shift_storage.storage [1407]),
    .S(_03614_),
    .X(_03618_));
 sg13g2_and2_1 _09275_ (.A(net131),
    .B(_03618_),
    .X(_00556_));
 sg13g2_mux2_1 _09276_ (.A0(\shift_storage.storage [1409]),
    .A1(\shift_storage.storage [1408]),
    .S(net130),
    .X(_03619_));
 sg13g2_and2_1 _09277_ (.A(net131),
    .B(_03619_),
    .X(_00557_));
 sg13g2_mux2_1 _09278_ (.A0(\shift_storage.storage [140]),
    .A1(\shift_storage.storage [139]),
    .S(net130),
    .X(_03620_));
 sg13g2_and2_1 _09279_ (.A(net131),
    .B(_03620_),
    .X(_00558_));
 sg13g2_buf_1 _09280_ (.A(net363),
    .X(_03621_));
 sg13g2_mux2_1 _09281_ (.A0(\shift_storage.storage [1410]),
    .A1(\shift_storage.storage [1409]),
    .S(net130),
    .X(_03622_));
 sg13g2_and2_1 _09282_ (.A(net129),
    .B(_03622_),
    .X(_00559_));
 sg13g2_mux2_1 _09283_ (.A0(\shift_storage.storage [1411]),
    .A1(\shift_storage.storage [1410]),
    .S(net130),
    .X(_03623_));
 sg13g2_and2_1 _09284_ (.A(net129),
    .B(_03623_),
    .X(_00560_));
 sg13g2_mux2_1 _09285_ (.A0(\shift_storage.storage [1412]),
    .A1(\shift_storage.storage [1411]),
    .S(net130),
    .X(_03624_));
 sg13g2_and2_1 _09286_ (.A(net129),
    .B(_03624_),
    .X(_00561_));
 sg13g2_mux2_1 _09287_ (.A0(\shift_storage.storage [1413]),
    .A1(\shift_storage.storage [1412]),
    .S(net130),
    .X(_03625_));
 sg13g2_and2_1 _09288_ (.A(_03621_),
    .B(_03625_),
    .X(_00562_));
 sg13g2_buf_1 _09289_ (.A(net364),
    .X(_03626_));
 sg13g2_mux2_1 _09290_ (.A0(\shift_storage.storage [1414]),
    .A1(\shift_storage.storage [1413]),
    .S(net128),
    .X(_03627_));
 sg13g2_and2_1 _09291_ (.A(_03621_),
    .B(_03627_),
    .X(_00563_));
 sg13g2_mux2_1 _09292_ (.A0(\shift_storage.storage [1415]),
    .A1(\shift_storage.storage [1414]),
    .S(net128),
    .X(_03628_));
 sg13g2_and2_1 _09293_ (.A(net129),
    .B(_03628_),
    .X(_00564_));
 sg13g2_mux2_1 _09294_ (.A0(\shift_storage.storage [1416]),
    .A1(\shift_storage.storage [1415]),
    .S(net128),
    .X(_03629_));
 sg13g2_and2_1 _09295_ (.A(net129),
    .B(_03629_),
    .X(_00565_));
 sg13g2_mux2_1 _09296_ (.A0(\shift_storage.storage [1417]),
    .A1(\shift_storage.storage [1416]),
    .S(net128),
    .X(_03630_));
 sg13g2_and2_1 _09297_ (.A(net129),
    .B(_03630_),
    .X(_00566_));
 sg13g2_mux2_1 _09298_ (.A0(\shift_storage.storage [1418]),
    .A1(\shift_storage.storage [1417]),
    .S(_03626_),
    .X(_03631_));
 sg13g2_and2_1 _09299_ (.A(net129),
    .B(_03631_),
    .X(_00567_));
 sg13g2_mux2_1 _09300_ (.A0(\shift_storage.storage [1419]),
    .A1(\shift_storage.storage [1418]),
    .S(_03626_),
    .X(_03632_));
 sg13g2_and2_1 _09301_ (.A(net129),
    .B(_03632_),
    .X(_00568_));
 sg13g2_buf_1 _09302_ (.A(net363),
    .X(_03633_));
 sg13g2_mux2_1 _09303_ (.A0(\shift_storage.storage [141]),
    .A1(\shift_storage.storage [140]),
    .S(net128),
    .X(_03634_));
 sg13g2_and2_1 _09304_ (.A(net127),
    .B(_03634_),
    .X(_00569_));
 sg13g2_mux2_1 _09305_ (.A0(\shift_storage.storage [1420]),
    .A1(\shift_storage.storage [1419]),
    .S(net128),
    .X(_03635_));
 sg13g2_and2_1 _09306_ (.A(net127),
    .B(_03635_),
    .X(_00570_));
 sg13g2_mux2_1 _09307_ (.A0(\shift_storage.storage [1421]),
    .A1(\shift_storage.storage [1420]),
    .S(net128),
    .X(_03636_));
 sg13g2_and2_1 _09308_ (.A(_03633_),
    .B(_03636_),
    .X(_00571_));
 sg13g2_mux2_1 _09309_ (.A0(\shift_storage.storage [1422]),
    .A1(\shift_storage.storage [1421]),
    .S(net128),
    .X(_03637_));
 sg13g2_and2_1 _09310_ (.A(_03633_),
    .B(_03637_),
    .X(_00572_));
 sg13g2_buf_1 _09311_ (.A(net364),
    .X(_03638_));
 sg13g2_mux2_1 _09312_ (.A0(\shift_storage.storage [1423]),
    .A1(\shift_storage.storage [1422]),
    .S(net126),
    .X(_03639_));
 sg13g2_and2_1 _09313_ (.A(net127),
    .B(_03639_),
    .X(_00573_));
 sg13g2_mux2_1 _09314_ (.A0(\shift_storage.storage [1424]),
    .A1(\shift_storage.storage [1423]),
    .S(net126),
    .X(_03640_));
 sg13g2_and2_1 _09315_ (.A(net127),
    .B(_03640_),
    .X(_00574_));
 sg13g2_mux2_1 _09316_ (.A0(\shift_storage.storage [1425]),
    .A1(\shift_storage.storage [1424]),
    .S(net126),
    .X(_03641_));
 sg13g2_and2_1 _09317_ (.A(net127),
    .B(_03641_),
    .X(_00575_));
 sg13g2_mux2_1 _09318_ (.A0(\shift_storage.storage [1426]),
    .A1(\shift_storage.storage [1425]),
    .S(net126),
    .X(_03642_));
 sg13g2_and2_1 _09319_ (.A(net127),
    .B(_03642_),
    .X(_00576_));
 sg13g2_mux2_1 _09320_ (.A0(\shift_storage.storage [1427]),
    .A1(\shift_storage.storage [1426]),
    .S(net126),
    .X(_03643_));
 sg13g2_and2_1 _09321_ (.A(net127),
    .B(_03643_),
    .X(_00577_));
 sg13g2_mux2_1 _09322_ (.A0(\shift_storage.storage [1428]),
    .A1(\shift_storage.storage [1427]),
    .S(net126),
    .X(_03644_));
 sg13g2_and2_1 _09323_ (.A(net127),
    .B(_03644_),
    .X(_00578_));
 sg13g2_buf_1 _09324_ (.A(net363),
    .X(_03645_));
 sg13g2_mux2_1 _09325_ (.A0(\shift_storage.storage [1429]),
    .A1(\shift_storage.storage [1428]),
    .S(net126),
    .X(_03646_));
 sg13g2_and2_1 _09326_ (.A(net125),
    .B(_03646_),
    .X(_00579_));
 sg13g2_mux2_1 _09327_ (.A0(\shift_storage.storage [142]),
    .A1(\shift_storage.storage [141]),
    .S(net126),
    .X(_03647_));
 sg13g2_and2_1 _09328_ (.A(net125),
    .B(_03647_),
    .X(_00580_));
 sg13g2_mux2_1 _09329_ (.A0(\shift_storage.storage [1430]),
    .A1(\shift_storage.storage [1429]),
    .S(_03638_),
    .X(_03648_));
 sg13g2_and2_1 _09330_ (.A(net125),
    .B(_03648_),
    .X(_00581_));
 sg13g2_mux2_1 _09331_ (.A0(\shift_storage.storage [1431]),
    .A1(\shift_storage.storage [1430]),
    .S(_03638_),
    .X(_03649_));
 sg13g2_and2_1 _09332_ (.A(net125),
    .B(_03649_),
    .X(_00582_));
 sg13g2_buf_1 _09333_ (.A(net364),
    .X(_03650_));
 sg13g2_mux2_1 _09334_ (.A0(\shift_storage.storage [1432]),
    .A1(\shift_storage.storage [1431]),
    .S(net124),
    .X(_03651_));
 sg13g2_and2_1 _09335_ (.A(net125),
    .B(_03651_),
    .X(_00583_));
 sg13g2_mux2_1 _09336_ (.A0(\shift_storage.storage [1433]),
    .A1(\shift_storage.storage [1432]),
    .S(net124),
    .X(_03652_));
 sg13g2_and2_1 _09337_ (.A(net125),
    .B(_03652_),
    .X(_00584_));
 sg13g2_mux2_1 _09338_ (.A0(\shift_storage.storage [1434]),
    .A1(\shift_storage.storage [1433]),
    .S(net124),
    .X(_03653_));
 sg13g2_and2_1 _09339_ (.A(net125),
    .B(_03653_),
    .X(_00585_));
 sg13g2_mux2_1 _09340_ (.A0(\shift_storage.storage [1435]),
    .A1(\shift_storage.storage [1434]),
    .S(net124),
    .X(_03654_));
 sg13g2_and2_1 _09341_ (.A(net125),
    .B(_03654_),
    .X(_00586_));
 sg13g2_mux2_1 _09342_ (.A0(\shift_storage.storage [1436]),
    .A1(\shift_storage.storage [1435]),
    .S(net124),
    .X(_03655_));
 sg13g2_and2_1 _09343_ (.A(_03645_),
    .B(_03655_),
    .X(_00587_));
 sg13g2_mux2_1 _09344_ (.A0(\shift_storage.storage [1437]),
    .A1(\shift_storage.storage [1436]),
    .S(net124),
    .X(_03656_));
 sg13g2_and2_1 _09345_ (.A(_03645_),
    .B(_03656_),
    .X(_00588_));
 sg13g2_buf_1 _09346_ (.A(net363),
    .X(_03657_));
 sg13g2_mux2_1 _09347_ (.A0(\shift_storage.storage [1438]),
    .A1(\shift_storage.storage [1437]),
    .S(net124),
    .X(_03658_));
 sg13g2_and2_1 _09348_ (.A(net123),
    .B(_03658_),
    .X(_00589_));
 sg13g2_mux2_1 _09349_ (.A0(\shift_storage.storage [1439]),
    .A1(\shift_storage.storage [1438]),
    .S(net124),
    .X(_03659_));
 sg13g2_and2_1 _09350_ (.A(net123),
    .B(_03659_),
    .X(_00590_));
 sg13g2_mux2_1 _09351_ (.A0(\shift_storage.storage [143]),
    .A1(\shift_storage.storage [142]),
    .S(_03650_),
    .X(_03660_));
 sg13g2_and2_1 _09352_ (.A(net123),
    .B(_03660_),
    .X(_00591_));
 sg13g2_mux2_1 _09353_ (.A0(\shift_storage.storage [1440]),
    .A1(\shift_storage.storage [1439]),
    .S(_03650_),
    .X(_03661_));
 sg13g2_and2_1 _09354_ (.A(net123),
    .B(_03661_),
    .X(_00592_));
 sg13g2_buf_1 _09355_ (.A(net410),
    .X(_03662_));
 sg13g2_buf_1 _09356_ (.A(net362),
    .X(_03663_));
 sg13g2_mux2_1 _09357_ (.A0(\shift_storage.storage [1441]),
    .A1(\shift_storage.storage [1440]),
    .S(net122),
    .X(_03664_));
 sg13g2_and2_1 _09358_ (.A(net123),
    .B(_03664_),
    .X(_00593_));
 sg13g2_mux2_1 _09359_ (.A0(\shift_storage.storage [1442]),
    .A1(\shift_storage.storage [1441]),
    .S(net122),
    .X(_03665_));
 sg13g2_and2_1 _09360_ (.A(net123),
    .B(_03665_),
    .X(_00594_));
 sg13g2_mux2_1 _09361_ (.A0(\shift_storage.storage [1443]),
    .A1(\shift_storage.storage [1442]),
    .S(net122),
    .X(_03666_));
 sg13g2_and2_1 _09362_ (.A(net123),
    .B(_03666_),
    .X(_00595_));
 sg13g2_mux2_1 _09363_ (.A0(\shift_storage.storage [1444]),
    .A1(\shift_storage.storage [1443]),
    .S(net122),
    .X(_03667_));
 sg13g2_and2_1 _09364_ (.A(net123),
    .B(_03667_),
    .X(_00596_));
 sg13g2_mux2_1 _09365_ (.A0(\shift_storage.storage [1445]),
    .A1(\shift_storage.storage [1444]),
    .S(net122),
    .X(_03668_));
 sg13g2_and2_1 _09366_ (.A(_03657_),
    .B(_03668_),
    .X(_00597_));
 sg13g2_mux2_1 _09367_ (.A0(\shift_storage.storage [1446]),
    .A1(\shift_storage.storage [1445]),
    .S(_03663_),
    .X(_03669_));
 sg13g2_and2_1 _09368_ (.A(_03657_),
    .B(_03669_),
    .X(_00598_));
 sg13g2_buf_1 _09369_ (.A(net411),
    .X(_03670_));
 sg13g2_buf_1 _09370_ (.A(net361),
    .X(_03671_));
 sg13g2_mux2_1 _09371_ (.A0(\shift_storage.storage [1447]),
    .A1(\shift_storage.storage [1446]),
    .S(net122),
    .X(_03672_));
 sg13g2_and2_1 _09372_ (.A(net121),
    .B(_03672_),
    .X(_00599_));
 sg13g2_mux2_1 _09373_ (.A0(\shift_storage.storage [1448]),
    .A1(\shift_storage.storage [1447]),
    .S(net122),
    .X(_03673_));
 sg13g2_and2_1 _09374_ (.A(net121),
    .B(_03673_),
    .X(_00600_));
 sg13g2_mux2_1 _09375_ (.A0(\shift_storage.storage [1449]),
    .A1(\shift_storage.storage [1448]),
    .S(net122),
    .X(_03674_));
 sg13g2_and2_1 _09376_ (.A(net121),
    .B(_03674_),
    .X(_00601_));
 sg13g2_mux2_1 _09377_ (.A0(\shift_storage.storage [144]),
    .A1(\shift_storage.storage [143]),
    .S(_03663_),
    .X(_03675_));
 sg13g2_and2_1 _09378_ (.A(_03671_),
    .B(_03675_),
    .X(_00602_));
 sg13g2_buf_1 _09379_ (.A(net362),
    .X(_03676_));
 sg13g2_mux2_1 _09380_ (.A0(\shift_storage.storage [1450]),
    .A1(\shift_storage.storage [1449]),
    .S(net120),
    .X(_03677_));
 sg13g2_and2_1 _09381_ (.A(_03671_),
    .B(_03677_),
    .X(_00603_));
 sg13g2_mux2_1 _09382_ (.A0(\shift_storage.storage [1451]),
    .A1(\shift_storage.storage [1450]),
    .S(net120),
    .X(_03678_));
 sg13g2_and2_1 _09383_ (.A(net121),
    .B(_03678_),
    .X(_00604_));
 sg13g2_mux2_1 _09384_ (.A0(\shift_storage.storage [1452]),
    .A1(\shift_storage.storage [1451]),
    .S(net120),
    .X(_03679_));
 sg13g2_and2_1 _09385_ (.A(net121),
    .B(_03679_),
    .X(_00605_));
 sg13g2_mux2_1 _09386_ (.A0(\shift_storage.storage [1453]),
    .A1(\shift_storage.storage [1452]),
    .S(net120),
    .X(_03680_));
 sg13g2_and2_1 _09387_ (.A(net121),
    .B(_03680_),
    .X(_00606_));
 sg13g2_mux2_1 _09388_ (.A0(\shift_storage.storage [1454]),
    .A1(\shift_storage.storage [1453]),
    .S(net120),
    .X(_03681_));
 sg13g2_and2_1 _09389_ (.A(net121),
    .B(_03681_),
    .X(_00607_));
 sg13g2_mux2_1 _09390_ (.A0(\shift_storage.storage [1455]),
    .A1(\shift_storage.storage [1454]),
    .S(net120),
    .X(_03682_));
 sg13g2_and2_1 _09391_ (.A(net121),
    .B(_03682_),
    .X(_00608_));
 sg13g2_buf_1 _09392_ (.A(net361),
    .X(_03683_));
 sg13g2_mux2_1 _09393_ (.A0(\shift_storage.storage [1456]),
    .A1(\shift_storage.storage [1455]),
    .S(net120),
    .X(_03684_));
 sg13g2_and2_1 _09394_ (.A(net119),
    .B(_03684_),
    .X(_00609_));
 sg13g2_mux2_1 _09395_ (.A0(\shift_storage.storage [1457]),
    .A1(\shift_storage.storage [1456]),
    .S(net120),
    .X(_03685_));
 sg13g2_and2_1 _09396_ (.A(net119),
    .B(_03685_),
    .X(_00610_));
 sg13g2_mux2_1 _09397_ (.A0(\shift_storage.storage [1458]),
    .A1(\shift_storage.storage [1457]),
    .S(_03676_),
    .X(_03686_));
 sg13g2_and2_1 _09398_ (.A(net119),
    .B(_03686_),
    .X(_00611_));
 sg13g2_mux2_1 _09399_ (.A0(\shift_storage.storage [1459]),
    .A1(\shift_storage.storage [1458]),
    .S(_03676_),
    .X(_03687_));
 sg13g2_and2_1 _09400_ (.A(_03683_),
    .B(_03687_),
    .X(_00612_));
 sg13g2_buf_1 _09401_ (.A(net362),
    .X(_03688_));
 sg13g2_mux2_1 _09402_ (.A0(\shift_storage.storage [145]),
    .A1(\shift_storage.storage [144]),
    .S(_03688_),
    .X(_03689_));
 sg13g2_and2_1 _09403_ (.A(_03683_),
    .B(_03689_),
    .X(_00613_));
 sg13g2_mux2_1 _09404_ (.A0(\shift_storage.storage [1460]),
    .A1(\shift_storage.storage [1459]),
    .S(net118),
    .X(_03690_));
 sg13g2_and2_1 _09405_ (.A(net119),
    .B(_03690_),
    .X(_00614_));
 sg13g2_mux2_1 _09406_ (.A0(\shift_storage.storage [1461]),
    .A1(\shift_storage.storage [1460]),
    .S(net118),
    .X(_03691_));
 sg13g2_and2_1 _09407_ (.A(net119),
    .B(_03691_),
    .X(_00615_));
 sg13g2_mux2_1 _09408_ (.A0(\shift_storage.storage [1462]),
    .A1(\shift_storage.storage [1461]),
    .S(net118),
    .X(_03692_));
 sg13g2_and2_1 _09409_ (.A(net119),
    .B(_03692_),
    .X(_00616_));
 sg13g2_mux2_1 _09410_ (.A0(\shift_storage.storage [1463]),
    .A1(\shift_storage.storage [1462]),
    .S(net118),
    .X(_03693_));
 sg13g2_and2_1 _09411_ (.A(net119),
    .B(_03693_),
    .X(_00617_));
 sg13g2_mux2_1 _09412_ (.A0(\shift_storage.storage [1464]),
    .A1(\shift_storage.storage [1463]),
    .S(net118),
    .X(_03694_));
 sg13g2_and2_1 _09413_ (.A(net119),
    .B(_03694_),
    .X(_00618_));
 sg13g2_buf_1 _09414_ (.A(net361),
    .X(_03695_));
 sg13g2_mux2_1 _09415_ (.A0(\shift_storage.storage [1465]),
    .A1(\shift_storage.storage [1464]),
    .S(net118),
    .X(_03696_));
 sg13g2_and2_1 _09416_ (.A(net117),
    .B(_03696_),
    .X(_00619_));
 sg13g2_mux2_1 _09417_ (.A0(\shift_storage.storage [1466]),
    .A1(\shift_storage.storage [1465]),
    .S(net118),
    .X(_03697_));
 sg13g2_and2_1 _09418_ (.A(net117),
    .B(_03697_),
    .X(_00620_));
 sg13g2_mux2_1 _09419_ (.A0(\shift_storage.storage [1467]),
    .A1(\shift_storage.storage [1466]),
    .S(net118),
    .X(_03698_));
 sg13g2_and2_1 _09420_ (.A(net117),
    .B(_03698_),
    .X(_00621_));
 sg13g2_mux2_1 _09421_ (.A0(\shift_storage.storage [1468]),
    .A1(\shift_storage.storage [1467]),
    .S(_03688_),
    .X(_03699_));
 sg13g2_and2_1 _09422_ (.A(net117),
    .B(_03699_),
    .X(_00622_));
 sg13g2_buf_1 _09423_ (.A(net362),
    .X(_03700_));
 sg13g2_mux2_1 _09424_ (.A0(\shift_storage.storage [1469]),
    .A1(\shift_storage.storage [1468]),
    .S(net116),
    .X(_03701_));
 sg13g2_and2_1 _09425_ (.A(net117),
    .B(_03701_),
    .X(_00623_));
 sg13g2_mux2_1 _09426_ (.A0(\shift_storage.storage [146]),
    .A1(\shift_storage.storage [145]),
    .S(net116),
    .X(_03702_));
 sg13g2_and2_1 _09427_ (.A(_03695_),
    .B(_03702_),
    .X(_00624_));
 sg13g2_mux2_1 _09428_ (.A0(\shift_storage.storage [1470]),
    .A1(\shift_storage.storage [1469]),
    .S(net116),
    .X(_03703_));
 sg13g2_and2_1 _09429_ (.A(_03695_),
    .B(_03703_),
    .X(_00625_));
 sg13g2_mux2_1 _09430_ (.A0(\shift_storage.storage [1471]),
    .A1(\shift_storage.storage [1470]),
    .S(net116),
    .X(_03704_));
 sg13g2_and2_1 _09431_ (.A(net117),
    .B(_03704_),
    .X(_00626_));
 sg13g2_mux2_1 _09432_ (.A0(\shift_storage.storage [1472]),
    .A1(\shift_storage.storage [1471]),
    .S(net116),
    .X(_03705_));
 sg13g2_and2_1 _09433_ (.A(net117),
    .B(_03705_),
    .X(_00627_));
 sg13g2_mux2_1 _09434_ (.A0(\shift_storage.storage [1473]),
    .A1(\shift_storage.storage [1472]),
    .S(net116),
    .X(_03706_));
 sg13g2_and2_1 _09435_ (.A(net117),
    .B(_03706_),
    .X(_00628_));
 sg13g2_buf_1 _09436_ (.A(net361),
    .X(_03707_));
 sg13g2_mux2_1 _09437_ (.A0(\shift_storage.storage [1474]),
    .A1(\shift_storage.storage [1473]),
    .S(net116),
    .X(_03708_));
 sg13g2_and2_1 _09438_ (.A(net115),
    .B(_03708_),
    .X(_00629_));
 sg13g2_mux2_1 _09439_ (.A0(\shift_storage.storage [1475]),
    .A1(\shift_storage.storage [1474]),
    .S(net116),
    .X(_03709_));
 sg13g2_and2_1 _09440_ (.A(net115),
    .B(_03709_),
    .X(_00630_));
 sg13g2_mux2_1 _09441_ (.A0(\shift_storage.storage [1476]),
    .A1(\shift_storage.storage [1475]),
    .S(_03700_),
    .X(_03710_));
 sg13g2_and2_1 _09442_ (.A(net115),
    .B(_03710_),
    .X(_00631_));
 sg13g2_mux2_1 _09443_ (.A0(\shift_storage.storage [1477]),
    .A1(\shift_storage.storage [1476]),
    .S(_03700_),
    .X(_03711_));
 sg13g2_and2_1 _09444_ (.A(net115),
    .B(_03711_),
    .X(_00632_));
 sg13g2_buf_1 _09445_ (.A(net362),
    .X(_03712_));
 sg13g2_mux2_1 _09446_ (.A0(\shift_storage.storage [1478]),
    .A1(\shift_storage.storage [1477]),
    .S(net114),
    .X(_03713_));
 sg13g2_and2_1 _09447_ (.A(net115),
    .B(_03713_),
    .X(_00633_));
 sg13g2_mux2_1 _09448_ (.A0(\shift_storage.storage [1479]),
    .A1(\shift_storage.storage [1478]),
    .S(net114),
    .X(_03714_));
 sg13g2_and2_1 _09449_ (.A(net115),
    .B(_03714_),
    .X(_00634_));
 sg13g2_mux2_1 _09450_ (.A0(\shift_storage.storage [147]),
    .A1(\shift_storage.storage [146]),
    .S(net114),
    .X(_03715_));
 sg13g2_and2_1 _09451_ (.A(net115),
    .B(_03715_),
    .X(_00635_));
 sg13g2_mux2_1 _09452_ (.A0(\shift_storage.storage [1480]),
    .A1(\shift_storage.storage [1479]),
    .S(net114),
    .X(_03716_));
 sg13g2_and2_1 _09453_ (.A(net115),
    .B(_03716_),
    .X(_00636_));
 sg13g2_mux2_1 _09454_ (.A0(\shift_storage.storage [1481]),
    .A1(\shift_storage.storage [1480]),
    .S(net114),
    .X(_03717_));
 sg13g2_and2_1 _09455_ (.A(_03707_),
    .B(_03717_),
    .X(_00637_));
 sg13g2_mux2_1 _09456_ (.A0(\shift_storage.storage [1482]),
    .A1(\shift_storage.storage [1481]),
    .S(net114),
    .X(_03718_));
 sg13g2_and2_1 _09457_ (.A(_03707_),
    .B(_03718_),
    .X(_00638_));
 sg13g2_buf_1 _09458_ (.A(net361),
    .X(_03719_));
 sg13g2_mux2_1 _09459_ (.A0(\shift_storage.storage [1483]),
    .A1(\shift_storage.storage [1482]),
    .S(net114),
    .X(_03720_));
 sg13g2_and2_1 _09460_ (.A(net113),
    .B(_03720_),
    .X(_00639_));
 sg13g2_mux2_1 _09461_ (.A0(\shift_storage.storage [1484]),
    .A1(\shift_storage.storage [1483]),
    .S(net114),
    .X(_03721_));
 sg13g2_and2_1 _09462_ (.A(net113),
    .B(_03721_),
    .X(_00640_));
 sg13g2_mux2_1 _09463_ (.A0(\shift_storage.storage [1485]),
    .A1(\shift_storage.storage [1484]),
    .S(_03712_),
    .X(_03722_));
 sg13g2_and2_1 _09464_ (.A(_03719_),
    .B(_03722_),
    .X(_00641_));
 sg13g2_mux2_1 _09465_ (.A0(\shift_storage.storage [1486]),
    .A1(\shift_storage.storage [1485]),
    .S(_03712_),
    .X(_03723_));
 sg13g2_and2_1 _09466_ (.A(_03719_),
    .B(_03723_),
    .X(_00642_));
 sg13g2_buf_1 _09467_ (.A(net362),
    .X(_03724_));
 sg13g2_mux2_1 _09468_ (.A0(\shift_storage.storage [1487]),
    .A1(\shift_storage.storage [1486]),
    .S(net112),
    .X(_03725_));
 sg13g2_and2_1 _09469_ (.A(net113),
    .B(_03725_),
    .X(_00643_));
 sg13g2_mux2_1 _09470_ (.A0(\shift_storage.storage [1488]),
    .A1(\shift_storage.storage [1487]),
    .S(net112),
    .X(_03726_));
 sg13g2_and2_1 _09471_ (.A(net113),
    .B(_03726_),
    .X(_00644_));
 sg13g2_mux2_1 _09472_ (.A0(\shift_storage.storage [1489]),
    .A1(\shift_storage.storage [1488]),
    .S(net112),
    .X(_03727_));
 sg13g2_and2_1 _09473_ (.A(net113),
    .B(_03727_),
    .X(_00645_));
 sg13g2_mux2_1 _09474_ (.A0(\shift_storage.storage [148]),
    .A1(\shift_storage.storage [147]),
    .S(net112),
    .X(_03728_));
 sg13g2_and2_1 _09475_ (.A(net113),
    .B(_03728_),
    .X(_00646_));
 sg13g2_mux2_1 _09476_ (.A0(\shift_storage.storage [1490]),
    .A1(\shift_storage.storage [1489]),
    .S(_03724_),
    .X(_03729_));
 sg13g2_and2_1 _09477_ (.A(net113),
    .B(_03729_),
    .X(_00647_));
 sg13g2_mux2_1 _09478_ (.A0(\shift_storage.storage [1491]),
    .A1(\shift_storage.storage [1490]),
    .S(_03724_),
    .X(_03730_));
 sg13g2_and2_1 _09479_ (.A(net113),
    .B(_03730_),
    .X(_00648_));
 sg13g2_buf_1 _09480_ (.A(net361),
    .X(_03731_));
 sg13g2_mux2_1 _09481_ (.A0(\shift_storage.storage [1492]),
    .A1(\shift_storage.storage [1491]),
    .S(net112),
    .X(_03732_));
 sg13g2_and2_1 _09482_ (.A(net111),
    .B(_03732_),
    .X(_00649_));
 sg13g2_mux2_1 _09483_ (.A0(\shift_storage.storage [1493]),
    .A1(\shift_storage.storage [1492]),
    .S(net112),
    .X(_03733_));
 sg13g2_and2_1 _09484_ (.A(net111),
    .B(_03733_),
    .X(_00650_));
 sg13g2_mux2_1 _09485_ (.A0(\shift_storage.storage [1494]),
    .A1(\shift_storage.storage [1493]),
    .S(net112),
    .X(_03734_));
 sg13g2_and2_1 _09486_ (.A(net111),
    .B(_03734_),
    .X(_00651_));
 sg13g2_mux2_1 _09487_ (.A0(\shift_storage.storage [1495]),
    .A1(\shift_storage.storage [1494]),
    .S(net112),
    .X(_03735_));
 sg13g2_and2_1 _09488_ (.A(net111),
    .B(_03735_),
    .X(_00652_));
 sg13g2_buf_1 _09489_ (.A(net362),
    .X(_03736_));
 sg13g2_mux2_1 _09490_ (.A0(\shift_storage.storage [1496]),
    .A1(\shift_storage.storage [1495]),
    .S(net110),
    .X(_03737_));
 sg13g2_and2_1 _09491_ (.A(net111),
    .B(_03737_),
    .X(_00653_));
 sg13g2_mux2_1 _09492_ (.A0(\shift_storage.storage [1497]),
    .A1(\shift_storage.storage [1496]),
    .S(net110),
    .X(_03738_));
 sg13g2_and2_1 _09493_ (.A(net111),
    .B(_03738_),
    .X(_00654_));
 sg13g2_mux2_1 _09494_ (.A0(\shift_storage.storage [1498]),
    .A1(\shift_storage.storage [1497]),
    .S(net110),
    .X(_03739_));
 sg13g2_and2_1 _09495_ (.A(net111),
    .B(_03739_),
    .X(_00655_));
 sg13g2_mux2_1 _09496_ (.A0(\shift_storage.storage [1499]),
    .A1(\shift_storage.storage [1498]),
    .S(net110),
    .X(_03740_));
 sg13g2_and2_1 _09497_ (.A(net111),
    .B(_03740_),
    .X(_00656_));
 sg13g2_mux2_1 _09498_ (.A0(\shift_storage.storage [149]),
    .A1(\shift_storage.storage [148]),
    .S(_03736_),
    .X(_03741_));
 sg13g2_and2_1 _09499_ (.A(_03731_),
    .B(_03741_),
    .X(_00657_));
 sg13g2_mux2_1 _09500_ (.A0(\shift_storage.storage [14]),
    .A1(\shift_storage.storage [13]),
    .S(_03736_),
    .X(_03742_));
 sg13g2_and2_1 _09501_ (.A(_03731_),
    .B(_03742_),
    .X(_00658_));
 sg13g2_buf_1 _09502_ (.A(net361),
    .X(_03743_));
 sg13g2_mux2_1 _09503_ (.A0(\shift_storage.storage [1500]),
    .A1(\shift_storage.storage [1499]),
    .S(net110),
    .X(_03744_));
 sg13g2_and2_1 _09504_ (.A(net109),
    .B(_03744_),
    .X(_00659_));
 sg13g2_mux2_1 _09505_ (.A0(\shift_storage.storage [1501]),
    .A1(\shift_storage.storage [1500]),
    .S(net110),
    .X(_03745_));
 sg13g2_and2_1 _09506_ (.A(net109),
    .B(_03745_),
    .X(_00660_));
 sg13g2_mux2_1 _09507_ (.A0(\shift_storage.storage [1502]),
    .A1(\shift_storage.storage [1501]),
    .S(net110),
    .X(_03746_));
 sg13g2_and2_1 _09508_ (.A(net109),
    .B(_03746_),
    .X(_00661_));
 sg13g2_mux2_1 _09509_ (.A0(\shift_storage.storage [1503]),
    .A1(\shift_storage.storage [1502]),
    .S(net110),
    .X(_03747_));
 sg13g2_and2_1 _09510_ (.A(net109),
    .B(_03747_),
    .X(_00662_));
 sg13g2_buf_1 _09511_ (.A(net362),
    .X(_03748_));
 sg13g2_mux2_1 _09512_ (.A0(\shift_storage.storage [1504]),
    .A1(\shift_storage.storage [1503]),
    .S(net108),
    .X(_03749_));
 sg13g2_and2_1 _09513_ (.A(net109),
    .B(_03749_),
    .X(_00663_));
 sg13g2_mux2_1 _09514_ (.A0(\shift_storage.storage [1505]),
    .A1(\shift_storage.storage [1504]),
    .S(net108),
    .X(_03750_));
 sg13g2_and2_1 _09515_ (.A(net109),
    .B(_03750_),
    .X(_00664_));
 sg13g2_mux2_1 _09516_ (.A0(\shift_storage.storage [1506]),
    .A1(\shift_storage.storage [1505]),
    .S(net108),
    .X(_03751_));
 sg13g2_and2_1 _09517_ (.A(net109),
    .B(_03751_),
    .X(_00665_));
 sg13g2_mux2_1 _09518_ (.A0(\shift_storage.storage [1507]),
    .A1(\shift_storage.storage [1506]),
    .S(net108),
    .X(_03752_));
 sg13g2_and2_1 _09519_ (.A(net109),
    .B(_03752_),
    .X(_00666_));
 sg13g2_mux2_1 _09520_ (.A0(\shift_storage.storage [1508]),
    .A1(\shift_storage.storage [1507]),
    .S(net108),
    .X(_03753_));
 sg13g2_and2_1 _09521_ (.A(_03743_),
    .B(_03753_),
    .X(_00667_));
 sg13g2_mux2_1 _09522_ (.A0(\shift_storage.storage [1509]),
    .A1(\shift_storage.storage [1508]),
    .S(net108),
    .X(_03754_));
 sg13g2_and2_1 _09523_ (.A(_03743_),
    .B(_03754_),
    .X(_00668_));
 sg13g2_buf_1 _09524_ (.A(net361),
    .X(_03755_));
 sg13g2_mux2_1 _09525_ (.A0(\shift_storage.storage [150]),
    .A1(\shift_storage.storage [149]),
    .S(net108),
    .X(_03756_));
 sg13g2_and2_1 _09526_ (.A(net107),
    .B(_03756_),
    .X(_00669_));
 sg13g2_mux2_1 _09527_ (.A0(\shift_storage.storage [1510]),
    .A1(\shift_storage.storage [1509]),
    .S(_03748_),
    .X(_03757_));
 sg13g2_and2_1 _09528_ (.A(net107),
    .B(_03757_),
    .X(_00670_));
 sg13g2_mux2_1 _09529_ (.A0(\shift_storage.storage [1511]),
    .A1(\shift_storage.storage [1510]),
    .S(_03748_),
    .X(_03758_));
 sg13g2_and2_1 _09530_ (.A(net107),
    .B(_03758_),
    .X(_00671_));
 sg13g2_mux2_1 _09531_ (.A0(\shift_storage.storage [1512]),
    .A1(\shift_storage.storage [1511]),
    .S(net108),
    .X(_03759_));
 sg13g2_and2_1 _09532_ (.A(net107),
    .B(_03759_),
    .X(_00672_));
 sg13g2_buf_1 _09533_ (.A(_03662_),
    .X(_03760_));
 sg13g2_mux2_1 _09534_ (.A0(\shift_storage.storage [1513]),
    .A1(\shift_storage.storage [1512]),
    .S(net106),
    .X(_03761_));
 sg13g2_and2_1 _09535_ (.A(net107),
    .B(_03761_),
    .X(_00673_));
 sg13g2_mux2_1 _09536_ (.A0(\shift_storage.storage [1514]),
    .A1(\shift_storage.storage [1513]),
    .S(net106),
    .X(_03762_));
 sg13g2_and2_1 _09537_ (.A(net107),
    .B(_03762_),
    .X(_00674_));
 sg13g2_mux2_1 _09538_ (.A0(\shift_storage.storage [1515]),
    .A1(\shift_storage.storage [1514]),
    .S(net106),
    .X(_03763_));
 sg13g2_and2_1 _09539_ (.A(net107),
    .B(_03763_),
    .X(_00675_));
 sg13g2_mux2_1 _09540_ (.A0(\shift_storage.storage [1516]),
    .A1(\shift_storage.storage [1515]),
    .S(net106),
    .X(_03764_));
 sg13g2_and2_1 _09541_ (.A(net107),
    .B(_03764_),
    .X(_00676_));
 sg13g2_mux2_1 _09542_ (.A0(\shift_storage.storage [1517]),
    .A1(\shift_storage.storage [1516]),
    .S(net106),
    .X(_03765_));
 sg13g2_and2_1 _09543_ (.A(_03755_),
    .B(_03765_),
    .X(_00677_));
 sg13g2_mux2_1 _09544_ (.A0(\shift_storage.storage [1518]),
    .A1(\shift_storage.storage [1517]),
    .S(net106),
    .X(_03766_));
 sg13g2_and2_1 _09545_ (.A(_03755_),
    .B(_03766_),
    .X(_00678_));
 sg13g2_buf_1 _09546_ (.A(_03670_),
    .X(_03767_));
 sg13g2_mux2_1 _09547_ (.A0(\shift_storage.storage [1519]),
    .A1(\shift_storage.storage [1518]),
    .S(net106),
    .X(_03768_));
 sg13g2_and2_1 _09548_ (.A(net105),
    .B(_03768_),
    .X(_00679_));
 sg13g2_mux2_1 _09549_ (.A0(\shift_storage.storage [151]),
    .A1(\shift_storage.storage [150]),
    .S(net106),
    .X(_03769_));
 sg13g2_and2_1 _09550_ (.A(net105),
    .B(_03769_),
    .X(_00680_));
 sg13g2_mux2_1 _09551_ (.A0(\shift_storage.storage [1520]),
    .A1(\shift_storage.storage [1519]),
    .S(_03760_),
    .X(_03770_));
 sg13g2_and2_1 _09552_ (.A(net105),
    .B(_03770_),
    .X(_00681_));
 sg13g2_mux2_1 _09553_ (.A0(\shift_storage.storage [1521]),
    .A1(\shift_storage.storage [1520]),
    .S(_03760_),
    .X(_03771_));
 sg13g2_and2_1 _09554_ (.A(net105),
    .B(_03771_),
    .X(_00682_));
 sg13g2_buf_1 _09555_ (.A(_03662_),
    .X(_03772_));
 sg13g2_mux2_1 _09556_ (.A0(\shift_storage.storage [1522]),
    .A1(\shift_storage.storage [1521]),
    .S(net104),
    .X(_03773_));
 sg13g2_and2_1 _09557_ (.A(net105),
    .B(_03773_),
    .X(_00683_));
 sg13g2_mux2_1 _09558_ (.A0(\shift_storage.storage [1523]),
    .A1(\shift_storage.storage [1522]),
    .S(net104),
    .X(_03774_));
 sg13g2_and2_1 _09559_ (.A(_03767_),
    .B(_03774_),
    .X(_00684_));
 sg13g2_mux2_1 _09560_ (.A0(\shift_storage.storage [1524]),
    .A1(\shift_storage.storage [1523]),
    .S(net104),
    .X(_03775_));
 sg13g2_and2_1 _09561_ (.A(_03767_),
    .B(_03775_),
    .X(_00685_));
 sg13g2_mux2_1 _09562_ (.A0(\shift_storage.storage [1525]),
    .A1(\shift_storage.storage [1524]),
    .S(_03772_),
    .X(_03776_));
 sg13g2_and2_1 _09563_ (.A(net105),
    .B(_03776_),
    .X(_00686_));
 sg13g2_mux2_1 _09564_ (.A0(\shift_storage.storage [1526]),
    .A1(\shift_storage.storage [1525]),
    .S(_03772_),
    .X(_03777_));
 sg13g2_and2_1 _09565_ (.A(net105),
    .B(_03777_),
    .X(_00687_));
 sg13g2_mux2_1 _09566_ (.A0(\shift_storage.storage [1527]),
    .A1(\shift_storage.storage [1526]),
    .S(net104),
    .X(_03778_));
 sg13g2_and2_1 _09567_ (.A(net105),
    .B(_03778_),
    .X(_00688_));
 sg13g2_buf_1 _09568_ (.A(_03670_),
    .X(_03779_));
 sg13g2_mux2_1 _09569_ (.A0(\shift_storage.storage [1528]),
    .A1(\shift_storage.storage [1527]),
    .S(net104),
    .X(_03780_));
 sg13g2_and2_1 _09570_ (.A(net103),
    .B(_03780_),
    .X(_00689_));
 sg13g2_mux2_1 _09571_ (.A0(\shift_storage.storage [1529]),
    .A1(\shift_storage.storage [1528]),
    .S(net104),
    .X(_03781_));
 sg13g2_and2_1 _09572_ (.A(net103),
    .B(_03781_),
    .X(_00690_));
 sg13g2_mux2_1 _09573_ (.A0(\shift_storage.storage [152]),
    .A1(\shift_storage.storage [151]),
    .S(net104),
    .X(_03782_));
 sg13g2_and2_1 _09574_ (.A(net103),
    .B(_03782_),
    .X(_00691_));
 sg13g2_mux2_1 _09575_ (.A0(\shift_storage.storage [1530]),
    .A1(\shift_storage.storage [1529]),
    .S(net104),
    .X(_03783_));
 sg13g2_and2_1 _09576_ (.A(net103),
    .B(_03783_),
    .X(_00692_));
 sg13g2_buf_1 _09577_ (.A(net410),
    .X(_03784_));
 sg13g2_buf_1 _09578_ (.A(net360),
    .X(_03785_));
 sg13g2_mux2_1 _09579_ (.A0(\shift_storage.storage [1531]),
    .A1(\shift_storage.storage [1530]),
    .S(net102),
    .X(_03786_));
 sg13g2_and2_1 _09580_ (.A(net103),
    .B(_03786_),
    .X(_00693_));
 sg13g2_mux2_1 _09581_ (.A0(\shift_storage.storage [1532]),
    .A1(\shift_storage.storage [1531]),
    .S(net102),
    .X(_03787_));
 sg13g2_and2_1 _09582_ (.A(net103),
    .B(_03787_),
    .X(_00694_));
 sg13g2_mux2_1 _09583_ (.A0(\shift_storage.storage [1533]),
    .A1(\shift_storage.storage [1532]),
    .S(net102),
    .X(_03788_));
 sg13g2_and2_1 _09584_ (.A(net103),
    .B(_03788_),
    .X(_00695_));
 sg13g2_mux2_1 _09585_ (.A0(\shift_storage.storage [1534]),
    .A1(\shift_storage.storage [1533]),
    .S(net102),
    .X(_03789_));
 sg13g2_and2_1 _09586_ (.A(net103),
    .B(_03789_),
    .X(_00696_));
 sg13g2_mux2_1 _09587_ (.A0(\shift_storage.storage [1535]),
    .A1(\shift_storage.storage [1534]),
    .S(net102),
    .X(_03790_));
 sg13g2_and2_1 _09588_ (.A(_03779_),
    .B(_03790_),
    .X(_00697_));
 sg13g2_mux2_1 _09589_ (.A0(\shift_storage.storage [1536]),
    .A1(\shift_storage.storage [1535]),
    .S(net102),
    .X(_03791_));
 sg13g2_and2_1 _09590_ (.A(_03779_),
    .B(_03791_),
    .X(_00698_));
 sg13g2_buf_1 _09591_ (.A(net411),
    .X(_03792_));
 sg13g2_buf_1 _09592_ (.A(net359),
    .X(_03793_));
 sg13g2_mux2_1 _09593_ (.A0(\shift_storage.storage [1537]),
    .A1(\shift_storage.storage [1536]),
    .S(net102),
    .X(_03794_));
 sg13g2_and2_1 _09594_ (.A(net101),
    .B(_03794_),
    .X(_00699_));
 sg13g2_mux2_1 _09595_ (.A0(\shift_storage.storage [1538]),
    .A1(\shift_storage.storage [1537]),
    .S(_03785_),
    .X(_03795_));
 sg13g2_and2_1 _09596_ (.A(net101),
    .B(_03795_),
    .X(_00700_));
 sg13g2_mux2_1 _09597_ (.A0(\shift_storage.storage [1539]),
    .A1(\shift_storage.storage [1538]),
    .S(_03785_),
    .X(_03796_));
 sg13g2_and2_1 _09598_ (.A(net101),
    .B(_03796_),
    .X(_00701_));
 sg13g2_mux2_1 _09599_ (.A0(\shift_storage.storage [153]),
    .A1(\shift_storage.storage [152]),
    .S(net102),
    .X(_03797_));
 sg13g2_and2_1 _09600_ (.A(net101),
    .B(_03797_),
    .X(_00702_));
 sg13g2_buf_1 _09601_ (.A(net360),
    .X(_03798_));
 sg13g2_mux2_1 _09602_ (.A0(\shift_storage.storage [1540]),
    .A1(\shift_storage.storage [1539]),
    .S(net100),
    .X(_03799_));
 sg13g2_and2_1 _09603_ (.A(net101),
    .B(_03799_),
    .X(_00703_));
 sg13g2_mux2_1 _09604_ (.A0(\shift_storage.storage [1541]),
    .A1(\shift_storage.storage [1540]),
    .S(net100),
    .X(_03800_));
 sg13g2_and2_1 _09605_ (.A(net101),
    .B(_03800_),
    .X(_00704_));
 sg13g2_mux2_1 _09606_ (.A0(\shift_storage.storage [1542]),
    .A1(\shift_storage.storage [1541]),
    .S(net100),
    .X(_03801_));
 sg13g2_and2_1 _09607_ (.A(net101),
    .B(_03801_),
    .X(_00705_));
 sg13g2_mux2_1 _09608_ (.A0(\shift_storage.storage [1543]),
    .A1(\shift_storage.storage [1542]),
    .S(net100),
    .X(_03802_));
 sg13g2_and2_1 _09609_ (.A(net101),
    .B(_03802_),
    .X(_00706_));
 sg13g2_mux2_1 _09610_ (.A0(\shift_storage.storage [1544]),
    .A1(\shift_storage.storage [1543]),
    .S(net100),
    .X(_03803_));
 sg13g2_and2_1 _09611_ (.A(_03793_),
    .B(_03803_),
    .X(_00707_));
 sg13g2_mux2_1 _09612_ (.A0(\shift_storage.storage [1545]),
    .A1(\shift_storage.storage [1544]),
    .S(net100),
    .X(_03804_));
 sg13g2_and2_1 _09613_ (.A(_03793_),
    .B(_03804_),
    .X(_00708_));
 sg13g2_buf_1 _09614_ (.A(net359),
    .X(_03805_));
 sg13g2_mux2_1 _09615_ (.A0(\shift_storage.storage [1546]),
    .A1(\shift_storage.storage [1545]),
    .S(net100),
    .X(_03806_));
 sg13g2_and2_1 _09616_ (.A(net99),
    .B(_03806_),
    .X(_00709_));
 sg13g2_mux2_1 _09617_ (.A0(\shift_storage.storage [1547]),
    .A1(\shift_storage.storage [1546]),
    .S(net100),
    .X(_03807_));
 sg13g2_and2_1 _09618_ (.A(net99),
    .B(_03807_),
    .X(_00710_));
 sg13g2_mux2_1 _09619_ (.A0(\shift_storage.storage [1548]),
    .A1(\shift_storage.storage [1547]),
    .S(_03798_),
    .X(_03808_));
 sg13g2_and2_1 _09620_ (.A(_03805_),
    .B(_03808_),
    .X(_00711_));
 sg13g2_mux2_1 _09621_ (.A0(\shift_storage.storage [1549]),
    .A1(\shift_storage.storage [1548]),
    .S(_03798_),
    .X(_03809_));
 sg13g2_and2_1 _09622_ (.A(_03805_),
    .B(_03809_),
    .X(_00712_));
 sg13g2_buf_1 _09623_ (.A(net360),
    .X(_03810_));
 sg13g2_mux2_1 _09624_ (.A0(\shift_storage.storage [154]),
    .A1(\shift_storage.storage [153]),
    .S(net98),
    .X(_03811_));
 sg13g2_and2_1 _09625_ (.A(net99),
    .B(_03811_),
    .X(_00713_));
 sg13g2_mux2_1 _09626_ (.A0(\shift_storage.storage [1550]),
    .A1(\shift_storage.storage [1549]),
    .S(net98),
    .X(_03812_));
 sg13g2_and2_1 _09627_ (.A(net99),
    .B(_03812_),
    .X(_00714_));
 sg13g2_mux2_1 _09628_ (.A0(\shift_storage.storage [1551]),
    .A1(\shift_storage.storage [1550]),
    .S(net98),
    .X(_03813_));
 sg13g2_and2_1 _09629_ (.A(net99),
    .B(_03813_),
    .X(_00715_));
 sg13g2_mux2_1 _09630_ (.A0(\shift_storage.storage [1552]),
    .A1(\shift_storage.storage [1551]),
    .S(net98),
    .X(_03814_));
 sg13g2_and2_1 _09631_ (.A(net99),
    .B(_03814_),
    .X(_00716_));
 sg13g2_mux2_1 _09632_ (.A0(\shift_storage.storage [1553]),
    .A1(\shift_storage.storage [1552]),
    .S(net98),
    .X(_03815_));
 sg13g2_and2_1 _09633_ (.A(net99),
    .B(_03815_),
    .X(_00717_));
 sg13g2_mux2_1 _09634_ (.A0(\shift_storage.storage [1554]),
    .A1(\shift_storage.storage [1553]),
    .S(net98),
    .X(_03816_));
 sg13g2_and2_1 _09635_ (.A(net99),
    .B(_03816_),
    .X(_00718_));
 sg13g2_buf_1 _09636_ (.A(net359),
    .X(_03817_));
 sg13g2_mux2_1 _09637_ (.A0(\shift_storage.storage [1555]),
    .A1(\shift_storage.storage [1554]),
    .S(net98),
    .X(_03818_));
 sg13g2_and2_1 _09638_ (.A(net97),
    .B(_03818_),
    .X(_00719_));
 sg13g2_mux2_1 _09639_ (.A0(\shift_storage.storage [1556]),
    .A1(\shift_storage.storage [1555]),
    .S(net98),
    .X(_03819_));
 sg13g2_and2_1 _09640_ (.A(net97),
    .B(_03819_),
    .X(_00720_));
 sg13g2_mux2_1 _09641_ (.A0(\shift_storage.storage [1557]),
    .A1(\shift_storage.storage [1556]),
    .S(_03810_),
    .X(_03820_));
 sg13g2_and2_1 _09642_ (.A(net97),
    .B(_03820_),
    .X(_00721_));
 sg13g2_mux2_1 _09643_ (.A0(\shift_storage.storage [1558]),
    .A1(\shift_storage.storage [1557]),
    .S(_03810_),
    .X(_03821_));
 sg13g2_and2_1 _09644_ (.A(net97),
    .B(_03821_),
    .X(_00722_));
 sg13g2_buf_1 _09645_ (.A(net360),
    .X(_03822_));
 sg13g2_mux2_1 _09646_ (.A0(\shift_storage.storage [1559]),
    .A1(\shift_storage.storage [1558]),
    .S(net96),
    .X(_03823_));
 sg13g2_and2_1 _09647_ (.A(net97),
    .B(_03823_),
    .X(_00723_));
 sg13g2_mux2_1 _09648_ (.A0(\shift_storage.storage [155]),
    .A1(\shift_storage.storage [154]),
    .S(net96),
    .X(_03824_));
 sg13g2_and2_1 _09649_ (.A(net97),
    .B(_03824_),
    .X(_00724_));
 sg13g2_mux2_1 _09650_ (.A0(\shift_storage.storage [1560]),
    .A1(\shift_storage.storage [1559]),
    .S(net96),
    .X(_03825_));
 sg13g2_and2_1 _09651_ (.A(net97),
    .B(_03825_),
    .X(_00725_));
 sg13g2_mux2_1 _09652_ (.A0(\shift_storage.storage [1561]),
    .A1(\shift_storage.storage [1560]),
    .S(net96),
    .X(_03826_));
 sg13g2_and2_1 _09653_ (.A(net97),
    .B(_03826_),
    .X(_00726_));
 sg13g2_mux2_1 _09654_ (.A0(\shift_storage.storage [1562]),
    .A1(\shift_storage.storage [1561]),
    .S(net96),
    .X(_03827_));
 sg13g2_and2_1 _09655_ (.A(_03817_),
    .B(_03827_),
    .X(_00727_));
 sg13g2_mux2_1 _09656_ (.A0(\shift_storage.storage [1563]),
    .A1(\shift_storage.storage [1562]),
    .S(net96),
    .X(_03828_));
 sg13g2_and2_1 _09657_ (.A(_03817_),
    .B(_03828_),
    .X(_00728_));
 sg13g2_buf_1 _09658_ (.A(net359),
    .X(_03829_));
 sg13g2_mux2_1 _09659_ (.A0(\shift_storage.storage [1564]),
    .A1(\shift_storage.storage [1563]),
    .S(net96),
    .X(_03830_));
 sg13g2_and2_1 _09660_ (.A(net95),
    .B(_03830_),
    .X(_00729_));
 sg13g2_mux2_1 _09661_ (.A0(\shift_storage.storage [1565]),
    .A1(\shift_storage.storage [1564]),
    .S(net96),
    .X(_03831_));
 sg13g2_and2_1 _09662_ (.A(net95),
    .B(_03831_),
    .X(_00730_));
 sg13g2_mux2_1 _09663_ (.A0(\shift_storage.storage [1566]),
    .A1(\shift_storage.storage [1565]),
    .S(_03822_),
    .X(_03832_));
 sg13g2_and2_1 _09664_ (.A(net95),
    .B(_03832_),
    .X(_00731_));
 sg13g2_mux2_1 _09665_ (.A0(\shift_storage.storage [1567]),
    .A1(\shift_storage.storage [1566]),
    .S(_03822_),
    .X(_03833_));
 sg13g2_and2_1 _09666_ (.A(net95),
    .B(_03833_),
    .X(_00732_));
 sg13g2_buf_1 _09667_ (.A(net360),
    .X(_03834_));
 sg13g2_mux2_1 _09668_ (.A0(\shift_storage.storage [1568]),
    .A1(\shift_storage.storage [1567]),
    .S(net94),
    .X(_03835_));
 sg13g2_and2_1 _09669_ (.A(net95),
    .B(_03835_),
    .X(_00733_));
 sg13g2_mux2_1 _09670_ (.A0(\shift_storage.storage [1569]),
    .A1(\shift_storage.storage [1568]),
    .S(net94),
    .X(_03836_));
 sg13g2_and2_1 _09671_ (.A(_03829_),
    .B(_03836_),
    .X(_00734_));
 sg13g2_mux2_1 _09672_ (.A0(\shift_storage.storage [156]),
    .A1(\shift_storage.storage [155]),
    .S(net94),
    .X(_03837_));
 sg13g2_and2_1 _09673_ (.A(net95),
    .B(_03837_),
    .X(_00735_));
 sg13g2_mux2_1 _09674_ (.A0(\shift_storage.storage [1570]),
    .A1(\shift_storage.storage [1569]),
    .S(net94),
    .X(_03838_));
 sg13g2_and2_1 _09675_ (.A(_03829_),
    .B(_03838_),
    .X(_00736_));
 sg13g2_mux2_1 _09676_ (.A0(\shift_storage.storage [1571]),
    .A1(\shift_storage.storage [1570]),
    .S(net94),
    .X(_03839_));
 sg13g2_and2_1 _09677_ (.A(net95),
    .B(_03839_),
    .X(_00737_));
 sg13g2_mux2_1 _09678_ (.A0(\shift_storage.storage [1572]),
    .A1(\shift_storage.storage [1571]),
    .S(net94),
    .X(_03840_));
 sg13g2_and2_1 _09679_ (.A(net95),
    .B(_03840_),
    .X(_00738_));
 sg13g2_buf_1 _09680_ (.A(_03792_),
    .X(_03841_));
 sg13g2_mux2_1 _09681_ (.A0(\shift_storage.storage [1573]),
    .A1(\shift_storage.storage [1572]),
    .S(net94),
    .X(_03842_));
 sg13g2_and2_1 _09682_ (.A(net93),
    .B(_03842_),
    .X(_00739_));
 sg13g2_mux2_1 _09683_ (.A0(\shift_storage.storage [1574]),
    .A1(\shift_storage.storage [1573]),
    .S(net94),
    .X(_03843_));
 sg13g2_and2_1 _09684_ (.A(net93),
    .B(_03843_),
    .X(_00740_));
 sg13g2_mux2_1 _09685_ (.A0(\shift_storage.storage [1575]),
    .A1(\shift_storage.storage [1574]),
    .S(_03834_),
    .X(_03844_));
 sg13g2_and2_1 _09686_ (.A(net93),
    .B(_03844_),
    .X(_00741_));
 sg13g2_mux2_1 _09687_ (.A0(\shift_storage.storage [1576]),
    .A1(\shift_storage.storage [1575]),
    .S(_03834_),
    .X(_03845_));
 sg13g2_and2_1 _09688_ (.A(net93),
    .B(_03845_),
    .X(_00742_));
 sg13g2_buf_1 _09689_ (.A(_03784_),
    .X(_03846_));
 sg13g2_mux2_1 _09690_ (.A0(\shift_storage.storage [1577]),
    .A1(\shift_storage.storage [1576]),
    .S(net92),
    .X(_03847_));
 sg13g2_and2_1 _09691_ (.A(net93),
    .B(_03847_),
    .X(_00743_));
 sg13g2_mux2_1 _09692_ (.A0(\shift_storage.storage [1578]),
    .A1(\shift_storage.storage [1577]),
    .S(net92),
    .X(_03848_));
 sg13g2_and2_1 _09693_ (.A(net93),
    .B(_03848_),
    .X(_00744_));
 sg13g2_mux2_1 _09694_ (.A0(\shift_storage.storage [1579]),
    .A1(\shift_storage.storage [1578]),
    .S(net92),
    .X(_03849_));
 sg13g2_and2_1 _09695_ (.A(_03841_),
    .B(_03849_),
    .X(_00745_));
 sg13g2_mux2_1 _09696_ (.A0(\shift_storage.storage [157]),
    .A1(\shift_storage.storage [156]),
    .S(net92),
    .X(_03850_));
 sg13g2_and2_1 _09697_ (.A(net93),
    .B(_03850_),
    .X(_00746_));
 sg13g2_mux2_1 _09698_ (.A0(\shift_storage.storage [1580]),
    .A1(\shift_storage.storage [1579]),
    .S(_03846_),
    .X(_03851_));
 sg13g2_and2_1 _09699_ (.A(_03841_),
    .B(_03851_),
    .X(_00747_));
 sg13g2_mux2_1 _09700_ (.A0(\shift_storage.storage [1581]),
    .A1(\shift_storage.storage [1580]),
    .S(_03846_),
    .X(_03852_));
 sg13g2_and2_1 _09701_ (.A(net93),
    .B(_03852_),
    .X(_00748_));
 sg13g2_buf_1 _09702_ (.A(_03792_),
    .X(_03853_));
 sg13g2_mux2_1 _09703_ (.A0(\shift_storage.storage [1582]),
    .A1(\shift_storage.storage [1581]),
    .S(net92),
    .X(_03854_));
 sg13g2_and2_1 _09704_ (.A(net91),
    .B(_03854_),
    .X(_00749_));
 sg13g2_mux2_1 _09705_ (.A0(\shift_storage.storage [1583]),
    .A1(\shift_storage.storage [1582]),
    .S(net92),
    .X(_03855_));
 sg13g2_and2_1 _09706_ (.A(net91),
    .B(_03855_),
    .X(_00750_));
 sg13g2_mux2_1 _09707_ (.A0(\shift_storage.storage [1584]),
    .A1(\shift_storage.storage [1583]),
    .S(net92),
    .X(_03856_));
 sg13g2_and2_1 _09708_ (.A(net91),
    .B(_03856_),
    .X(_00751_));
 sg13g2_mux2_1 _09709_ (.A0(\shift_storage.storage [1585]),
    .A1(\shift_storage.storage [1584]),
    .S(net92),
    .X(_03857_));
 sg13g2_and2_1 _09710_ (.A(net91),
    .B(_03857_),
    .X(_00752_));
 sg13g2_buf_1 _09711_ (.A(_03784_),
    .X(_03858_));
 sg13g2_mux2_1 _09712_ (.A0(\shift_storage.storage [1586]),
    .A1(\shift_storage.storage [1585]),
    .S(net90),
    .X(_03859_));
 sg13g2_and2_1 _09713_ (.A(net91),
    .B(_03859_),
    .X(_00753_));
 sg13g2_mux2_1 _09714_ (.A0(\shift_storage.storage [1587]),
    .A1(\shift_storage.storage [1586]),
    .S(net90),
    .X(_03860_));
 sg13g2_and2_1 _09715_ (.A(_03853_),
    .B(_03860_),
    .X(_00754_));
 sg13g2_mux2_1 _09716_ (.A0(\shift_storage.storage [1588]),
    .A1(\shift_storage.storage [1587]),
    .S(_03858_),
    .X(_03861_));
 sg13g2_and2_1 _09717_ (.A(_03853_),
    .B(_03861_),
    .X(_00755_));
 sg13g2_mux2_1 _09718_ (.A0(\shift_storage.storage [1589]),
    .A1(\shift_storage.storage [1588]),
    .S(net90),
    .X(_03862_));
 sg13g2_and2_1 _09719_ (.A(net91),
    .B(_03862_),
    .X(_00756_));
 sg13g2_mux2_1 _09720_ (.A0(\shift_storage.storage [158]),
    .A1(\shift_storage.storage [157]),
    .S(net90),
    .X(_03863_));
 sg13g2_and2_1 _09721_ (.A(net91),
    .B(_03863_),
    .X(_00757_));
 sg13g2_mux2_1 _09722_ (.A0(\shift_storage.storage [1590]),
    .A1(\shift_storage.storage [1589]),
    .S(net90),
    .X(_03864_));
 sg13g2_and2_1 _09723_ (.A(net91),
    .B(_03864_),
    .X(_00758_));
 sg13g2_buf_1 _09724_ (.A(net359),
    .X(_03865_));
 sg13g2_mux2_1 _09725_ (.A0(\shift_storage.storage [1591]),
    .A1(\shift_storage.storage [1590]),
    .S(net90),
    .X(_03866_));
 sg13g2_and2_1 _09726_ (.A(net89),
    .B(_03866_),
    .X(_00759_));
 sg13g2_mux2_1 _09727_ (.A0(\shift_storage.storage [1592]),
    .A1(\shift_storage.storage [1591]),
    .S(net90),
    .X(_03867_));
 sg13g2_and2_1 _09728_ (.A(net89),
    .B(_03867_),
    .X(_00760_));
 sg13g2_mux2_1 _09729_ (.A0(\shift_storage.storage [1593]),
    .A1(\shift_storage.storage [1592]),
    .S(net90),
    .X(_03868_));
 sg13g2_and2_1 _09730_ (.A(net89),
    .B(_03868_),
    .X(_00761_));
 sg13g2_mux2_1 _09731_ (.A0(\shift_storage.storage [1594]),
    .A1(\shift_storage.storage [1593]),
    .S(_03858_),
    .X(_03869_));
 sg13g2_and2_1 _09732_ (.A(net89),
    .B(_03869_),
    .X(_00762_));
 sg13g2_buf_1 _09733_ (.A(net360),
    .X(_03870_));
 sg13g2_mux2_1 _09734_ (.A0(\shift_storage.storage [1595]),
    .A1(\shift_storage.storage [1594]),
    .S(net88),
    .X(_03871_));
 sg13g2_and2_1 _09735_ (.A(net89),
    .B(_03871_),
    .X(_00763_));
 sg13g2_mux2_1 _09736_ (.A0(\shift_storage.storage [1596]),
    .A1(\shift_storage.storage [1595]),
    .S(net88),
    .X(_03872_));
 sg13g2_and2_1 _09737_ (.A(net89),
    .B(_03872_),
    .X(_00764_));
 sg13g2_mux2_1 _09738_ (.A0(\shift_storage.storage [1597]),
    .A1(\shift_storage.storage [1596]),
    .S(net88),
    .X(_03873_));
 sg13g2_and2_1 _09739_ (.A(net89),
    .B(_03873_),
    .X(_00765_));
 sg13g2_mux2_1 _09740_ (.A0(\shift_storage.storage [1598]),
    .A1(\shift_storage.storage [1597]),
    .S(_03870_),
    .X(_03874_));
 sg13g2_and2_1 _09741_ (.A(_03865_),
    .B(_03874_),
    .X(_00766_));
 sg13g2_mux2_1 _09742_ (.A0(\shift_storage.shreg_out ),
    .A1(\shift_storage.storage [1598]),
    .S(_03870_),
    .X(_03875_));
 sg13g2_and2_1 _09743_ (.A(_03865_),
    .B(_03875_),
    .X(_00767_));
 sg13g2_mux2_1 _09744_ (.A0(\shift_storage.storage [159]),
    .A1(\shift_storage.storage [158]),
    .S(net88),
    .X(_03876_));
 sg13g2_and2_1 _09745_ (.A(net89),
    .B(_03876_),
    .X(_00768_));
 sg13g2_buf_1 _09746_ (.A(net359),
    .X(_03877_));
 sg13g2_mux2_1 _09747_ (.A0(\shift_storage.storage [15]),
    .A1(\shift_storage.storage [14]),
    .S(net88),
    .X(_03878_));
 sg13g2_and2_1 _09748_ (.A(net87),
    .B(_03878_),
    .X(_00769_));
 sg13g2_mux2_1 _09749_ (.A0(\shift_storage.storage [160]),
    .A1(\shift_storage.storage [159]),
    .S(net88),
    .X(_03879_));
 sg13g2_and2_1 _09750_ (.A(net87),
    .B(_03879_),
    .X(_00770_));
 sg13g2_mux2_1 _09751_ (.A0(\shift_storage.storage [161]),
    .A1(\shift_storage.storage [160]),
    .S(net88),
    .X(_03880_));
 sg13g2_and2_1 _09752_ (.A(net87),
    .B(_03880_),
    .X(_00771_));
 sg13g2_mux2_1 _09753_ (.A0(\shift_storage.storage [162]),
    .A1(\shift_storage.storage [161]),
    .S(net88),
    .X(_03881_));
 sg13g2_and2_1 _09754_ (.A(net87),
    .B(_03881_),
    .X(_00772_));
 sg13g2_buf_1 _09755_ (.A(net360),
    .X(_03882_));
 sg13g2_mux2_1 _09756_ (.A0(\shift_storage.storage [163]),
    .A1(\shift_storage.storage [162]),
    .S(net86),
    .X(_03883_));
 sg13g2_and2_1 _09757_ (.A(net87),
    .B(_03883_),
    .X(_00773_));
 sg13g2_mux2_1 _09758_ (.A0(\shift_storage.storage [164]),
    .A1(\shift_storage.storage [163]),
    .S(net86),
    .X(_03884_));
 sg13g2_and2_1 _09759_ (.A(net87),
    .B(_03884_),
    .X(_00774_));
 sg13g2_mux2_1 _09760_ (.A0(\shift_storage.storage [165]),
    .A1(\shift_storage.storage [164]),
    .S(net86),
    .X(_03885_));
 sg13g2_and2_1 _09761_ (.A(net87),
    .B(_03885_),
    .X(_00775_));
 sg13g2_mux2_1 _09762_ (.A0(\shift_storage.storage [166]),
    .A1(\shift_storage.storage [165]),
    .S(net86),
    .X(_03886_));
 sg13g2_and2_1 _09763_ (.A(_03877_),
    .B(_03886_),
    .X(_00776_));
 sg13g2_mux2_1 _09764_ (.A0(\shift_storage.storage [167]),
    .A1(\shift_storage.storage [166]),
    .S(_03882_),
    .X(_03887_));
 sg13g2_and2_1 _09765_ (.A(_03877_),
    .B(_03887_),
    .X(_00777_));
 sg13g2_mux2_1 _09766_ (.A0(\shift_storage.storage [168]),
    .A1(\shift_storage.storage [167]),
    .S(_03882_),
    .X(_03888_));
 sg13g2_and2_1 _09767_ (.A(net87),
    .B(_03888_),
    .X(_00778_));
 sg13g2_buf_1 _09768_ (.A(net359),
    .X(_03889_));
 sg13g2_mux2_1 _09769_ (.A0(\shift_storage.storage [169]),
    .A1(\shift_storage.storage [168]),
    .S(net86),
    .X(_03890_));
 sg13g2_and2_1 _09770_ (.A(net85),
    .B(_03890_),
    .X(_00779_));
 sg13g2_mux2_1 _09771_ (.A0(\shift_storage.storage [16]),
    .A1(\shift_storage.storage [15]),
    .S(net86),
    .X(_03891_));
 sg13g2_and2_1 _09772_ (.A(net85),
    .B(_03891_),
    .X(_00780_));
 sg13g2_mux2_1 _09773_ (.A0(\shift_storage.storage [170]),
    .A1(\shift_storage.storage [169]),
    .S(net86),
    .X(_03892_));
 sg13g2_and2_1 _09774_ (.A(_03889_),
    .B(_03892_),
    .X(_00781_));
 sg13g2_mux2_1 _09775_ (.A0(\shift_storage.storage [171]),
    .A1(\shift_storage.storage [170]),
    .S(net86),
    .X(_03893_));
 sg13g2_and2_1 _09776_ (.A(_03889_),
    .B(_03893_),
    .X(_00782_));
 sg13g2_buf_1 _09777_ (.A(net360),
    .X(_03894_));
 sg13g2_mux2_1 _09778_ (.A0(\shift_storage.storage [172]),
    .A1(\shift_storage.storage [171]),
    .S(net84),
    .X(_03895_));
 sg13g2_and2_1 _09779_ (.A(net85),
    .B(_03895_),
    .X(_00783_));
 sg13g2_mux2_1 _09780_ (.A0(\shift_storage.storage [173]),
    .A1(\shift_storage.storage [172]),
    .S(net84),
    .X(_03896_));
 sg13g2_and2_1 _09781_ (.A(net85),
    .B(_03896_),
    .X(_00784_));
 sg13g2_mux2_1 _09782_ (.A0(\shift_storage.storage [174]),
    .A1(\shift_storage.storage [173]),
    .S(net84),
    .X(_03897_));
 sg13g2_and2_1 _09783_ (.A(net85),
    .B(_03897_),
    .X(_00785_));
 sg13g2_mux2_1 _09784_ (.A0(\shift_storage.storage [175]),
    .A1(\shift_storage.storage [174]),
    .S(net84),
    .X(_03898_));
 sg13g2_and2_1 _09785_ (.A(net85),
    .B(_03898_),
    .X(_00786_));
 sg13g2_mux2_1 _09786_ (.A0(\shift_storage.storage [176]),
    .A1(\shift_storage.storage [175]),
    .S(_03894_),
    .X(_03899_));
 sg13g2_and2_1 _09787_ (.A(net85),
    .B(_03899_),
    .X(_00787_));
 sg13g2_mux2_1 _09788_ (.A0(\shift_storage.storage [177]),
    .A1(\shift_storage.storage [176]),
    .S(_03894_),
    .X(_03900_));
 sg13g2_and2_1 _09789_ (.A(net85),
    .B(_03900_),
    .X(_00788_));
 sg13g2_buf_1 _09790_ (.A(net359),
    .X(_03901_));
 sg13g2_mux2_1 _09791_ (.A0(\shift_storage.storage [178]),
    .A1(\shift_storage.storage [177]),
    .S(net84),
    .X(_03902_));
 sg13g2_and2_1 _09792_ (.A(net83),
    .B(_03902_),
    .X(_00789_));
 sg13g2_mux2_1 _09793_ (.A0(\shift_storage.storage [179]),
    .A1(\shift_storage.storage [178]),
    .S(net84),
    .X(_03903_));
 sg13g2_and2_1 _09794_ (.A(net83),
    .B(_03903_),
    .X(_00790_));
 sg13g2_mux2_1 _09795_ (.A0(\shift_storage.storage [17]),
    .A1(\shift_storage.storage [16]),
    .S(net84),
    .X(_03904_));
 sg13g2_and2_1 _09796_ (.A(net83),
    .B(_03904_),
    .X(_00791_));
 sg13g2_mux2_1 _09797_ (.A0(\shift_storage.storage [180]),
    .A1(\shift_storage.storage [179]),
    .S(net84),
    .X(_03905_));
 sg13g2_and2_1 _09798_ (.A(_03901_),
    .B(_03905_),
    .X(_00792_));
 sg13g2_buf_1 _09799_ (.A(_03059_),
    .X(_03906_));
 sg13g2_buf_1 _09800_ (.A(net358),
    .X(_03907_));
 sg13g2_mux2_1 _09801_ (.A0(\shift_storage.storage [181]),
    .A1(\shift_storage.storage [180]),
    .S(net82),
    .X(_03908_));
 sg13g2_and2_1 _09802_ (.A(_03901_),
    .B(_03908_),
    .X(_00793_));
 sg13g2_mux2_1 _09803_ (.A0(\shift_storage.storage [182]),
    .A1(\shift_storage.storage [181]),
    .S(net82),
    .X(_03909_));
 sg13g2_and2_1 _09804_ (.A(net83),
    .B(_03909_),
    .X(_00794_));
 sg13g2_mux2_1 _09805_ (.A0(\shift_storage.storage [183]),
    .A1(\shift_storage.storage [182]),
    .S(net82),
    .X(_03910_));
 sg13g2_and2_1 _09806_ (.A(net83),
    .B(_03910_),
    .X(_00795_));
 sg13g2_mux2_1 _09807_ (.A0(\shift_storage.storage [184]),
    .A1(\shift_storage.storage [183]),
    .S(net82),
    .X(_03911_));
 sg13g2_and2_1 _09808_ (.A(net83),
    .B(_03911_),
    .X(_00796_));
 sg13g2_mux2_1 _09809_ (.A0(\shift_storage.storage [185]),
    .A1(\shift_storage.storage [184]),
    .S(_03907_),
    .X(_03912_));
 sg13g2_and2_1 _09810_ (.A(net83),
    .B(_03912_),
    .X(_00797_));
 sg13g2_mux2_1 _09811_ (.A0(\shift_storage.storage [186]),
    .A1(\shift_storage.storage [185]),
    .S(_03907_),
    .X(_03913_));
 sg13g2_and2_1 _09812_ (.A(net83),
    .B(_03913_),
    .X(_00798_));
 sg13g2_buf_1 _09813_ (.A(net411),
    .X(_03914_));
 sg13g2_buf_1 _09814_ (.A(net357),
    .X(_03915_));
 sg13g2_mux2_1 _09815_ (.A0(\shift_storage.storage [187]),
    .A1(\shift_storage.storage [186]),
    .S(net82),
    .X(_03916_));
 sg13g2_and2_1 _09816_ (.A(net81),
    .B(_03916_),
    .X(_00799_));
 sg13g2_mux2_1 _09817_ (.A0(\shift_storage.storage [188]),
    .A1(\shift_storage.storage [187]),
    .S(net82),
    .X(_03917_));
 sg13g2_and2_1 _09818_ (.A(net81),
    .B(_03917_),
    .X(_00800_));
 sg13g2_mux2_1 _09819_ (.A0(\shift_storage.storage [189]),
    .A1(\shift_storage.storage [188]),
    .S(net82),
    .X(_03918_));
 sg13g2_and2_1 _09820_ (.A(_03915_),
    .B(_03918_),
    .X(_00801_));
 sg13g2_mux2_1 _09821_ (.A0(\shift_storage.storage [18]),
    .A1(\shift_storage.storage [17]),
    .S(net82),
    .X(_03919_));
 sg13g2_and2_1 _09822_ (.A(_03915_),
    .B(_03919_),
    .X(_00802_));
 sg13g2_buf_1 _09823_ (.A(net358),
    .X(_03920_));
 sg13g2_mux2_1 _09824_ (.A0(\shift_storage.storage [190]),
    .A1(\shift_storage.storage [189]),
    .S(net80),
    .X(_03921_));
 sg13g2_and2_1 _09825_ (.A(net81),
    .B(_03921_),
    .X(_00803_));
 sg13g2_mux2_1 _09826_ (.A0(\shift_storage.storage [191]),
    .A1(\shift_storage.storage [190]),
    .S(net80),
    .X(_03922_));
 sg13g2_and2_1 _09827_ (.A(net81),
    .B(_03922_),
    .X(_00804_));
 sg13g2_mux2_1 _09828_ (.A0(\shift_storage.storage [192]),
    .A1(\shift_storage.storage [191]),
    .S(net80),
    .X(_03923_));
 sg13g2_and2_1 _09829_ (.A(net81),
    .B(_03923_),
    .X(_00805_));
 sg13g2_mux2_1 _09830_ (.A0(\shift_storage.storage [193]),
    .A1(\shift_storage.storage [192]),
    .S(_03920_),
    .X(_03924_));
 sg13g2_and2_1 _09831_ (.A(net81),
    .B(_03924_),
    .X(_00806_));
 sg13g2_mux2_1 _09832_ (.A0(\shift_storage.storage [194]),
    .A1(\shift_storage.storage [193]),
    .S(_03920_),
    .X(_03925_));
 sg13g2_and2_1 _09833_ (.A(net81),
    .B(_03925_),
    .X(_00807_));
 sg13g2_mux2_1 _09834_ (.A0(\shift_storage.storage [195]),
    .A1(\shift_storage.storage [194]),
    .S(net80),
    .X(_03926_));
 sg13g2_and2_1 _09835_ (.A(net81),
    .B(_03926_),
    .X(_00808_));
 sg13g2_buf_1 _09836_ (.A(net357),
    .X(_03927_));
 sg13g2_mux2_1 _09837_ (.A0(\shift_storage.storage [196]),
    .A1(\shift_storage.storage [195]),
    .S(net80),
    .X(_03928_));
 sg13g2_and2_1 _09838_ (.A(net79),
    .B(_03928_),
    .X(_00809_));
 sg13g2_mux2_1 _09839_ (.A0(\shift_storage.storage [197]),
    .A1(\shift_storage.storage [196]),
    .S(net80),
    .X(_03929_));
 sg13g2_and2_1 _09840_ (.A(_03927_),
    .B(_03929_),
    .X(_00810_));
 sg13g2_mux2_1 _09841_ (.A0(\shift_storage.storage [198]),
    .A1(\shift_storage.storage [197]),
    .S(net80),
    .X(_03930_));
 sg13g2_and2_1 _09842_ (.A(net79),
    .B(_03930_),
    .X(_00811_));
 sg13g2_mux2_1 _09843_ (.A0(\shift_storage.storage [199]),
    .A1(\shift_storage.storage [198]),
    .S(net80),
    .X(_03931_));
 sg13g2_and2_1 _09844_ (.A(net79),
    .B(_03931_),
    .X(_00812_));
 sg13g2_buf_1 _09845_ (.A(net358),
    .X(_03932_));
 sg13g2_mux2_1 _09846_ (.A0(\shift_storage.storage [19]),
    .A1(\shift_storage.storage [18]),
    .S(net78),
    .X(_03933_));
 sg13g2_and2_1 _09847_ (.A(_03927_),
    .B(_03933_),
    .X(_00813_));
 sg13g2_mux2_1 _09848_ (.A0(\shift_storage.storage [1]),
    .A1(\shift_storage.storage [0]),
    .S(net78),
    .X(_03934_));
 sg13g2_and2_1 _09849_ (.A(net79),
    .B(_03934_),
    .X(_00814_));
 sg13g2_mux2_1 _09850_ (.A0(\shift_storage.storage [200]),
    .A1(\shift_storage.storage [199]),
    .S(net78),
    .X(_03935_));
 sg13g2_and2_1 _09851_ (.A(net79),
    .B(_03935_),
    .X(_00815_));
 sg13g2_mux2_1 _09852_ (.A0(\shift_storage.storage [201]),
    .A1(\shift_storage.storage [200]),
    .S(net78),
    .X(_03936_));
 sg13g2_and2_1 _09853_ (.A(net79),
    .B(_03936_),
    .X(_00816_));
 sg13g2_mux2_1 _09854_ (.A0(\shift_storage.storage [202]),
    .A1(\shift_storage.storage [201]),
    .S(net78),
    .X(_03937_));
 sg13g2_and2_1 _09855_ (.A(net79),
    .B(_03937_),
    .X(_00817_));
 sg13g2_mux2_1 _09856_ (.A0(\shift_storage.storage [203]),
    .A1(\shift_storage.storage [202]),
    .S(net78),
    .X(_03938_));
 sg13g2_and2_1 _09857_ (.A(net79),
    .B(_03938_),
    .X(_00818_));
 sg13g2_buf_1 _09858_ (.A(net357),
    .X(_03939_));
 sg13g2_mux2_1 _09859_ (.A0(\shift_storage.storage [204]),
    .A1(\shift_storage.storage [203]),
    .S(net78),
    .X(_03940_));
 sg13g2_and2_1 _09860_ (.A(net77),
    .B(_03940_),
    .X(_00819_));
 sg13g2_mux2_1 _09861_ (.A0(\shift_storage.storage [205]),
    .A1(\shift_storage.storage [204]),
    .S(net78),
    .X(_03941_));
 sg13g2_and2_1 _09862_ (.A(net77),
    .B(_03941_),
    .X(_00820_));
 sg13g2_mux2_1 _09863_ (.A0(\shift_storage.storage [206]),
    .A1(\shift_storage.storage [205]),
    .S(_03932_),
    .X(_03942_));
 sg13g2_and2_1 _09864_ (.A(net77),
    .B(_03942_),
    .X(_00821_));
 sg13g2_mux2_1 _09865_ (.A0(\shift_storage.storage [207]),
    .A1(\shift_storage.storage [206]),
    .S(_03932_),
    .X(_03943_));
 sg13g2_and2_1 _09866_ (.A(net77),
    .B(_03943_),
    .X(_00822_));
 sg13g2_buf_1 _09867_ (.A(net358),
    .X(_03944_));
 sg13g2_mux2_1 _09868_ (.A0(\shift_storage.storage [208]),
    .A1(\shift_storage.storage [207]),
    .S(net76),
    .X(_03945_));
 sg13g2_and2_1 _09869_ (.A(net77),
    .B(_03945_),
    .X(_00823_));
 sg13g2_mux2_1 _09870_ (.A0(\shift_storage.storage [209]),
    .A1(\shift_storage.storage [208]),
    .S(net76),
    .X(_03946_));
 sg13g2_and2_1 _09871_ (.A(net77),
    .B(_03946_),
    .X(_00824_));
 sg13g2_mux2_1 _09872_ (.A0(\shift_storage.storage [20]),
    .A1(\shift_storage.storage [19]),
    .S(net76),
    .X(_03947_));
 sg13g2_and2_1 _09873_ (.A(net77),
    .B(_03947_),
    .X(_00825_));
 sg13g2_mux2_1 _09874_ (.A0(\shift_storage.storage [210]),
    .A1(\shift_storage.storage [209]),
    .S(net76),
    .X(_03948_));
 sg13g2_and2_1 _09875_ (.A(net77),
    .B(_03948_),
    .X(_00826_));
 sg13g2_mux2_1 _09876_ (.A0(\shift_storage.storage [211]),
    .A1(\shift_storage.storage [210]),
    .S(net76),
    .X(_03949_));
 sg13g2_and2_1 _09877_ (.A(_03939_),
    .B(_03949_),
    .X(_00827_));
 sg13g2_mux2_1 _09878_ (.A0(\shift_storage.storage [212]),
    .A1(\shift_storage.storage [211]),
    .S(net76),
    .X(_03950_));
 sg13g2_and2_1 _09879_ (.A(_03939_),
    .B(_03950_),
    .X(_00828_));
 sg13g2_buf_1 _09880_ (.A(net357),
    .X(_03951_));
 sg13g2_mux2_1 _09881_ (.A0(\shift_storage.storage [213]),
    .A1(\shift_storage.storage [212]),
    .S(net76),
    .X(_03952_));
 sg13g2_and2_1 _09882_ (.A(net75),
    .B(_03952_),
    .X(_00829_));
 sg13g2_mux2_1 _09883_ (.A0(\shift_storage.storage [214]),
    .A1(\shift_storage.storage [213]),
    .S(net76),
    .X(_03953_));
 sg13g2_and2_1 _09884_ (.A(net75),
    .B(_03953_),
    .X(_00830_));
 sg13g2_mux2_1 _09885_ (.A0(\shift_storage.storage [215]),
    .A1(\shift_storage.storage [214]),
    .S(_03944_),
    .X(_03954_));
 sg13g2_and2_1 _09886_ (.A(net75),
    .B(_03954_),
    .X(_00831_));
 sg13g2_mux2_1 _09887_ (.A0(\shift_storage.storage [216]),
    .A1(\shift_storage.storage [215]),
    .S(_03944_),
    .X(_03955_));
 sg13g2_and2_1 _09888_ (.A(net75),
    .B(_03955_),
    .X(_00832_));
 sg13g2_buf_1 _09889_ (.A(net358),
    .X(_03956_));
 sg13g2_mux2_1 _09890_ (.A0(\shift_storage.storage [217]),
    .A1(\shift_storage.storage [216]),
    .S(net74),
    .X(_03957_));
 sg13g2_and2_1 _09891_ (.A(net75),
    .B(_03957_),
    .X(_00833_));
 sg13g2_mux2_1 _09892_ (.A0(\shift_storage.storage [218]),
    .A1(\shift_storage.storage [217]),
    .S(net74),
    .X(_03958_));
 sg13g2_and2_1 _09893_ (.A(net75),
    .B(_03958_),
    .X(_00834_));
 sg13g2_mux2_1 _09894_ (.A0(\shift_storage.storage [219]),
    .A1(\shift_storage.storage [218]),
    .S(net74),
    .X(_03959_));
 sg13g2_and2_1 _09895_ (.A(net75),
    .B(_03959_),
    .X(_00835_));
 sg13g2_mux2_1 _09896_ (.A0(\shift_storage.storage [21]),
    .A1(\shift_storage.storage [20]),
    .S(net74),
    .X(_03960_));
 sg13g2_and2_1 _09897_ (.A(net75),
    .B(_03960_),
    .X(_00836_));
 sg13g2_mux2_1 _09898_ (.A0(\shift_storage.storage [220]),
    .A1(\shift_storage.storage [219]),
    .S(net74),
    .X(_03961_));
 sg13g2_and2_1 _09899_ (.A(_03951_),
    .B(_03961_),
    .X(_00837_));
 sg13g2_mux2_1 _09900_ (.A0(\shift_storage.storage [221]),
    .A1(\shift_storage.storage [220]),
    .S(net74),
    .X(_03962_));
 sg13g2_and2_1 _09901_ (.A(_03951_),
    .B(_03962_),
    .X(_00838_));
 sg13g2_buf_1 _09902_ (.A(net357),
    .X(_03963_));
 sg13g2_mux2_1 _09903_ (.A0(\shift_storage.storage [222]),
    .A1(\shift_storage.storage [221]),
    .S(net74),
    .X(_03964_));
 sg13g2_and2_1 _09904_ (.A(net73),
    .B(_03964_),
    .X(_00839_));
 sg13g2_mux2_1 _09905_ (.A0(\shift_storage.storage [223]),
    .A1(\shift_storage.storage [222]),
    .S(net74),
    .X(_03965_));
 sg13g2_and2_1 _09906_ (.A(net73),
    .B(_03965_),
    .X(_00840_));
 sg13g2_mux2_1 _09907_ (.A0(\shift_storage.storage [224]),
    .A1(\shift_storage.storage [223]),
    .S(_03956_),
    .X(_03966_));
 sg13g2_and2_1 _09908_ (.A(net73),
    .B(_03966_),
    .X(_00841_));
 sg13g2_mux2_1 _09909_ (.A0(\shift_storage.storage [225]),
    .A1(\shift_storage.storage [224]),
    .S(_03956_),
    .X(_03967_));
 sg13g2_and2_1 _09910_ (.A(net73),
    .B(_03967_),
    .X(_00842_));
 sg13g2_buf_1 _09911_ (.A(net358),
    .X(_03968_));
 sg13g2_mux2_1 _09912_ (.A0(\shift_storage.storage [226]),
    .A1(\shift_storage.storage [225]),
    .S(net72),
    .X(_03969_));
 sg13g2_and2_1 _09913_ (.A(net73),
    .B(_03969_),
    .X(_00843_));
 sg13g2_mux2_1 _09914_ (.A0(\shift_storage.storage [227]),
    .A1(\shift_storage.storage [226]),
    .S(net72),
    .X(_03970_));
 sg13g2_and2_1 _09915_ (.A(net73),
    .B(_03970_),
    .X(_00844_));
 sg13g2_mux2_1 _09916_ (.A0(\shift_storage.storage [228]),
    .A1(\shift_storage.storage [227]),
    .S(net72),
    .X(_03971_));
 sg13g2_and2_1 _09917_ (.A(net73),
    .B(_03971_),
    .X(_00845_));
 sg13g2_mux2_1 _09918_ (.A0(\shift_storage.storage [229]),
    .A1(\shift_storage.storage [228]),
    .S(net72),
    .X(_03972_));
 sg13g2_and2_1 _09919_ (.A(_03963_),
    .B(_03972_),
    .X(_00846_));
 sg13g2_mux2_1 _09920_ (.A0(\shift_storage.storage [22]),
    .A1(\shift_storage.storage [21]),
    .S(net72),
    .X(_03973_));
 sg13g2_and2_1 _09921_ (.A(net73),
    .B(_03973_),
    .X(_00847_));
 sg13g2_mux2_1 _09922_ (.A0(\shift_storage.storage [230]),
    .A1(\shift_storage.storage [229]),
    .S(net72),
    .X(_03974_));
 sg13g2_and2_1 _09923_ (.A(_03963_),
    .B(_03974_),
    .X(_00848_));
 sg13g2_buf_1 _09924_ (.A(net357),
    .X(_03975_));
 sg13g2_mux2_1 _09925_ (.A0(\shift_storage.storage [231]),
    .A1(\shift_storage.storage [230]),
    .S(net72),
    .X(_03976_));
 sg13g2_and2_1 _09926_ (.A(net71),
    .B(_03976_),
    .X(_00849_));
 sg13g2_mux2_1 _09927_ (.A0(\shift_storage.storage [232]),
    .A1(\shift_storage.storage [231]),
    .S(net72),
    .X(_03977_));
 sg13g2_and2_1 _09928_ (.A(net71),
    .B(_03977_),
    .X(_00850_));
 sg13g2_mux2_1 _09929_ (.A0(\shift_storage.storage [233]),
    .A1(\shift_storage.storage [232]),
    .S(_03968_),
    .X(_03978_));
 sg13g2_and2_1 _09930_ (.A(net71),
    .B(_03978_),
    .X(_00851_));
 sg13g2_mux2_1 _09931_ (.A0(\shift_storage.storage [234]),
    .A1(\shift_storage.storage [233]),
    .S(_03968_),
    .X(_03979_));
 sg13g2_and2_1 _09932_ (.A(net71),
    .B(_03979_),
    .X(_00852_));
 sg13g2_buf_1 _09933_ (.A(_03906_),
    .X(_03980_));
 sg13g2_mux2_1 _09934_ (.A0(\shift_storage.storage [235]),
    .A1(\shift_storage.storage [234]),
    .S(net70),
    .X(_03981_));
 sg13g2_and2_1 _09935_ (.A(net71),
    .B(_03981_),
    .X(_00853_));
 sg13g2_mux2_1 _09936_ (.A0(\shift_storage.storage [236]),
    .A1(\shift_storage.storage [235]),
    .S(net70),
    .X(_03982_));
 sg13g2_and2_1 _09937_ (.A(net71),
    .B(_03982_),
    .X(_00854_));
 sg13g2_mux2_1 _09938_ (.A0(\shift_storage.storage [237]),
    .A1(\shift_storage.storage [236]),
    .S(net70),
    .X(_03983_));
 sg13g2_and2_1 _09939_ (.A(net71),
    .B(_03983_),
    .X(_00855_));
 sg13g2_mux2_1 _09940_ (.A0(\shift_storage.storage [238]),
    .A1(\shift_storage.storage [237]),
    .S(_03980_),
    .X(_03984_));
 sg13g2_and2_1 _09941_ (.A(_03975_),
    .B(_03984_),
    .X(_00856_));
 sg13g2_mux2_1 _09942_ (.A0(\shift_storage.storage [239]),
    .A1(\shift_storage.storage [238]),
    .S(_03980_),
    .X(_03985_));
 sg13g2_and2_1 _09943_ (.A(_03975_),
    .B(_03985_),
    .X(_00857_));
 sg13g2_mux2_1 _09944_ (.A0(\shift_storage.storage [23]),
    .A1(\shift_storage.storage [22]),
    .S(net70),
    .X(_03986_));
 sg13g2_and2_1 _09945_ (.A(net71),
    .B(_03986_),
    .X(_00858_));
 sg13g2_buf_1 _09946_ (.A(_03914_),
    .X(_03987_));
 sg13g2_mux2_1 _09947_ (.A0(\shift_storage.storage [240]),
    .A1(\shift_storage.storage [239]),
    .S(net70),
    .X(_03988_));
 sg13g2_and2_1 _09948_ (.A(net69),
    .B(_03988_),
    .X(_00859_));
 sg13g2_mux2_1 _09949_ (.A0(\shift_storage.storage [241]),
    .A1(\shift_storage.storage [240]),
    .S(net70),
    .X(_03989_));
 sg13g2_and2_1 _09950_ (.A(net69),
    .B(_03989_),
    .X(_00860_));
 sg13g2_mux2_1 _09951_ (.A0(\shift_storage.storage [242]),
    .A1(\shift_storage.storage [241]),
    .S(net70),
    .X(_03990_));
 sg13g2_and2_1 _09952_ (.A(net69),
    .B(_03990_),
    .X(_00861_));
 sg13g2_mux2_1 _09953_ (.A0(\shift_storage.storage [243]),
    .A1(\shift_storage.storage [242]),
    .S(net70),
    .X(_03991_));
 sg13g2_and2_1 _09954_ (.A(net69),
    .B(_03991_),
    .X(_00862_));
 sg13g2_buf_1 _09955_ (.A(_03906_),
    .X(_03992_));
 sg13g2_mux2_1 _09956_ (.A0(\shift_storage.storage [244]),
    .A1(\shift_storage.storage [243]),
    .S(net68),
    .X(_03993_));
 sg13g2_and2_1 _09957_ (.A(net69),
    .B(_03993_),
    .X(_00863_));
 sg13g2_mux2_1 _09958_ (.A0(\shift_storage.storage [245]),
    .A1(\shift_storage.storage [244]),
    .S(net68),
    .X(_03994_));
 sg13g2_and2_1 _09959_ (.A(net69),
    .B(_03994_),
    .X(_00864_));
 sg13g2_mux2_1 _09960_ (.A0(\shift_storage.storage [246]),
    .A1(\shift_storage.storage [245]),
    .S(net68),
    .X(_03995_));
 sg13g2_and2_1 _09961_ (.A(net69),
    .B(_03995_),
    .X(_00865_));
 sg13g2_mux2_1 _09962_ (.A0(\shift_storage.storage [247]),
    .A1(\shift_storage.storage [246]),
    .S(net68),
    .X(_03996_));
 sg13g2_and2_1 _09963_ (.A(net69),
    .B(_03996_),
    .X(_00866_));
 sg13g2_mux2_1 _09964_ (.A0(\shift_storage.storage [248]),
    .A1(\shift_storage.storage [247]),
    .S(net68),
    .X(_03997_));
 sg13g2_and2_1 _09965_ (.A(_03987_),
    .B(_03997_),
    .X(_00867_));
 sg13g2_mux2_1 _09966_ (.A0(\shift_storage.storage [249]),
    .A1(\shift_storage.storage [248]),
    .S(net68),
    .X(_03998_));
 sg13g2_and2_1 _09967_ (.A(_03987_),
    .B(_03998_),
    .X(_00868_));
 sg13g2_buf_1 _09968_ (.A(_03914_),
    .X(_03999_));
 sg13g2_mux2_1 _09969_ (.A0(\shift_storage.storage [24]),
    .A1(\shift_storage.storage [23]),
    .S(net68),
    .X(_04000_));
 sg13g2_and2_1 _09970_ (.A(net67),
    .B(_04000_),
    .X(_00869_));
 sg13g2_mux2_1 _09971_ (.A0(\shift_storage.storage [250]),
    .A1(\shift_storage.storage [249]),
    .S(net68),
    .X(_04001_));
 sg13g2_and2_1 _09972_ (.A(net67),
    .B(_04001_),
    .X(_00870_));
 sg13g2_mux2_1 _09973_ (.A0(\shift_storage.storage [251]),
    .A1(\shift_storage.storage [250]),
    .S(_03992_),
    .X(_04002_));
 sg13g2_and2_1 _09974_ (.A(net67),
    .B(_04002_),
    .X(_00871_));
 sg13g2_mux2_1 _09975_ (.A0(\shift_storage.storage [252]),
    .A1(\shift_storage.storage [251]),
    .S(_03992_),
    .X(_04003_));
 sg13g2_and2_1 _09976_ (.A(net67),
    .B(_04003_),
    .X(_00872_));
 sg13g2_buf_1 _09977_ (.A(net358),
    .X(_04004_));
 sg13g2_mux2_1 _09978_ (.A0(\shift_storage.storage [253]),
    .A1(\shift_storage.storage [252]),
    .S(net66),
    .X(_04005_));
 sg13g2_and2_1 _09979_ (.A(net67),
    .B(_04005_),
    .X(_00873_));
 sg13g2_mux2_1 _09980_ (.A0(\shift_storage.storage [254]),
    .A1(\shift_storage.storage [253]),
    .S(net66),
    .X(_04006_));
 sg13g2_and2_1 _09981_ (.A(_03999_),
    .B(_04006_),
    .X(_00874_));
 sg13g2_mux2_1 _09982_ (.A0(\shift_storage.storage [255]),
    .A1(\shift_storage.storage [254]),
    .S(net66),
    .X(_04007_));
 sg13g2_and2_1 _09983_ (.A(_03999_),
    .B(_04007_),
    .X(_00875_));
 sg13g2_mux2_1 _09984_ (.A0(\shift_storage.storage [256]),
    .A1(\shift_storage.storage [255]),
    .S(net66),
    .X(_04008_));
 sg13g2_and2_1 _09985_ (.A(net67),
    .B(_04008_),
    .X(_00876_));
 sg13g2_mux2_1 _09986_ (.A0(\shift_storage.storage [257]),
    .A1(\shift_storage.storage [256]),
    .S(net66),
    .X(_04009_));
 sg13g2_and2_1 _09987_ (.A(net67),
    .B(_04009_),
    .X(_00877_));
 sg13g2_mux2_1 _09988_ (.A0(\shift_storage.storage [258]),
    .A1(\shift_storage.storage [257]),
    .S(net66),
    .X(_04010_));
 sg13g2_and2_1 _09989_ (.A(net67),
    .B(_04010_),
    .X(_00878_));
 sg13g2_buf_1 _09990_ (.A(net357),
    .X(_04011_));
 sg13g2_mux2_1 _09991_ (.A0(\shift_storage.storage [259]),
    .A1(\shift_storage.storage [258]),
    .S(net66),
    .X(_04012_));
 sg13g2_and2_1 _09992_ (.A(net65),
    .B(_04012_),
    .X(_00879_));
 sg13g2_mux2_1 _09993_ (.A0(\shift_storage.storage [25]),
    .A1(\shift_storage.storage [24]),
    .S(net66),
    .X(_04013_));
 sg13g2_and2_1 _09994_ (.A(net65),
    .B(_04013_),
    .X(_00880_));
 sg13g2_mux2_1 _09995_ (.A0(\shift_storage.storage [260]),
    .A1(\shift_storage.storage [259]),
    .S(_04004_),
    .X(_04014_));
 sg13g2_and2_1 _09996_ (.A(net65),
    .B(_04014_),
    .X(_00881_));
 sg13g2_mux2_1 _09997_ (.A0(\shift_storage.storage [261]),
    .A1(\shift_storage.storage [260]),
    .S(_04004_),
    .X(_04015_));
 sg13g2_and2_1 _09998_ (.A(net65),
    .B(_04015_),
    .X(_00882_));
 sg13g2_buf_1 _09999_ (.A(net358),
    .X(_04016_));
 sg13g2_mux2_1 _10000_ (.A0(\shift_storage.storage [262]),
    .A1(\shift_storage.storage [261]),
    .S(net64),
    .X(_04017_));
 sg13g2_and2_1 _10001_ (.A(net65),
    .B(_04017_),
    .X(_00883_));
 sg13g2_mux2_1 _10002_ (.A0(\shift_storage.storage [263]),
    .A1(\shift_storage.storage [262]),
    .S(net64),
    .X(_04018_));
 sg13g2_and2_1 _10003_ (.A(_04011_),
    .B(_04018_),
    .X(_00884_));
 sg13g2_mux2_1 _10004_ (.A0(\shift_storage.storage [264]),
    .A1(\shift_storage.storage [263]),
    .S(_04016_),
    .X(_04019_));
 sg13g2_and2_1 _10005_ (.A(_04011_),
    .B(_04019_),
    .X(_00885_));
 sg13g2_mux2_1 _10006_ (.A0(\shift_storage.storage [265]),
    .A1(\shift_storage.storage [264]),
    .S(_04016_),
    .X(_04020_));
 sg13g2_and2_1 _10007_ (.A(net65),
    .B(_04020_),
    .X(_00886_));
 sg13g2_mux2_1 _10008_ (.A0(\shift_storage.storage [266]),
    .A1(\shift_storage.storage [265]),
    .S(net64),
    .X(_04021_));
 sg13g2_and2_1 _10009_ (.A(net65),
    .B(_04021_),
    .X(_00887_));
 sg13g2_mux2_1 _10010_ (.A0(\shift_storage.storage [267]),
    .A1(\shift_storage.storage [266]),
    .S(net64),
    .X(_04022_));
 sg13g2_and2_1 _10011_ (.A(net65),
    .B(_04022_),
    .X(_00888_));
 sg13g2_buf_1 _10012_ (.A(net357),
    .X(_04023_));
 sg13g2_mux2_1 _10013_ (.A0(\shift_storage.storage [268]),
    .A1(\shift_storage.storage [267]),
    .S(net64),
    .X(_04024_));
 sg13g2_and2_1 _10014_ (.A(net63),
    .B(_04024_),
    .X(_00889_));
 sg13g2_mux2_1 _10015_ (.A0(\shift_storage.storage [269]),
    .A1(\shift_storage.storage [268]),
    .S(net64),
    .X(_04025_));
 sg13g2_and2_1 _10016_ (.A(_04023_),
    .B(_04025_),
    .X(_00890_));
 sg13g2_mux2_1 _10017_ (.A0(\shift_storage.storage [26]),
    .A1(\shift_storage.storage [25]),
    .S(net64),
    .X(_04026_));
 sg13g2_and2_1 _10018_ (.A(_04023_),
    .B(_04026_),
    .X(_00891_));
 sg13g2_mux2_1 _10019_ (.A0(\shift_storage.storage [270]),
    .A1(\shift_storage.storage [269]),
    .S(net64),
    .X(_04027_));
 sg13g2_and2_1 _10020_ (.A(net63),
    .B(_04027_),
    .X(_00892_));
 sg13g2_buf_1 _10021_ (.A(_03059_),
    .X(_04028_));
 sg13g2_buf_1 _10022_ (.A(net356),
    .X(_04029_));
 sg13g2_mux2_1 _10023_ (.A0(\shift_storage.storage [271]),
    .A1(\shift_storage.storage [270]),
    .S(net62),
    .X(_04030_));
 sg13g2_and2_1 _10024_ (.A(net63),
    .B(_04030_),
    .X(_00893_));
 sg13g2_mux2_1 _10025_ (.A0(\shift_storage.storage [272]),
    .A1(\shift_storage.storage [271]),
    .S(net62),
    .X(_04031_));
 sg13g2_and2_1 _10026_ (.A(net63),
    .B(_04031_),
    .X(_00894_));
 sg13g2_mux2_1 _10027_ (.A0(\shift_storage.storage [273]),
    .A1(\shift_storage.storage [272]),
    .S(net62),
    .X(_04032_));
 sg13g2_and2_1 _10028_ (.A(net63),
    .B(_04032_),
    .X(_00895_));
 sg13g2_mux2_1 _10029_ (.A0(\shift_storage.storage [274]),
    .A1(\shift_storage.storage [273]),
    .S(net62),
    .X(_04033_));
 sg13g2_and2_1 _10030_ (.A(net63),
    .B(_04033_),
    .X(_00896_));
 sg13g2_mux2_1 _10031_ (.A0(\shift_storage.storage [275]),
    .A1(\shift_storage.storage [274]),
    .S(_04029_),
    .X(_04034_));
 sg13g2_and2_1 _10032_ (.A(net63),
    .B(_04034_),
    .X(_00897_));
 sg13g2_mux2_1 _10033_ (.A0(\shift_storage.storage [276]),
    .A1(\shift_storage.storage [275]),
    .S(_04029_),
    .X(_04035_));
 sg13g2_and2_1 _10034_ (.A(net63),
    .B(_04035_),
    .X(_00898_));
 sg13g2_buf_1 _10035_ (.A(_03050_),
    .X(_04036_));
 sg13g2_buf_1 _10036_ (.A(net355),
    .X(_04037_));
 sg13g2_mux2_1 _10037_ (.A0(\shift_storage.storage [277]),
    .A1(\shift_storage.storage [276]),
    .S(net62),
    .X(_04038_));
 sg13g2_and2_1 _10038_ (.A(net61),
    .B(_04038_),
    .X(_00899_));
 sg13g2_mux2_1 _10039_ (.A0(\shift_storage.storage [278]),
    .A1(\shift_storage.storage [277]),
    .S(net62),
    .X(_04039_));
 sg13g2_and2_1 _10040_ (.A(net61),
    .B(_04039_),
    .X(_00900_));
 sg13g2_mux2_1 _10041_ (.A0(\shift_storage.storage [279]),
    .A1(\shift_storage.storage [278]),
    .S(net62),
    .X(_04040_));
 sg13g2_and2_1 _10042_ (.A(net61),
    .B(_04040_),
    .X(_00901_));
 sg13g2_mux2_1 _10043_ (.A0(\shift_storage.storage [27]),
    .A1(\shift_storage.storage [26]),
    .S(net62),
    .X(_04041_));
 sg13g2_and2_1 _10044_ (.A(_04037_),
    .B(_04041_),
    .X(_00902_));
 sg13g2_buf_1 _10045_ (.A(net356),
    .X(_04042_));
 sg13g2_mux2_1 _10046_ (.A0(\shift_storage.storage [280]),
    .A1(\shift_storage.storage [279]),
    .S(net60),
    .X(_04043_));
 sg13g2_and2_1 _10047_ (.A(_04037_),
    .B(_04043_),
    .X(_00903_));
 sg13g2_mux2_1 _10048_ (.A0(\shift_storage.storage [281]),
    .A1(\shift_storage.storage [280]),
    .S(net60),
    .X(_04044_));
 sg13g2_and2_1 _10049_ (.A(net61),
    .B(_04044_),
    .X(_00904_));
 sg13g2_mux2_1 _10050_ (.A0(\shift_storage.storage [282]),
    .A1(\shift_storage.storage [281]),
    .S(net60),
    .X(_04045_));
 sg13g2_and2_1 _10051_ (.A(net61),
    .B(_04045_),
    .X(_00905_));
 sg13g2_mux2_1 _10052_ (.A0(\shift_storage.storage [283]),
    .A1(\shift_storage.storage [282]),
    .S(net60),
    .X(_04046_));
 sg13g2_and2_1 _10053_ (.A(net61),
    .B(_04046_),
    .X(_00906_));
 sg13g2_mux2_1 _10054_ (.A0(\shift_storage.storage [284]),
    .A1(\shift_storage.storage [283]),
    .S(net60),
    .X(_04047_));
 sg13g2_and2_1 _10055_ (.A(net61),
    .B(_04047_),
    .X(_00907_));
 sg13g2_mux2_1 _10056_ (.A0(\shift_storage.storage [285]),
    .A1(\shift_storage.storage [284]),
    .S(net60),
    .X(_04048_));
 sg13g2_and2_1 _10057_ (.A(net61),
    .B(_04048_),
    .X(_00908_));
 sg13g2_buf_1 _10058_ (.A(net355),
    .X(_04049_));
 sg13g2_mux2_1 _10059_ (.A0(\shift_storage.storage [286]),
    .A1(\shift_storage.storage [285]),
    .S(net60),
    .X(_04050_));
 sg13g2_and2_1 _10060_ (.A(net59),
    .B(_04050_),
    .X(_00909_));
 sg13g2_mux2_1 _10061_ (.A0(\shift_storage.storage [287]),
    .A1(\shift_storage.storage [286]),
    .S(net60),
    .X(_04051_));
 sg13g2_and2_1 _10062_ (.A(net59),
    .B(_04051_),
    .X(_00910_));
 sg13g2_mux2_1 _10063_ (.A0(\shift_storage.storage [288]),
    .A1(\shift_storage.storage [287]),
    .S(_04042_),
    .X(_04052_));
 sg13g2_and2_1 _10064_ (.A(net59),
    .B(_04052_),
    .X(_00911_));
 sg13g2_mux2_1 _10065_ (.A0(\shift_storage.storage [289]),
    .A1(\shift_storage.storage [288]),
    .S(_04042_),
    .X(_04053_));
 sg13g2_and2_1 _10066_ (.A(net59),
    .B(_04053_),
    .X(_00912_));
 sg13g2_buf_1 _10067_ (.A(net356),
    .X(_04054_));
 sg13g2_mux2_1 _10068_ (.A0(\shift_storage.storage [28]),
    .A1(\shift_storage.storage [27]),
    .S(net58),
    .X(_04055_));
 sg13g2_and2_1 _10069_ (.A(net59),
    .B(_04055_),
    .X(_00913_));
 sg13g2_mux2_1 _10070_ (.A0(\shift_storage.storage [290]),
    .A1(\shift_storage.storage [289]),
    .S(net58),
    .X(_04056_));
 sg13g2_and2_1 _10071_ (.A(_04049_),
    .B(_04056_),
    .X(_00914_));
 sg13g2_mux2_1 _10072_ (.A0(\shift_storage.storage [291]),
    .A1(\shift_storage.storage [290]),
    .S(_04054_),
    .X(_04057_));
 sg13g2_and2_1 _10073_ (.A(_04049_),
    .B(_04057_),
    .X(_00915_));
 sg13g2_mux2_1 _10074_ (.A0(\shift_storage.storage [292]),
    .A1(\shift_storage.storage [291]),
    .S(_04054_),
    .X(_04058_));
 sg13g2_and2_1 _10075_ (.A(net59),
    .B(_04058_),
    .X(_00916_));
 sg13g2_mux2_1 _10076_ (.A0(\shift_storage.storage [293]),
    .A1(\shift_storage.storage [292]),
    .S(net58),
    .X(_04059_));
 sg13g2_and2_1 _10077_ (.A(net59),
    .B(_04059_),
    .X(_00917_));
 sg13g2_mux2_1 _10078_ (.A0(\shift_storage.storage [294]),
    .A1(\shift_storage.storage [293]),
    .S(net58),
    .X(_04060_));
 sg13g2_and2_1 _10079_ (.A(net59),
    .B(_04060_),
    .X(_00918_));
 sg13g2_buf_1 _10080_ (.A(net355),
    .X(_04061_));
 sg13g2_mux2_1 _10081_ (.A0(\shift_storage.storage [295]),
    .A1(\shift_storage.storage [294]),
    .S(net58),
    .X(_04062_));
 sg13g2_and2_1 _10082_ (.A(net57),
    .B(_04062_),
    .X(_00919_));
 sg13g2_mux2_1 _10083_ (.A0(\shift_storage.storage [296]),
    .A1(\shift_storage.storage [295]),
    .S(net58),
    .X(_04063_));
 sg13g2_and2_1 _10084_ (.A(net57),
    .B(_04063_),
    .X(_00920_));
 sg13g2_mux2_1 _10085_ (.A0(\shift_storage.storage [297]),
    .A1(\shift_storage.storage [296]),
    .S(net58),
    .X(_04064_));
 sg13g2_and2_1 _10086_ (.A(net57),
    .B(_04064_),
    .X(_00921_));
 sg13g2_mux2_1 _10087_ (.A0(\shift_storage.storage [298]),
    .A1(\shift_storage.storage [297]),
    .S(net58),
    .X(_04065_));
 sg13g2_and2_1 _10088_ (.A(_04061_),
    .B(_04065_),
    .X(_00922_));
 sg13g2_buf_1 _10089_ (.A(net356),
    .X(_04066_));
 sg13g2_mux2_1 _10090_ (.A0(\shift_storage.storage [299]),
    .A1(\shift_storage.storage [298]),
    .S(net56),
    .X(_04067_));
 sg13g2_and2_1 _10091_ (.A(net57),
    .B(_04067_),
    .X(_00923_));
 sg13g2_mux2_1 _10092_ (.A0(\shift_storage.storage [29]),
    .A1(\shift_storage.storage [28]),
    .S(net56),
    .X(_04068_));
 sg13g2_and2_1 _10093_ (.A(_04061_),
    .B(_04068_),
    .X(_00924_));
 sg13g2_mux2_1 _10094_ (.A0(\shift_storage.storage [2]),
    .A1(\shift_storage.storage [1]),
    .S(net56),
    .X(_04069_));
 sg13g2_and2_1 _10095_ (.A(net57),
    .B(_04069_),
    .X(_00925_));
 sg13g2_mux2_1 _10096_ (.A0(\shift_storage.storage [300]),
    .A1(\shift_storage.storage [299]),
    .S(net56),
    .X(_04070_));
 sg13g2_and2_1 _10097_ (.A(net57),
    .B(_04070_),
    .X(_00926_));
 sg13g2_mux2_1 _10098_ (.A0(\shift_storage.storage [301]),
    .A1(\shift_storage.storage [300]),
    .S(net56),
    .X(_04071_));
 sg13g2_and2_1 _10099_ (.A(net57),
    .B(_04071_),
    .X(_00927_));
 sg13g2_mux2_1 _10100_ (.A0(\shift_storage.storage [302]),
    .A1(\shift_storage.storage [301]),
    .S(net56),
    .X(_04072_));
 sg13g2_and2_1 _10101_ (.A(net57),
    .B(_04072_),
    .X(_00928_));
 sg13g2_buf_1 _10102_ (.A(net355),
    .X(_04073_));
 sg13g2_mux2_1 _10103_ (.A0(\shift_storage.storage [303]),
    .A1(\shift_storage.storage [302]),
    .S(net56),
    .X(_04074_));
 sg13g2_and2_1 _10104_ (.A(net55),
    .B(_04074_),
    .X(_00929_));
 sg13g2_mux2_1 _10105_ (.A0(\shift_storage.storage [304]),
    .A1(\shift_storage.storage [303]),
    .S(net56),
    .X(_04075_));
 sg13g2_and2_1 _10106_ (.A(net55),
    .B(_04075_),
    .X(_00930_));
 sg13g2_mux2_1 _10107_ (.A0(\shift_storage.storage [305]),
    .A1(\shift_storage.storage [304]),
    .S(_04066_),
    .X(_04076_));
 sg13g2_and2_1 _10108_ (.A(net55),
    .B(_04076_),
    .X(_00931_));
 sg13g2_mux2_1 _10109_ (.A0(\shift_storage.storage [306]),
    .A1(\shift_storage.storage [305]),
    .S(_04066_),
    .X(_04077_));
 sg13g2_and2_1 _10110_ (.A(net55),
    .B(_04077_),
    .X(_00932_));
 sg13g2_buf_1 _10111_ (.A(net356),
    .X(_04078_));
 sg13g2_mux2_1 _10112_ (.A0(\shift_storage.storage [307]),
    .A1(\shift_storage.storage [306]),
    .S(net54),
    .X(_04079_));
 sg13g2_and2_1 _10113_ (.A(net55),
    .B(_04079_),
    .X(_00933_));
 sg13g2_mux2_1 _10114_ (.A0(\shift_storage.storage [308]),
    .A1(\shift_storage.storage [307]),
    .S(net54),
    .X(_04080_));
 sg13g2_and2_1 _10115_ (.A(net55),
    .B(_04080_),
    .X(_00934_));
 sg13g2_mux2_1 _10116_ (.A0(\shift_storage.storage [309]),
    .A1(\shift_storage.storage [308]),
    .S(net54),
    .X(_04081_));
 sg13g2_and2_1 _10117_ (.A(net55),
    .B(_04081_),
    .X(_00935_));
 sg13g2_mux2_1 _10118_ (.A0(\shift_storage.storage [30]),
    .A1(\shift_storage.storage [29]),
    .S(net54),
    .X(_04082_));
 sg13g2_and2_1 _10119_ (.A(net55),
    .B(_04082_),
    .X(_00936_));
 sg13g2_mux2_1 _10120_ (.A0(\shift_storage.storage [310]),
    .A1(\shift_storage.storage [309]),
    .S(net54),
    .X(_04083_));
 sg13g2_and2_1 _10121_ (.A(_04073_),
    .B(_04083_),
    .X(_00937_));
 sg13g2_mux2_1 _10122_ (.A0(\shift_storage.storage [311]),
    .A1(\shift_storage.storage [310]),
    .S(net54),
    .X(_04084_));
 sg13g2_and2_1 _10123_ (.A(_04073_),
    .B(_04084_),
    .X(_00938_));
 sg13g2_buf_1 _10124_ (.A(_04036_),
    .X(_04085_));
 sg13g2_mux2_1 _10125_ (.A0(\shift_storage.storage [312]),
    .A1(\shift_storage.storage [311]),
    .S(net54),
    .X(_04086_));
 sg13g2_and2_1 _10126_ (.A(net53),
    .B(_04086_),
    .X(_00939_));
 sg13g2_mux2_1 _10127_ (.A0(\shift_storage.storage [313]),
    .A1(\shift_storage.storage [312]),
    .S(net54),
    .X(_04087_));
 sg13g2_and2_1 _10128_ (.A(net53),
    .B(_04087_),
    .X(_00940_));
 sg13g2_mux2_1 _10129_ (.A0(\shift_storage.storage [314]),
    .A1(\shift_storage.storage [313]),
    .S(_04078_),
    .X(_04088_));
 sg13g2_and2_1 _10130_ (.A(net53),
    .B(_04088_),
    .X(_00941_));
 sg13g2_mux2_1 _10131_ (.A0(\shift_storage.storage [315]),
    .A1(\shift_storage.storage [314]),
    .S(_04078_),
    .X(_04089_));
 sg13g2_and2_1 _10132_ (.A(net53),
    .B(_04089_),
    .X(_00942_));
 sg13g2_buf_1 _10133_ (.A(_04028_),
    .X(_04090_));
 sg13g2_mux2_1 _10134_ (.A0(\shift_storage.storage [316]),
    .A1(\shift_storage.storage [315]),
    .S(net52),
    .X(_04091_));
 sg13g2_and2_1 _10135_ (.A(net53),
    .B(_04091_),
    .X(_00943_));
 sg13g2_mux2_1 _10136_ (.A0(\shift_storage.storage [317]),
    .A1(\shift_storage.storage [316]),
    .S(net52),
    .X(_04092_));
 sg13g2_and2_1 _10137_ (.A(net53),
    .B(_04092_),
    .X(_00944_));
 sg13g2_mux2_1 _10138_ (.A0(\shift_storage.storage [318]),
    .A1(\shift_storage.storage [317]),
    .S(net52),
    .X(_04093_));
 sg13g2_and2_1 _10139_ (.A(net53),
    .B(_04093_),
    .X(_00945_));
 sg13g2_mux2_1 _10140_ (.A0(\shift_storage.storage [319]),
    .A1(\shift_storage.storage [318]),
    .S(net52),
    .X(_04094_));
 sg13g2_and2_1 _10141_ (.A(net53),
    .B(_04094_),
    .X(_00946_));
 sg13g2_mux2_1 _10142_ (.A0(\shift_storage.storage [31]),
    .A1(\shift_storage.storage [30]),
    .S(net52),
    .X(_04095_));
 sg13g2_and2_1 _10143_ (.A(_04085_),
    .B(_04095_),
    .X(_00947_));
 sg13g2_mux2_1 _10144_ (.A0(\shift_storage.storage [320]),
    .A1(\shift_storage.storage [319]),
    .S(net52),
    .X(_04096_));
 sg13g2_and2_1 _10145_ (.A(_04085_),
    .B(_04096_),
    .X(_00948_));
 sg13g2_buf_1 _10146_ (.A(_04036_),
    .X(_04097_));
 sg13g2_mux2_1 _10147_ (.A0(\shift_storage.storage [321]),
    .A1(\shift_storage.storage [320]),
    .S(net52),
    .X(_04098_));
 sg13g2_and2_1 _10148_ (.A(net51),
    .B(_04098_),
    .X(_00949_));
 sg13g2_mux2_1 _10149_ (.A0(\shift_storage.storage [322]),
    .A1(\shift_storage.storage [321]),
    .S(net52),
    .X(_04099_));
 sg13g2_and2_1 _10150_ (.A(net51),
    .B(_04099_),
    .X(_00950_));
 sg13g2_mux2_1 _10151_ (.A0(\shift_storage.storage [323]),
    .A1(\shift_storage.storage [322]),
    .S(_04090_),
    .X(_04100_));
 sg13g2_and2_1 _10152_ (.A(net51),
    .B(_04100_),
    .X(_00951_));
 sg13g2_mux2_1 _10153_ (.A0(\shift_storage.storage [324]),
    .A1(\shift_storage.storage [323]),
    .S(_04090_),
    .X(_04101_));
 sg13g2_and2_1 _10154_ (.A(net51),
    .B(_04101_),
    .X(_00952_));
 sg13g2_buf_1 _10155_ (.A(_04028_),
    .X(_04102_));
 sg13g2_mux2_1 _10156_ (.A0(\shift_storage.storage [325]),
    .A1(\shift_storage.storage [324]),
    .S(net50),
    .X(_04103_));
 sg13g2_and2_1 _10157_ (.A(_04097_),
    .B(_04103_),
    .X(_00953_));
 sg13g2_mux2_1 _10158_ (.A0(\shift_storage.storage [326]),
    .A1(\shift_storage.storage [325]),
    .S(_04102_),
    .X(_04104_));
 sg13g2_and2_1 _10159_ (.A(_04097_),
    .B(_04104_),
    .X(_00954_));
 sg13g2_mux2_1 _10160_ (.A0(\shift_storage.storage [327]),
    .A1(\shift_storage.storage [326]),
    .S(_04102_),
    .X(_04105_));
 sg13g2_and2_1 _10161_ (.A(net51),
    .B(_04105_),
    .X(_00955_));
 sg13g2_mux2_1 _10162_ (.A0(\shift_storage.storage [328]),
    .A1(\shift_storage.storage [327]),
    .S(net50),
    .X(_04106_));
 sg13g2_and2_1 _10163_ (.A(net51),
    .B(_04106_),
    .X(_00956_));
 sg13g2_mux2_1 _10164_ (.A0(\shift_storage.storage [329]),
    .A1(\shift_storage.storage [328]),
    .S(net50),
    .X(_04107_));
 sg13g2_and2_1 _10165_ (.A(net51),
    .B(_04107_),
    .X(_00957_));
 sg13g2_mux2_1 _10166_ (.A0(\shift_storage.storage [32]),
    .A1(\shift_storage.storage [31]),
    .S(net50),
    .X(_04108_));
 sg13g2_and2_1 _10167_ (.A(net51),
    .B(_04108_),
    .X(_00958_));
 sg13g2_buf_1 _10168_ (.A(net355),
    .X(_04109_));
 sg13g2_mux2_1 _10169_ (.A0(\shift_storage.storage [330]),
    .A1(\shift_storage.storage [329]),
    .S(net50),
    .X(_04110_));
 sg13g2_and2_1 _10170_ (.A(net49),
    .B(_04110_),
    .X(_00959_));
 sg13g2_mux2_1 _10171_ (.A0(\shift_storage.storage [331]),
    .A1(\shift_storage.storage [330]),
    .S(net50),
    .X(_04111_));
 sg13g2_and2_1 _10172_ (.A(net49),
    .B(_04111_),
    .X(_00960_));
 sg13g2_mux2_1 _10173_ (.A0(\shift_storage.storage [332]),
    .A1(\shift_storage.storage [331]),
    .S(net50),
    .X(_04112_));
 sg13g2_and2_1 _10174_ (.A(net49),
    .B(_04112_),
    .X(_00961_));
 sg13g2_mux2_1 _10175_ (.A0(\shift_storage.storage [333]),
    .A1(\shift_storage.storage [332]),
    .S(net50),
    .X(_04113_));
 sg13g2_and2_1 _10176_ (.A(net49),
    .B(_04113_),
    .X(_00962_));
 sg13g2_buf_1 _10177_ (.A(net356),
    .X(_04114_));
 sg13g2_mux2_1 _10178_ (.A0(\shift_storage.storage [334]),
    .A1(\shift_storage.storage [333]),
    .S(net48),
    .X(_04115_));
 sg13g2_and2_1 _10179_ (.A(net49),
    .B(_04115_),
    .X(_00963_));
 sg13g2_mux2_1 _10180_ (.A0(\shift_storage.storage [335]),
    .A1(\shift_storage.storage [334]),
    .S(net48),
    .X(_04116_));
 sg13g2_and2_1 _10181_ (.A(net49),
    .B(_04116_),
    .X(_00964_));
 sg13g2_mux2_1 _10182_ (.A0(\shift_storage.storage [336]),
    .A1(\shift_storage.storage [335]),
    .S(net48),
    .X(_04117_));
 sg13g2_and2_1 _10183_ (.A(net49),
    .B(_04117_),
    .X(_00965_));
 sg13g2_mux2_1 _10184_ (.A0(\shift_storage.storage [337]),
    .A1(\shift_storage.storage [336]),
    .S(net48),
    .X(_04118_));
 sg13g2_and2_1 _10185_ (.A(net49),
    .B(_04118_),
    .X(_00966_));
 sg13g2_mux2_1 _10186_ (.A0(\shift_storage.storage [338]),
    .A1(\shift_storage.storage [337]),
    .S(net48),
    .X(_04119_));
 sg13g2_and2_1 _10187_ (.A(_04109_),
    .B(_04119_),
    .X(_00967_));
 sg13g2_mux2_1 _10188_ (.A0(\shift_storage.storage [339]),
    .A1(\shift_storage.storage [338]),
    .S(net48),
    .X(_04120_));
 sg13g2_and2_1 _10189_ (.A(_04109_),
    .B(_04120_),
    .X(_00968_));
 sg13g2_buf_1 _10190_ (.A(net355),
    .X(_04121_));
 sg13g2_mux2_1 _10191_ (.A0(\shift_storage.storage [33]),
    .A1(\shift_storage.storage [32]),
    .S(net48),
    .X(_04122_));
 sg13g2_and2_1 _10192_ (.A(net47),
    .B(_04122_),
    .X(_00969_));
 sg13g2_mux2_1 _10193_ (.A0(\shift_storage.storage [340]),
    .A1(\shift_storage.storage [339]),
    .S(net48),
    .X(_04123_));
 sg13g2_and2_1 _10194_ (.A(net47),
    .B(_04123_),
    .X(_00970_));
 sg13g2_mux2_1 _10195_ (.A0(\shift_storage.storage [341]),
    .A1(\shift_storage.storage [340]),
    .S(_04114_),
    .X(_04124_));
 sg13g2_and2_1 _10196_ (.A(net47),
    .B(_04124_),
    .X(_00971_));
 sg13g2_mux2_1 _10197_ (.A0(\shift_storage.storage [342]),
    .A1(\shift_storage.storage [341]),
    .S(_04114_),
    .X(_04125_));
 sg13g2_and2_1 _10198_ (.A(_04121_),
    .B(_04125_),
    .X(_00972_));
 sg13g2_buf_1 _10199_ (.A(net356),
    .X(_04126_));
 sg13g2_mux2_1 _10200_ (.A0(\shift_storage.storage [343]),
    .A1(\shift_storage.storage [342]),
    .S(net46),
    .X(_04127_));
 sg13g2_and2_1 _10201_ (.A(_04121_),
    .B(_04127_),
    .X(_00973_));
 sg13g2_mux2_1 _10202_ (.A0(\shift_storage.storage [344]),
    .A1(\shift_storage.storage [343]),
    .S(net46),
    .X(_04128_));
 sg13g2_and2_1 _10203_ (.A(net47),
    .B(_04128_),
    .X(_00974_));
 sg13g2_mux2_1 _10204_ (.A0(\shift_storage.storage [345]),
    .A1(\shift_storage.storage [344]),
    .S(net46),
    .X(_04129_));
 sg13g2_and2_1 _10205_ (.A(net47),
    .B(_04129_),
    .X(_00975_));
 sg13g2_mux2_1 _10206_ (.A0(\shift_storage.storage [346]),
    .A1(\shift_storage.storage [345]),
    .S(net46),
    .X(_04130_));
 sg13g2_and2_1 _10207_ (.A(net47),
    .B(_04130_),
    .X(_00976_));
 sg13g2_mux2_1 _10208_ (.A0(\shift_storage.storage [347]),
    .A1(\shift_storage.storage [346]),
    .S(_04126_),
    .X(_04131_));
 sg13g2_and2_1 _10209_ (.A(net47),
    .B(_04131_),
    .X(_00977_));
 sg13g2_mux2_1 _10210_ (.A0(\shift_storage.storage [348]),
    .A1(\shift_storage.storage [347]),
    .S(_04126_),
    .X(_04132_));
 sg13g2_and2_1 _10211_ (.A(net47),
    .B(_04132_),
    .X(_00978_));
 sg13g2_buf_1 _10212_ (.A(net355),
    .X(_04133_));
 sg13g2_mux2_1 _10213_ (.A0(\shift_storage.storage [349]),
    .A1(\shift_storage.storage [348]),
    .S(net46),
    .X(_04134_));
 sg13g2_and2_1 _10214_ (.A(net45),
    .B(_04134_),
    .X(_00979_));
 sg13g2_mux2_1 _10215_ (.A0(\shift_storage.storage [34]),
    .A1(\shift_storage.storage [33]),
    .S(net46),
    .X(_04135_));
 sg13g2_and2_1 _10216_ (.A(net45),
    .B(_04135_),
    .X(_00980_));
 sg13g2_mux2_1 _10217_ (.A0(\shift_storage.storage [350]),
    .A1(\shift_storage.storage [349]),
    .S(net46),
    .X(_04136_));
 sg13g2_and2_1 _10218_ (.A(net45),
    .B(_04136_),
    .X(_00981_));
 sg13g2_mux2_1 _10219_ (.A0(\shift_storage.storage [351]),
    .A1(\shift_storage.storage [350]),
    .S(net46),
    .X(_04137_));
 sg13g2_and2_1 _10220_ (.A(net45),
    .B(_04137_),
    .X(_00982_));
 sg13g2_buf_1 _10221_ (.A(net356),
    .X(_04138_));
 sg13g2_mux2_1 _10222_ (.A0(\shift_storage.storage [352]),
    .A1(\shift_storage.storage [351]),
    .S(net44),
    .X(_04139_));
 sg13g2_and2_1 _10223_ (.A(net45),
    .B(_04139_),
    .X(_00983_));
 sg13g2_mux2_1 _10224_ (.A0(\shift_storage.storage [353]),
    .A1(\shift_storage.storage [352]),
    .S(net44),
    .X(_04140_));
 sg13g2_and2_1 _10225_ (.A(net45),
    .B(_04140_),
    .X(_00984_));
 sg13g2_mux2_1 _10226_ (.A0(\shift_storage.storage [354]),
    .A1(\shift_storage.storage [353]),
    .S(net44),
    .X(_04141_));
 sg13g2_and2_1 _10227_ (.A(net45),
    .B(_04141_),
    .X(_00985_));
 sg13g2_mux2_1 _10228_ (.A0(\shift_storage.storage [355]),
    .A1(\shift_storage.storage [354]),
    .S(net44),
    .X(_04142_));
 sg13g2_and2_1 _10229_ (.A(net45),
    .B(_04142_),
    .X(_00986_));
 sg13g2_mux2_1 _10230_ (.A0(\shift_storage.storage [356]),
    .A1(\shift_storage.storage [355]),
    .S(net44),
    .X(_04143_));
 sg13g2_and2_1 _10231_ (.A(_04133_),
    .B(_04143_),
    .X(_00987_));
 sg13g2_mux2_1 _10232_ (.A0(\shift_storage.storage [357]),
    .A1(\shift_storage.storage [356]),
    .S(net44),
    .X(_04144_));
 sg13g2_and2_1 _10233_ (.A(_04133_),
    .B(_04144_),
    .X(_00988_));
 sg13g2_buf_1 _10234_ (.A(net355),
    .X(_04145_));
 sg13g2_mux2_1 _10235_ (.A0(\shift_storage.storage [358]),
    .A1(\shift_storage.storage [357]),
    .S(net44),
    .X(_04146_));
 sg13g2_and2_1 _10236_ (.A(net43),
    .B(_04146_),
    .X(_00989_));
 sg13g2_mux2_1 _10237_ (.A0(\shift_storage.storage [359]),
    .A1(\shift_storage.storage [358]),
    .S(_04138_),
    .X(_04147_));
 sg13g2_and2_1 _10238_ (.A(net43),
    .B(_04147_),
    .X(_00990_));
 sg13g2_mux2_1 _10239_ (.A0(\shift_storage.storage [35]),
    .A1(\shift_storage.storage [34]),
    .S(net44),
    .X(_04148_));
 sg13g2_and2_1 _10240_ (.A(net43),
    .B(_04148_),
    .X(_00991_));
 sg13g2_mux2_1 _10241_ (.A0(\shift_storage.storage [360]),
    .A1(\shift_storage.storage [359]),
    .S(_04138_),
    .X(_04149_));
 sg13g2_and2_1 _10242_ (.A(net43),
    .B(_04149_),
    .X(_00992_));
 sg13g2_buf_1 _10243_ (.A(_03058_),
    .X(_04150_));
 sg13g2_buf_1 _10244_ (.A(net409),
    .X(_04151_));
 sg13g2_mux2_1 _10245_ (.A0(\shift_storage.storage [361]),
    .A1(\shift_storage.storage [360]),
    .S(net354),
    .X(_04152_));
 sg13g2_and2_1 _10246_ (.A(net43),
    .B(_04152_),
    .X(_00993_));
 sg13g2_mux2_1 _10247_ (.A0(\shift_storage.storage [362]),
    .A1(\shift_storage.storage [361]),
    .S(net354),
    .X(_04153_));
 sg13g2_and2_1 _10248_ (.A(_04145_),
    .B(_04153_),
    .X(_00994_));
 sg13g2_mux2_1 _10249_ (.A0(\shift_storage.storage [363]),
    .A1(\shift_storage.storage [362]),
    .S(net354),
    .X(_04154_));
 sg13g2_and2_1 _10250_ (.A(_04145_),
    .B(_04154_),
    .X(_00995_));
 sg13g2_mux2_1 _10251_ (.A0(\shift_storage.storage [364]),
    .A1(\shift_storage.storage [363]),
    .S(net354),
    .X(_04155_));
 sg13g2_and2_1 _10252_ (.A(net43),
    .B(_04155_),
    .X(_00996_));
 sg13g2_mux2_1 _10253_ (.A0(\shift_storage.storage [365]),
    .A1(\shift_storage.storage [364]),
    .S(_04151_),
    .X(_04156_));
 sg13g2_and2_1 _10254_ (.A(net43),
    .B(_04156_),
    .X(_00997_));
 sg13g2_mux2_1 _10255_ (.A0(\shift_storage.storage [366]),
    .A1(\shift_storage.storage [365]),
    .S(_04151_),
    .X(_04157_));
 sg13g2_and2_1 _10256_ (.A(net43),
    .B(_04157_),
    .X(_00998_));
 sg13g2_buf_1 _10257_ (.A(_03050_),
    .X(_04158_));
 sg13g2_buf_1 _10258_ (.A(net353),
    .X(_04159_));
 sg13g2_mux2_1 _10259_ (.A0(\shift_storage.storage [367]),
    .A1(\shift_storage.storage [366]),
    .S(net354),
    .X(_04160_));
 sg13g2_and2_1 _10260_ (.A(net42),
    .B(_04160_),
    .X(_00999_));
 sg13g2_mux2_1 _10261_ (.A0(\shift_storage.storage [368]),
    .A1(\shift_storage.storage [367]),
    .S(net354),
    .X(_04161_));
 sg13g2_and2_1 _10262_ (.A(net42),
    .B(_04161_),
    .X(_01000_));
 sg13g2_mux2_1 _10263_ (.A0(\shift_storage.storage [369]),
    .A1(\shift_storage.storage [368]),
    .S(net354),
    .X(_04162_));
 sg13g2_and2_1 _10264_ (.A(net42),
    .B(_04162_),
    .X(_01001_));
 sg13g2_mux2_1 _10265_ (.A0(\shift_storage.storage [36]),
    .A1(\shift_storage.storage [35]),
    .S(net354),
    .X(_04163_));
 sg13g2_and2_1 _10266_ (.A(net42),
    .B(_04163_),
    .X(_01002_));
 sg13g2_buf_1 _10267_ (.A(net409),
    .X(_04164_));
 sg13g2_mux2_1 _10268_ (.A0(\shift_storage.storage [370]),
    .A1(\shift_storage.storage [369]),
    .S(net352),
    .X(_04165_));
 sg13g2_and2_1 _10269_ (.A(net42),
    .B(_04165_),
    .X(_01003_));
 sg13g2_mux2_1 _10270_ (.A0(\shift_storage.storage [371]),
    .A1(\shift_storage.storage [370]),
    .S(net352),
    .X(_04166_));
 sg13g2_and2_1 _10271_ (.A(net42),
    .B(_04166_),
    .X(_01004_));
 sg13g2_mux2_1 _10272_ (.A0(\shift_storage.storage [372]),
    .A1(\shift_storage.storage [371]),
    .S(net352),
    .X(_04167_));
 sg13g2_and2_1 _10273_ (.A(net42),
    .B(_04167_),
    .X(_01005_));
 sg13g2_mux2_1 _10274_ (.A0(\shift_storage.storage [373]),
    .A1(\shift_storage.storage [372]),
    .S(net352),
    .X(_04168_));
 sg13g2_and2_1 _10275_ (.A(net42),
    .B(_04168_),
    .X(_01006_));
 sg13g2_mux2_1 _10276_ (.A0(\shift_storage.storage [374]),
    .A1(\shift_storage.storage [373]),
    .S(net352),
    .X(_04169_));
 sg13g2_and2_1 _10277_ (.A(_04159_),
    .B(_04169_),
    .X(_01007_));
 sg13g2_mux2_1 _10278_ (.A0(\shift_storage.storage [375]),
    .A1(\shift_storage.storage [374]),
    .S(net352),
    .X(_04170_));
 sg13g2_and2_1 _10279_ (.A(_04159_),
    .B(_04170_),
    .X(_01008_));
 sg13g2_buf_1 _10280_ (.A(_04158_),
    .X(_04171_));
 sg13g2_mux2_1 _10281_ (.A0(\shift_storage.storage [376]),
    .A1(\shift_storage.storage [375]),
    .S(net352),
    .X(_04172_));
 sg13g2_and2_1 _10282_ (.A(net41),
    .B(_04172_),
    .X(_01009_));
 sg13g2_mux2_1 _10283_ (.A0(\shift_storage.storage [377]),
    .A1(\shift_storage.storage [376]),
    .S(net352),
    .X(_04173_));
 sg13g2_and2_1 _10284_ (.A(net41),
    .B(_04173_),
    .X(_01010_));
 sg13g2_mux2_1 _10285_ (.A0(\shift_storage.storage [378]),
    .A1(\shift_storage.storage [377]),
    .S(_04164_),
    .X(_04174_));
 sg13g2_and2_1 _10286_ (.A(net41),
    .B(_04174_),
    .X(_01011_));
 sg13g2_mux2_1 _10287_ (.A0(\shift_storage.storage [379]),
    .A1(\shift_storage.storage [378]),
    .S(_04164_),
    .X(_04175_));
 sg13g2_and2_1 _10288_ (.A(_04171_),
    .B(_04175_),
    .X(_01012_));
 sg13g2_buf_1 _10289_ (.A(net409),
    .X(_04176_));
 sg13g2_mux2_1 _10290_ (.A0(\shift_storage.storage [37]),
    .A1(\shift_storage.storage [36]),
    .S(net351),
    .X(_04177_));
 sg13g2_and2_1 _10291_ (.A(net41),
    .B(_04177_),
    .X(_01013_));
 sg13g2_mux2_1 _10292_ (.A0(\shift_storage.storage [380]),
    .A1(\shift_storage.storage [379]),
    .S(net351),
    .X(_04178_));
 sg13g2_and2_1 _10293_ (.A(net41),
    .B(_04178_),
    .X(_01014_));
 sg13g2_mux2_1 _10294_ (.A0(\shift_storage.storage [381]),
    .A1(\shift_storage.storage [380]),
    .S(_04176_),
    .X(_04179_));
 sg13g2_and2_1 _10295_ (.A(net41),
    .B(_04179_),
    .X(_01015_));
 sg13g2_mux2_1 _10296_ (.A0(\shift_storage.storage [382]),
    .A1(\shift_storage.storage [381]),
    .S(_04176_),
    .X(_04180_));
 sg13g2_and2_1 _10297_ (.A(net41),
    .B(_04180_),
    .X(_01016_));
 sg13g2_mux2_1 _10298_ (.A0(\shift_storage.storage [383]),
    .A1(\shift_storage.storage [382]),
    .S(net351),
    .X(_04181_));
 sg13g2_and2_1 _10299_ (.A(_04171_),
    .B(_04181_),
    .X(_01017_));
 sg13g2_mux2_1 _10300_ (.A0(\shift_storage.storage [384]),
    .A1(\shift_storage.storage [383]),
    .S(net351),
    .X(_04182_));
 sg13g2_and2_1 _10301_ (.A(net41),
    .B(_04182_),
    .X(_01018_));
 sg13g2_buf_1 _10302_ (.A(_04158_),
    .X(_04183_));
 sg13g2_mux2_1 _10303_ (.A0(\shift_storage.storage [385]),
    .A1(\shift_storage.storage [384]),
    .S(net351),
    .X(_04184_));
 sg13g2_and2_1 _10304_ (.A(net40),
    .B(_04184_),
    .X(_01019_));
 sg13g2_mux2_1 _10305_ (.A0(\shift_storage.storage [386]),
    .A1(\shift_storage.storage [385]),
    .S(net351),
    .X(_04185_));
 sg13g2_and2_1 _10306_ (.A(net40),
    .B(_04185_),
    .X(_01020_));
 sg13g2_mux2_1 _10307_ (.A0(\shift_storage.storage [387]),
    .A1(\shift_storage.storage [386]),
    .S(net351),
    .X(_04186_));
 sg13g2_and2_1 _10308_ (.A(net40),
    .B(_04186_),
    .X(_01021_));
 sg13g2_mux2_1 _10309_ (.A0(\shift_storage.storage [388]),
    .A1(\shift_storage.storage [387]),
    .S(net351),
    .X(_04187_));
 sg13g2_and2_1 _10310_ (.A(_04183_),
    .B(_04187_),
    .X(_01022_));
 sg13g2_buf_1 _10311_ (.A(_04150_),
    .X(_04188_));
 sg13g2_mux2_1 _10312_ (.A0(\shift_storage.storage [389]),
    .A1(\shift_storage.storage [388]),
    .S(_04188_),
    .X(_04189_));
 sg13g2_and2_1 _10313_ (.A(net40),
    .B(_04189_),
    .X(_01023_));
 sg13g2_mux2_1 _10314_ (.A0(\shift_storage.storage [38]),
    .A1(\shift_storage.storage [37]),
    .S(_04188_),
    .X(_04190_));
 sg13g2_and2_1 _10315_ (.A(_04183_),
    .B(_04190_),
    .X(_01024_));
 sg13g2_mux2_1 _10316_ (.A0(\shift_storage.storage [390]),
    .A1(\shift_storage.storage [389]),
    .S(net350),
    .X(_04191_));
 sg13g2_and2_1 _10317_ (.A(net40),
    .B(_04191_),
    .X(_01025_));
 sg13g2_mux2_1 _10318_ (.A0(\shift_storage.storage [391]),
    .A1(\shift_storage.storage [390]),
    .S(net350),
    .X(_04192_));
 sg13g2_and2_1 _10319_ (.A(net40),
    .B(_04192_),
    .X(_01026_));
 sg13g2_mux2_1 _10320_ (.A0(\shift_storage.storage [392]),
    .A1(\shift_storage.storage [391]),
    .S(net350),
    .X(_04193_));
 sg13g2_and2_1 _10321_ (.A(net40),
    .B(_04193_),
    .X(_01027_));
 sg13g2_mux2_1 _10322_ (.A0(\shift_storage.storage [393]),
    .A1(\shift_storage.storage [392]),
    .S(net350),
    .X(_04194_));
 sg13g2_and2_1 _10323_ (.A(net40),
    .B(_04194_),
    .X(_01028_));
 sg13g2_buf_1 _10324_ (.A(net353),
    .X(_04195_));
 sg13g2_mux2_1 _10325_ (.A0(\shift_storage.storage [394]),
    .A1(\shift_storage.storage [393]),
    .S(net350),
    .X(_04196_));
 sg13g2_and2_1 _10326_ (.A(net39),
    .B(_04196_),
    .X(_01029_));
 sg13g2_mux2_1 _10327_ (.A0(\shift_storage.storage [395]),
    .A1(\shift_storage.storage [394]),
    .S(net350),
    .X(_04197_));
 sg13g2_and2_1 _10328_ (.A(net39),
    .B(_04197_),
    .X(_01030_));
 sg13g2_mux2_1 _10329_ (.A0(\shift_storage.storage [396]),
    .A1(\shift_storage.storage [395]),
    .S(net350),
    .X(_04198_));
 sg13g2_and2_1 _10330_ (.A(net39),
    .B(_04198_),
    .X(_01031_));
 sg13g2_mux2_1 _10331_ (.A0(\shift_storage.storage [397]),
    .A1(\shift_storage.storage [396]),
    .S(net350),
    .X(_04199_));
 sg13g2_and2_1 _10332_ (.A(net39),
    .B(_04199_),
    .X(_01032_));
 sg13g2_buf_1 _10333_ (.A(_04150_),
    .X(_04200_));
 sg13g2_mux2_1 _10334_ (.A0(\shift_storage.storage [398]),
    .A1(\shift_storage.storage [397]),
    .S(net349),
    .X(_04201_));
 sg13g2_and2_1 _10335_ (.A(net39),
    .B(_04201_),
    .X(_01033_));
 sg13g2_mux2_1 _10336_ (.A0(\shift_storage.storage [399]),
    .A1(\shift_storage.storage [398]),
    .S(net349),
    .X(_04202_));
 sg13g2_and2_1 _10337_ (.A(net39),
    .B(_04202_),
    .X(_01034_));
 sg13g2_mux2_1 _10338_ (.A0(\shift_storage.storage [39]),
    .A1(\shift_storage.storage [38]),
    .S(net349),
    .X(_04203_));
 sg13g2_and2_1 _10339_ (.A(net39),
    .B(_04203_),
    .X(_01035_));
 sg13g2_mux2_1 _10340_ (.A0(\shift_storage.storage [3]),
    .A1(\shift_storage.storage [2]),
    .S(net349),
    .X(_04204_));
 sg13g2_and2_1 _10341_ (.A(net39),
    .B(_04204_),
    .X(_01036_));
 sg13g2_mux2_1 _10342_ (.A0(\shift_storage.storage [400]),
    .A1(\shift_storage.storage [399]),
    .S(net349),
    .X(_04205_));
 sg13g2_and2_1 _10343_ (.A(_04195_),
    .B(_04205_),
    .X(_01037_));
 sg13g2_mux2_1 _10344_ (.A0(\shift_storage.storage [401]),
    .A1(\shift_storage.storage [400]),
    .S(net349),
    .X(_04206_));
 sg13g2_and2_1 _10345_ (.A(_04195_),
    .B(_04206_),
    .X(_01038_));
 sg13g2_buf_1 _10346_ (.A(net353),
    .X(_04207_));
 sg13g2_mux2_1 _10347_ (.A0(\shift_storage.storage [402]),
    .A1(\shift_storage.storage [401]),
    .S(net349),
    .X(_04208_));
 sg13g2_and2_1 _10348_ (.A(net38),
    .B(_04208_),
    .X(_01039_));
 sg13g2_mux2_1 _10349_ (.A0(\shift_storage.storage [403]),
    .A1(\shift_storage.storage [402]),
    .S(net349),
    .X(_04209_));
 sg13g2_and2_1 _10350_ (.A(net38),
    .B(_04209_),
    .X(_01040_));
 sg13g2_mux2_1 _10351_ (.A0(\shift_storage.storage [404]),
    .A1(\shift_storage.storage [403]),
    .S(_04200_),
    .X(_04210_));
 sg13g2_and2_1 _10352_ (.A(net38),
    .B(_04210_),
    .X(_01041_));
 sg13g2_mux2_1 _10353_ (.A0(\shift_storage.storage [405]),
    .A1(\shift_storage.storage [404]),
    .S(_04200_),
    .X(_04211_));
 sg13g2_and2_1 _10354_ (.A(_04207_),
    .B(_04211_),
    .X(_01042_));
 sg13g2_buf_1 _10355_ (.A(net409),
    .X(_04212_));
 sg13g2_mux2_1 _10356_ (.A0(\shift_storage.storage [406]),
    .A1(\shift_storage.storage [405]),
    .S(net348),
    .X(_04213_));
 sg13g2_and2_1 _10357_ (.A(net38),
    .B(_04213_),
    .X(_01043_));
 sg13g2_mux2_1 _10358_ (.A0(\shift_storage.storage [407]),
    .A1(\shift_storage.storage [406]),
    .S(net348),
    .X(_04214_));
 sg13g2_and2_1 _10359_ (.A(net38),
    .B(_04214_),
    .X(_01044_));
 sg13g2_mux2_1 _10360_ (.A0(\shift_storage.storage [408]),
    .A1(\shift_storage.storage [407]),
    .S(net348),
    .X(_04215_));
 sg13g2_and2_1 _10361_ (.A(net38),
    .B(_04215_),
    .X(_01045_));
 sg13g2_mux2_1 _10362_ (.A0(\shift_storage.storage [409]),
    .A1(\shift_storage.storage [408]),
    .S(net348),
    .X(_04216_));
 sg13g2_and2_1 _10363_ (.A(net38),
    .B(_04216_),
    .X(_01046_));
 sg13g2_mux2_1 _10364_ (.A0(\shift_storage.storage [40]),
    .A1(\shift_storage.storage [39]),
    .S(net348),
    .X(_04217_));
 sg13g2_and2_1 _10365_ (.A(_04207_),
    .B(_04217_),
    .X(_01047_));
 sg13g2_mux2_1 _10366_ (.A0(\shift_storage.storage [410]),
    .A1(\shift_storage.storage [409]),
    .S(net348),
    .X(_04218_));
 sg13g2_and2_1 _10367_ (.A(net38),
    .B(_04218_),
    .X(_01048_));
 sg13g2_buf_1 _10368_ (.A(net353),
    .X(_04219_));
 sg13g2_mux2_1 _10369_ (.A0(\shift_storage.storage [411]),
    .A1(\shift_storage.storage [410]),
    .S(net348),
    .X(_04220_));
 sg13g2_and2_1 _10370_ (.A(net37),
    .B(_04220_),
    .X(_01049_));
 sg13g2_mux2_1 _10371_ (.A0(\shift_storage.storage [412]),
    .A1(\shift_storage.storage [411]),
    .S(net348),
    .X(_04221_));
 sg13g2_and2_1 _10372_ (.A(net37),
    .B(_04221_),
    .X(_01050_));
 sg13g2_mux2_1 _10373_ (.A0(\shift_storage.storage [413]),
    .A1(\shift_storage.storage [412]),
    .S(_04212_),
    .X(_04222_));
 sg13g2_and2_1 _10374_ (.A(net37),
    .B(_04222_),
    .X(_01051_));
 sg13g2_mux2_1 _10375_ (.A0(\shift_storage.storage [414]),
    .A1(\shift_storage.storage [413]),
    .S(_04212_),
    .X(_04223_));
 sg13g2_and2_1 _10376_ (.A(net37),
    .B(_04223_),
    .X(_01052_));
 sg13g2_buf_1 _10377_ (.A(net409),
    .X(_04224_));
 sg13g2_mux2_1 _10378_ (.A0(\shift_storage.storage [415]),
    .A1(\shift_storage.storage [414]),
    .S(net347),
    .X(_04225_));
 sg13g2_and2_1 _10379_ (.A(net37),
    .B(_04225_),
    .X(_01053_));
 sg13g2_mux2_1 _10380_ (.A0(\shift_storage.storage [416]),
    .A1(\shift_storage.storage [415]),
    .S(net347),
    .X(_04226_));
 sg13g2_and2_1 _10381_ (.A(net37),
    .B(_04226_),
    .X(_01054_));
 sg13g2_mux2_1 _10382_ (.A0(\shift_storage.storage [417]),
    .A1(\shift_storage.storage [416]),
    .S(net347),
    .X(_04227_));
 sg13g2_and2_1 _10383_ (.A(net37),
    .B(_04227_),
    .X(_01055_));
 sg13g2_mux2_1 _10384_ (.A0(\shift_storage.storage [418]),
    .A1(\shift_storage.storage [417]),
    .S(net347),
    .X(_04228_));
 sg13g2_and2_1 _10385_ (.A(_04219_),
    .B(_04228_),
    .X(_01056_));
 sg13g2_mux2_1 _10386_ (.A0(\shift_storage.storage [419]),
    .A1(\shift_storage.storage [418]),
    .S(net347),
    .X(_04229_));
 sg13g2_and2_1 _10387_ (.A(_04219_),
    .B(_04229_),
    .X(_01057_));
 sg13g2_mux2_1 _10388_ (.A0(\shift_storage.storage [41]),
    .A1(\shift_storage.storage [40]),
    .S(net347),
    .X(_04230_));
 sg13g2_and2_1 _10389_ (.A(net37),
    .B(_04230_),
    .X(_01058_));
 sg13g2_buf_1 _10390_ (.A(net353),
    .X(_04231_));
 sg13g2_mux2_1 _10391_ (.A0(\shift_storage.storage [420]),
    .A1(\shift_storage.storage [419]),
    .S(net347),
    .X(_04232_));
 sg13g2_and2_1 _10392_ (.A(net36),
    .B(_04232_),
    .X(_01059_));
 sg13g2_mux2_1 _10393_ (.A0(\shift_storage.storage [421]),
    .A1(\shift_storage.storage [420]),
    .S(net347),
    .X(_04233_));
 sg13g2_and2_1 _10394_ (.A(net36),
    .B(_04233_),
    .X(_01060_));
 sg13g2_mux2_1 _10395_ (.A0(\shift_storage.storage [422]),
    .A1(\shift_storage.storage [421]),
    .S(_04224_),
    .X(_04234_));
 sg13g2_and2_1 _10396_ (.A(net36),
    .B(_04234_),
    .X(_01061_));
 sg13g2_mux2_1 _10397_ (.A0(\shift_storage.storage [423]),
    .A1(\shift_storage.storage [422]),
    .S(_04224_),
    .X(_04235_));
 sg13g2_and2_1 _10398_ (.A(net36),
    .B(_04235_),
    .X(_01062_));
 sg13g2_buf_1 _10399_ (.A(net409),
    .X(_04236_));
 sg13g2_mux2_1 _10400_ (.A0(\shift_storage.storage [424]),
    .A1(\shift_storage.storage [423]),
    .S(net346),
    .X(_04237_));
 sg13g2_and2_1 _10401_ (.A(net36),
    .B(_04237_),
    .X(_01063_));
 sg13g2_mux2_1 _10402_ (.A0(\shift_storage.storage [425]),
    .A1(\shift_storage.storage [424]),
    .S(net346),
    .X(_04238_));
 sg13g2_and2_1 _10403_ (.A(net36),
    .B(_04238_),
    .X(_01064_));
 sg13g2_mux2_1 _10404_ (.A0(\shift_storage.storage [426]),
    .A1(\shift_storage.storage [425]),
    .S(net346),
    .X(_04239_));
 sg13g2_and2_1 _10405_ (.A(net36),
    .B(_04239_),
    .X(_01065_));
 sg13g2_mux2_1 _10406_ (.A0(\shift_storage.storage [427]),
    .A1(\shift_storage.storage [426]),
    .S(net346),
    .X(_04240_));
 sg13g2_and2_1 _10407_ (.A(_04231_),
    .B(_04240_),
    .X(_01066_));
 sg13g2_mux2_1 _10408_ (.A0(\shift_storage.storage [428]),
    .A1(\shift_storage.storage [427]),
    .S(_04236_),
    .X(_04241_));
 sg13g2_and2_1 _10409_ (.A(_04231_),
    .B(_04241_),
    .X(_01067_));
 sg13g2_mux2_1 _10410_ (.A0(\shift_storage.storage [429]),
    .A1(\shift_storage.storage [428]),
    .S(_04236_),
    .X(_04242_));
 sg13g2_and2_1 _10411_ (.A(net36),
    .B(_04242_),
    .X(_01068_));
 sg13g2_buf_1 _10412_ (.A(net353),
    .X(_04243_));
 sg13g2_mux2_1 _10413_ (.A0(\shift_storage.storage [42]),
    .A1(\shift_storage.storage [41]),
    .S(net346),
    .X(_04244_));
 sg13g2_and2_1 _10414_ (.A(net35),
    .B(_04244_),
    .X(_01069_));
 sg13g2_mux2_1 _10415_ (.A0(\shift_storage.storage [430]),
    .A1(\shift_storage.storage [429]),
    .S(net346),
    .X(_04245_));
 sg13g2_and2_1 _10416_ (.A(net35),
    .B(_04245_),
    .X(_01070_));
 sg13g2_mux2_1 _10417_ (.A0(\shift_storage.storage [431]),
    .A1(\shift_storage.storage [430]),
    .S(net346),
    .X(_04246_));
 sg13g2_and2_1 _10418_ (.A(net35),
    .B(_04246_),
    .X(_01071_));
 sg13g2_mux2_1 _10419_ (.A0(\shift_storage.storage [432]),
    .A1(\shift_storage.storage [431]),
    .S(net346),
    .X(_04247_));
 sg13g2_and2_1 _10420_ (.A(net35),
    .B(_04247_),
    .X(_01072_));
 sg13g2_buf_1 _10421_ (.A(net409),
    .X(_04248_));
 sg13g2_mux2_1 _10422_ (.A0(\shift_storage.storage [433]),
    .A1(\shift_storage.storage [432]),
    .S(net345),
    .X(_04249_));
 sg13g2_and2_1 _10423_ (.A(net35),
    .B(_04249_),
    .X(_01073_));
 sg13g2_mux2_1 _10424_ (.A0(\shift_storage.storage [434]),
    .A1(\shift_storage.storage [433]),
    .S(net345),
    .X(_04250_));
 sg13g2_and2_1 _10425_ (.A(net35),
    .B(_04250_),
    .X(_01074_));
 sg13g2_mux2_1 _10426_ (.A0(\shift_storage.storage [435]),
    .A1(\shift_storage.storage [434]),
    .S(net345),
    .X(_04251_));
 sg13g2_and2_1 _10427_ (.A(net35),
    .B(_04251_),
    .X(_01075_));
 sg13g2_mux2_1 _10428_ (.A0(\shift_storage.storage [436]),
    .A1(\shift_storage.storage [435]),
    .S(net345),
    .X(_04252_));
 sg13g2_and2_1 _10429_ (.A(net35),
    .B(_04252_),
    .X(_01076_));
 sg13g2_mux2_1 _10430_ (.A0(\shift_storage.storage [437]),
    .A1(\shift_storage.storage [436]),
    .S(net345),
    .X(_04253_));
 sg13g2_and2_1 _10431_ (.A(_04243_),
    .B(_04253_),
    .X(_01077_));
 sg13g2_mux2_1 _10432_ (.A0(\shift_storage.storage [438]),
    .A1(\shift_storage.storage [437]),
    .S(net345),
    .X(_04254_));
 sg13g2_and2_1 _10433_ (.A(_04243_),
    .B(_04254_),
    .X(_01078_));
 sg13g2_buf_1 _10434_ (.A(net353),
    .X(_04255_));
 sg13g2_mux2_1 _10435_ (.A0(\shift_storage.storage [439]),
    .A1(\shift_storage.storage [438]),
    .S(net345),
    .X(_04256_));
 sg13g2_and2_1 _10436_ (.A(net34),
    .B(_04256_),
    .X(_01079_));
 sg13g2_mux2_1 _10437_ (.A0(\shift_storage.storage [43]),
    .A1(\shift_storage.storage [42]),
    .S(net345),
    .X(_04257_));
 sg13g2_and2_1 _10438_ (.A(net34),
    .B(_04257_),
    .X(_01080_));
 sg13g2_mux2_1 _10439_ (.A0(\shift_storage.storage [440]),
    .A1(\shift_storage.storage [439]),
    .S(_04248_),
    .X(_04258_));
 sg13g2_and2_1 _10440_ (.A(net34),
    .B(_04258_),
    .X(_01081_));
 sg13g2_mux2_1 _10441_ (.A0(\shift_storage.storage [441]),
    .A1(\shift_storage.storage [440]),
    .S(_04248_),
    .X(_04259_));
 sg13g2_and2_1 _10442_ (.A(net34),
    .B(_04259_),
    .X(_01082_));
 sg13g2_buf_1 _10443_ (.A(net409),
    .X(_04260_));
 sg13g2_mux2_1 _10444_ (.A0(\shift_storage.storage [442]),
    .A1(\shift_storage.storage [441]),
    .S(net344),
    .X(_04261_));
 sg13g2_and2_1 _10445_ (.A(net34),
    .B(_04261_),
    .X(_01083_));
 sg13g2_mux2_1 _10446_ (.A0(\shift_storage.storage [443]),
    .A1(\shift_storage.storage [442]),
    .S(net344),
    .X(_04262_));
 sg13g2_and2_1 _10447_ (.A(_04255_),
    .B(_04262_),
    .X(_01084_));
 sg13g2_mux2_1 _10448_ (.A0(\shift_storage.storage [444]),
    .A1(\shift_storage.storage [443]),
    .S(net344),
    .X(_04263_));
 sg13g2_and2_1 _10449_ (.A(_04255_),
    .B(_04263_),
    .X(_01085_));
 sg13g2_mux2_1 _10450_ (.A0(\shift_storage.storage [445]),
    .A1(\shift_storage.storage [444]),
    .S(_04260_),
    .X(_04264_));
 sg13g2_and2_1 _10451_ (.A(net34),
    .B(_04264_),
    .X(_01086_));
 sg13g2_mux2_1 _10452_ (.A0(\shift_storage.storage [446]),
    .A1(\shift_storage.storage [445]),
    .S(_04260_),
    .X(_04265_));
 sg13g2_and2_1 _10453_ (.A(net34),
    .B(_04265_),
    .X(_01087_));
 sg13g2_mux2_1 _10454_ (.A0(\shift_storage.storage [447]),
    .A1(\shift_storage.storage [446]),
    .S(net344),
    .X(_04266_));
 sg13g2_and2_1 _10455_ (.A(net34),
    .B(_04266_),
    .X(_01088_));
 sg13g2_buf_1 _10456_ (.A(net353),
    .X(_04267_));
 sg13g2_mux2_1 _10457_ (.A0(\shift_storage.storage [448]),
    .A1(\shift_storage.storage [447]),
    .S(net344),
    .X(_04268_));
 sg13g2_and2_1 _10458_ (.A(net33),
    .B(_04268_),
    .X(_01089_));
 sg13g2_mux2_1 _10459_ (.A0(\shift_storage.storage [449]),
    .A1(\shift_storage.storage [448]),
    .S(net344),
    .X(_04269_));
 sg13g2_and2_1 _10460_ (.A(net33),
    .B(_04269_),
    .X(_01090_));
 sg13g2_mux2_1 _10461_ (.A0(\shift_storage.storage [44]),
    .A1(\shift_storage.storage [43]),
    .S(net344),
    .X(_04270_));
 sg13g2_and2_1 _10462_ (.A(_04267_),
    .B(_04270_),
    .X(_01091_));
 sg13g2_mux2_1 _10463_ (.A0(\shift_storage.storage [450]),
    .A1(\shift_storage.storage [449]),
    .S(net344),
    .X(_04271_));
 sg13g2_and2_1 _10464_ (.A(_04267_),
    .B(_04271_),
    .X(_01092_));
 sg13g2_buf_1 _10465_ (.A(_03058_),
    .X(_04272_));
 sg13g2_buf_1 _10466_ (.A(net408),
    .X(_04273_));
 sg13g2_mux2_1 _10467_ (.A0(\shift_storage.storage [451]),
    .A1(\shift_storage.storage [450]),
    .S(net343),
    .X(_04274_));
 sg13g2_and2_1 _10468_ (.A(net33),
    .B(_04274_),
    .X(_01093_));
 sg13g2_mux2_1 _10469_ (.A0(\shift_storage.storage [452]),
    .A1(\shift_storage.storage [451]),
    .S(net343),
    .X(_04275_));
 sg13g2_and2_1 _10470_ (.A(net33),
    .B(_04275_),
    .X(_01094_));
 sg13g2_mux2_1 _10471_ (.A0(\shift_storage.storage [453]),
    .A1(\shift_storage.storage [452]),
    .S(net343),
    .X(_04276_));
 sg13g2_and2_1 _10472_ (.A(net33),
    .B(_04276_),
    .X(_01095_));
 sg13g2_mux2_1 _10473_ (.A0(\shift_storage.storage [454]),
    .A1(\shift_storage.storage [453]),
    .S(_04273_),
    .X(_04277_));
 sg13g2_and2_1 _10474_ (.A(net33),
    .B(_04277_),
    .X(_01096_));
 sg13g2_mux2_1 _10475_ (.A0(\shift_storage.storage [455]),
    .A1(\shift_storage.storage [454]),
    .S(_04273_),
    .X(_04278_));
 sg13g2_and2_1 _10476_ (.A(net33),
    .B(_04278_),
    .X(_01097_));
 sg13g2_mux2_1 _10477_ (.A0(\shift_storage.storage [456]),
    .A1(\shift_storage.storage [455]),
    .S(net343),
    .X(_04279_));
 sg13g2_and2_1 _10478_ (.A(net33),
    .B(_04279_),
    .X(_01098_));
 sg13g2_buf_1 _10479_ (.A(_02909_),
    .X(_04280_));
 sg13g2_buf_1 _10480_ (.A(net407),
    .X(_04281_));
 sg13g2_mux2_1 _10481_ (.A0(\shift_storage.storage [457]),
    .A1(\shift_storage.storage [456]),
    .S(net343),
    .X(_04282_));
 sg13g2_and2_1 _10482_ (.A(net342),
    .B(_04282_),
    .X(_01099_));
 sg13g2_mux2_1 _10483_ (.A0(\shift_storage.storage [458]),
    .A1(\shift_storage.storage [457]),
    .S(net343),
    .X(_04283_));
 sg13g2_and2_1 _10484_ (.A(net342),
    .B(_04283_),
    .X(_01100_));
 sg13g2_mux2_1 _10485_ (.A0(\shift_storage.storage [459]),
    .A1(\shift_storage.storage [458]),
    .S(net343),
    .X(_04284_));
 sg13g2_and2_1 _10486_ (.A(_04281_),
    .B(_04284_),
    .X(_01101_));
 sg13g2_mux2_1 _10487_ (.A0(\shift_storage.storage [45]),
    .A1(\shift_storage.storage [44]),
    .S(net343),
    .X(_04285_));
 sg13g2_and2_1 _10488_ (.A(_04281_),
    .B(_04285_),
    .X(_01102_));
 sg13g2_buf_1 _10489_ (.A(net408),
    .X(_04286_));
 sg13g2_mux2_1 _10490_ (.A0(\shift_storage.storage [460]),
    .A1(\shift_storage.storage [459]),
    .S(net341),
    .X(_04287_));
 sg13g2_and2_1 _10491_ (.A(net342),
    .B(_04287_),
    .X(_01103_));
 sg13g2_mux2_1 _10492_ (.A0(\shift_storage.storage [461]),
    .A1(\shift_storage.storage [460]),
    .S(net341),
    .X(_04288_));
 sg13g2_and2_1 _10493_ (.A(net342),
    .B(_04288_),
    .X(_01104_));
 sg13g2_mux2_1 _10494_ (.A0(\shift_storage.storage [462]),
    .A1(\shift_storage.storage [461]),
    .S(net341),
    .X(_04289_));
 sg13g2_and2_1 _10495_ (.A(net342),
    .B(_04289_),
    .X(_01105_));
 sg13g2_mux2_1 _10496_ (.A0(\shift_storage.storage [463]),
    .A1(\shift_storage.storage [462]),
    .S(net341),
    .X(_04290_));
 sg13g2_and2_1 _10497_ (.A(net342),
    .B(_04290_),
    .X(_01106_));
 sg13g2_mux2_1 _10498_ (.A0(\shift_storage.storage [464]),
    .A1(\shift_storage.storage [463]),
    .S(_04286_),
    .X(_04291_));
 sg13g2_and2_1 _10499_ (.A(net342),
    .B(_04291_),
    .X(_01107_));
 sg13g2_mux2_1 _10500_ (.A0(\shift_storage.storage [465]),
    .A1(\shift_storage.storage [464]),
    .S(_04286_),
    .X(_04292_));
 sg13g2_and2_1 _10501_ (.A(net342),
    .B(_04292_),
    .X(_01108_));
 sg13g2_buf_1 _10502_ (.A(net407),
    .X(_04293_));
 sg13g2_mux2_1 _10503_ (.A0(\shift_storage.storage [466]),
    .A1(\shift_storage.storage [465]),
    .S(net341),
    .X(_04294_));
 sg13g2_and2_1 _10504_ (.A(net340),
    .B(_04294_),
    .X(_01109_));
 sg13g2_mux2_1 _10505_ (.A0(\shift_storage.storage [467]),
    .A1(\shift_storage.storage [466]),
    .S(net341),
    .X(_04295_));
 sg13g2_and2_1 _10506_ (.A(net340),
    .B(_04295_),
    .X(_01110_));
 sg13g2_mux2_1 _10507_ (.A0(\shift_storage.storage [468]),
    .A1(\shift_storage.storage [467]),
    .S(net341),
    .X(_04296_));
 sg13g2_and2_1 _10508_ (.A(_04293_),
    .B(_04296_),
    .X(_01111_));
 sg13g2_mux2_1 _10509_ (.A0(\shift_storage.storage [469]),
    .A1(\shift_storage.storage [468]),
    .S(net341),
    .X(_04297_));
 sg13g2_and2_1 _10510_ (.A(_04293_),
    .B(_04297_),
    .X(_01112_));
 sg13g2_buf_1 _10511_ (.A(_04272_),
    .X(_04298_));
 sg13g2_mux2_1 _10512_ (.A0(\shift_storage.storage [46]),
    .A1(\shift_storage.storage [45]),
    .S(net339),
    .X(_04299_));
 sg13g2_and2_1 _10513_ (.A(net340),
    .B(_04299_),
    .X(_01113_));
 sg13g2_mux2_1 _10514_ (.A0(\shift_storage.storage [470]),
    .A1(\shift_storage.storage [469]),
    .S(net339),
    .X(_04300_));
 sg13g2_and2_1 _10515_ (.A(net340),
    .B(_04300_),
    .X(_01114_));
 sg13g2_mux2_1 _10516_ (.A0(\shift_storage.storage [471]),
    .A1(\shift_storage.storage [470]),
    .S(net339),
    .X(_04301_));
 sg13g2_and2_1 _10517_ (.A(net340),
    .B(_04301_),
    .X(_01115_));
 sg13g2_mux2_1 _10518_ (.A0(\shift_storage.storage [472]),
    .A1(\shift_storage.storage [471]),
    .S(net339),
    .X(_04302_));
 sg13g2_and2_1 _10519_ (.A(net340),
    .B(_04302_),
    .X(_01116_));
 sg13g2_mux2_1 _10520_ (.A0(\shift_storage.storage [473]),
    .A1(\shift_storage.storage [472]),
    .S(net339),
    .X(_04303_));
 sg13g2_and2_1 _10521_ (.A(net340),
    .B(_04303_),
    .X(_01117_));
 sg13g2_mux2_1 _10522_ (.A0(\shift_storage.storage [474]),
    .A1(\shift_storage.storage [473]),
    .S(net339),
    .X(_04304_));
 sg13g2_and2_1 _10523_ (.A(net340),
    .B(_04304_),
    .X(_01118_));
 sg13g2_buf_1 _10524_ (.A(_04280_),
    .X(_04305_));
 sg13g2_mux2_1 _10525_ (.A0(\shift_storage.storage [475]),
    .A1(\shift_storage.storage [474]),
    .S(net339),
    .X(_04306_));
 sg13g2_and2_1 _10526_ (.A(net338),
    .B(_04306_),
    .X(_01119_));
 sg13g2_mux2_1 _10527_ (.A0(\shift_storage.storage [476]),
    .A1(\shift_storage.storage [475]),
    .S(net339),
    .X(_04307_));
 sg13g2_and2_1 _10528_ (.A(net338),
    .B(_04307_),
    .X(_01120_));
 sg13g2_mux2_1 _10529_ (.A0(\shift_storage.storage [477]),
    .A1(\shift_storage.storage [476]),
    .S(_04298_),
    .X(_04308_));
 sg13g2_and2_1 _10530_ (.A(net338),
    .B(_04308_),
    .X(_01121_));
 sg13g2_mux2_1 _10531_ (.A0(\shift_storage.storage [478]),
    .A1(\shift_storage.storage [477]),
    .S(_04298_),
    .X(_04309_));
 sg13g2_and2_1 _10532_ (.A(net338),
    .B(_04309_),
    .X(_01122_));
 sg13g2_buf_1 _10533_ (.A(_04272_),
    .X(_04310_));
 sg13g2_mux2_1 _10534_ (.A0(\shift_storage.storage [479]),
    .A1(\shift_storage.storage [478]),
    .S(net337),
    .X(_04311_));
 sg13g2_and2_1 _10535_ (.A(net338),
    .B(_04311_),
    .X(_01123_));
 sg13g2_mux2_1 _10536_ (.A0(\shift_storage.storage [47]),
    .A1(\shift_storage.storage [46]),
    .S(net337),
    .X(_04312_));
 sg13g2_and2_1 _10537_ (.A(net338),
    .B(_04312_),
    .X(_01124_));
 sg13g2_mux2_1 _10538_ (.A0(\shift_storage.storage [480]),
    .A1(\shift_storage.storage [479]),
    .S(net337),
    .X(_04313_));
 sg13g2_and2_1 _10539_ (.A(net338),
    .B(_04313_),
    .X(_01125_));
 sg13g2_mux2_1 _10540_ (.A0(\shift_storage.storage [481]),
    .A1(\shift_storage.storage [480]),
    .S(net337),
    .X(_04314_));
 sg13g2_and2_1 _10541_ (.A(net338),
    .B(_04314_),
    .X(_01126_));
 sg13g2_mux2_1 _10542_ (.A0(\shift_storage.storage [482]),
    .A1(\shift_storage.storage [481]),
    .S(_04310_),
    .X(_04315_));
 sg13g2_and2_1 _10543_ (.A(_04305_),
    .B(_04315_),
    .X(_01127_));
 sg13g2_mux2_1 _10544_ (.A0(\shift_storage.storage [483]),
    .A1(\shift_storage.storage [482]),
    .S(_04310_),
    .X(_04316_));
 sg13g2_and2_1 _10545_ (.A(_04305_),
    .B(_04316_),
    .X(_01128_));
 sg13g2_buf_1 _10546_ (.A(_04280_),
    .X(_04317_));
 sg13g2_mux2_1 _10547_ (.A0(\shift_storage.storage [484]),
    .A1(\shift_storage.storage [483]),
    .S(net337),
    .X(_04318_));
 sg13g2_and2_1 _10548_ (.A(net336),
    .B(_04318_),
    .X(_01129_));
 sg13g2_mux2_1 _10549_ (.A0(\shift_storage.storage [485]),
    .A1(\shift_storage.storage [484]),
    .S(net337),
    .X(_04319_));
 sg13g2_and2_1 _10550_ (.A(net336),
    .B(_04319_),
    .X(_01130_));
 sg13g2_mux2_1 _10551_ (.A0(\shift_storage.storage [486]),
    .A1(\shift_storage.storage [485]),
    .S(net337),
    .X(_04320_));
 sg13g2_and2_1 _10552_ (.A(net336),
    .B(_04320_),
    .X(_01131_));
 sg13g2_mux2_1 _10553_ (.A0(\shift_storage.storage [487]),
    .A1(\shift_storage.storage [486]),
    .S(net337),
    .X(_04321_));
 sg13g2_and2_1 _10554_ (.A(net336),
    .B(_04321_),
    .X(_01132_));
 sg13g2_buf_1 _10555_ (.A(net408),
    .X(_04322_));
 sg13g2_mux2_1 _10556_ (.A0(\shift_storage.storage [488]),
    .A1(\shift_storage.storage [487]),
    .S(net335),
    .X(_04323_));
 sg13g2_and2_1 _10557_ (.A(net336),
    .B(_04323_),
    .X(_01133_));
 sg13g2_mux2_1 _10558_ (.A0(\shift_storage.storage [489]),
    .A1(\shift_storage.storage [488]),
    .S(net335),
    .X(_04324_));
 sg13g2_and2_1 _10559_ (.A(net336),
    .B(_04324_),
    .X(_01134_));
 sg13g2_mux2_1 _10560_ (.A0(\shift_storage.storage [48]),
    .A1(\shift_storage.storage [47]),
    .S(_04322_),
    .X(_04325_));
 sg13g2_and2_1 _10561_ (.A(net336),
    .B(_04325_),
    .X(_01135_));
 sg13g2_mux2_1 _10562_ (.A0(\shift_storage.storage [490]),
    .A1(\shift_storage.storage [489]),
    .S(net335),
    .X(_04326_));
 sg13g2_and2_1 _10563_ (.A(net336),
    .B(_04326_),
    .X(_01136_));
 sg13g2_mux2_1 _10564_ (.A0(\shift_storage.storage [491]),
    .A1(\shift_storage.storage [490]),
    .S(net335),
    .X(_04327_));
 sg13g2_and2_1 _10565_ (.A(_04317_),
    .B(_04327_),
    .X(_01137_));
 sg13g2_mux2_1 _10566_ (.A0(\shift_storage.storage [492]),
    .A1(\shift_storage.storage [491]),
    .S(_04322_),
    .X(_04328_));
 sg13g2_and2_1 _10567_ (.A(_04317_),
    .B(_04328_),
    .X(_01138_));
 sg13g2_buf_1 _10568_ (.A(net407),
    .X(_04329_));
 sg13g2_mux2_1 _10569_ (.A0(\shift_storage.storage [493]),
    .A1(\shift_storage.storage [492]),
    .S(net335),
    .X(_04330_));
 sg13g2_and2_1 _10570_ (.A(net334),
    .B(_04330_),
    .X(_01139_));
 sg13g2_mux2_1 _10571_ (.A0(\shift_storage.storage [494]),
    .A1(\shift_storage.storage [493]),
    .S(net335),
    .X(_04331_));
 sg13g2_and2_1 _10572_ (.A(net334),
    .B(_04331_),
    .X(_01140_));
 sg13g2_mux2_1 _10573_ (.A0(\shift_storage.storage [495]),
    .A1(\shift_storage.storage [494]),
    .S(net335),
    .X(_04332_));
 sg13g2_and2_1 _10574_ (.A(net334),
    .B(_04332_),
    .X(_01141_));
 sg13g2_mux2_1 _10575_ (.A0(\shift_storage.storage [496]),
    .A1(\shift_storage.storage [495]),
    .S(net335),
    .X(_04333_));
 sg13g2_and2_1 _10576_ (.A(net334),
    .B(_04333_),
    .X(_01142_));
 sg13g2_buf_1 _10577_ (.A(net408),
    .X(_04334_));
 sg13g2_mux2_1 _10578_ (.A0(\shift_storage.storage [497]),
    .A1(\shift_storage.storage [496]),
    .S(net333),
    .X(_04335_));
 sg13g2_and2_1 _10579_ (.A(net334),
    .B(_04335_),
    .X(_01143_));
 sg13g2_mux2_1 _10580_ (.A0(\shift_storage.storage [498]),
    .A1(\shift_storage.storage [497]),
    .S(net333),
    .X(_04336_));
 sg13g2_and2_1 _10581_ (.A(net334),
    .B(_04336_),
    .X(_01144_));
 sg13g2_mux2_1 _10582_ (.A0(\shift_storage.storage [499]),
    .A1(\shift_storage.storage [498]),
    .S(net333),
    .X(_04337_));
 sg13g2_and2_1 _10583_ (.A(net334),
    .B(_04337_),
    .X(_01145_));
 sg13g2_mux2_1 _10584_ (.A0(\shift_storage.storage [49]),
    .A1(\shift_storage.storage [48]),
    .S(net333),
    .X(_04338_));
 sg13g2_and2_1 _10585_ (.A(net334),
    .B(_04338_),
    .X(_01146_));
 sg13g2_mux2_1 _10586_ (.A0(\shift_storage.storage [4]),
    .A1(\shift_storage.storage [3]),
    .S(_04334_),
    .X(_04339_));
 sg13g2_and2_1 _10587_ (.A(_04329_),
    .B(_04339_),
    .X(_01147_));
 sg13g2_mux2_1 _10588_ (.A0(\shift_storage.storage [500]),
    .A1(\shift_storage.storage [499]),
    .S(_04334_),
    .X(_04340_));
 sg13g2_and2_1 _10589_ (.A(_04329_),
    .B(_04340_),
    .X(_01148_));
 sg13g2_buf_1 _10590_ (.A(net407),
    .X(_04341_));
 sg13g2_mux2_1 _10591_ (.A0(\shift_storage.storage [501]),
    .A1(\shift_storage.storage [500]),
    .S(net333),
    .X(_04342_));
 sg13g2_and2_1 _10592_ (.A(net332),
    .B(_04342_),
    .X(_01149_));
 sg13g2_mux2_1 _10593_ (.A0(\shift_storage.storage [502]),
    .A1(\shift_storage.storage [501]),
    .S(net333),
    .X(_04343_));
 sg13g2_and2_1 _10594_ (.A(net332),
    .B(_04343_),
    .X(_01150_));
 sg13g2_mux2_1 _10595_ (.A0(\shift_storage.storage [503]),
    .A1(\shift_storage.storage [502]),
    .S(net333),
    .X(_04344_));
 sg13g2_and2_1 _10596_ (.A(_04341_),
    .B(_04344_),
    .X(_01151_));
 sg13g2_mux2_1 _10597_ (.A0(\shift_storage.storage [504]),
    .A1(\shift_storage.storage [503]),
    .S(net333),
    .X(_04345_));
 sg13g2_and2_1 _10598_ (.A(_04341_),
    .B(_04345_),
    .X(_01152_));
 sg13g2_buf_1 _10599_ (.A(net408),
    .X(_04346_));
 sg13g2_mux2_1 _10600_ (.A0(\shift_storage.storage [505]),
    .A1(\shift_storage.storage [504]),
    .S(net331),
    .X(_04347_));
 sg13g2_and2_1 _10601_ (.A(net332),
    .B(_04347_),
    .X(_01153_));
 sg13g2_mux2_1 _10602_ (.A0(\shift_storage.storage [506]),
    .A1(\shift_storage.storage [505]),
    .S(net331),
    .X(_04348_));
 sg13g2_and2_1 _10603_ (.A(net332),
    .B(_04348_),
    .X(_01154_));
 sg13g2_mux2_1 _10604_ (.A0(\shift_storage.storage [507]),
    .A1(\shift_storage.storage [506]),
    .S(net331),
    .X(_04349_));
 sg13g2_and2_1 _10605_ (.A(net332),
    .B(_04349_),
    .X(_01155_));
 sg13g2_mux2_1 _10606_ (.A0(\shift_storage.storage [508]),
    .A1(\shift_storage.storage [507]),
    .S(net331),
    .X(_04350_));
 sg13g2_and2_1 _10607_ (.A(net332),
    .B(_04350_),
    .X(_01156_));
 sg13g2_mux2_1 _10608_ (.A0(\shift_storage.storage [509]),
    .A1(\shift_storage.storage [508]),
    .S(_04346_),
    .X(_04351_));
 sg13g2_and2_1 _10609_ (.A(net332),
    .B(_04351_),
    .X(_01157_));
 sg13g2_mux2_1 _10610_ (.A0(\shift_storage.storage [50]),
    .A1(\shift_storage.storage [49]),
    .S(_04346_),
    .X(_04352_));
 sg13g2_and2_1 _10611_ (.A(net332),
    .B(_04352_),
    .X(_01158_));
 sg13g2_buf_1 _10612_ (.A(net407),
    .X(_04353_));
 sg13g2_mux2_1 _10613_ (.A0(\shift_storage.storage [510]),
    .A1(\shift_storage.storage [509]),
    .S(net331),
    .X(_04354_));
 sg13g2_and2_1 _10614_ (.A(net330),
    .B(_04354_),
    .X(_01159_));
 sg13g2_mux2_1 _10615_ (.A0(\shift_storage.storage [511]),
    .A1(\shift_storage.storage [510]),
    .S(net331),
    .X(_04355_));
 sg13g2_and2_1 _10616_ (.A(net330),
    .B(_04355_),
    .X(_01160_));
 sg13g2_mux2_1 _10617_ (.A0(\shift_storage.storage [512]),
    .A1(\shift_storage.storage [511]),
    .S(net331),
    .X(_04356_));
 sg13g2_and2_1 _10618_ (.A(_04353_),
    .B(_04356_),
    .X(_01161_));
 sg13g2_mux2_1 _10619_ (.A0(\shift_storage.storage [513]),
    .A1(\shift_storage.storage [512]),
    .S(net331),
    .X(_04357_));
 sg13g2_and2_1 _10620_ (.A(_04353_),
    .B(_04357_),
    .X(_01162_));
 sg13g2_buf_1 _10621_ (.A(net408),
    .X(_04358_));
 sg13g2_mux2_1 _10622_ (.A0(\shift_storage.storage [514]),
    .A1(\shift_storage.storage [513]),
    .S(net329),
    .X(_04359_));
 sg13g2_and2_1 _10623_ (.A(net330),
    .B(_04359_),
    .X(_01163_));
 sg13g2_mux2_1 _10624_ (.A0(\shift_storage.storage [515]),
    .A1(\shift_storage.storage [514]),
    .S(net329),
    .X(_04360_));
 sg13g2_and2_1 _10625_ (.A(net330),
    .B(_04360_),
    .X(_01164_));
 sg13g2_mux2_1 _10626_ (.A0(\shift_storage.storage [516]),
    .A1(\shift_storage.storage [515]),
    .S(net329),
    .X(_04361_));
 sg13g2_and2_1 _10627_ (.A(net330),
    .B(_04361_),
    .X(_01165_));
 sg13g2_mux2_1 _10628_ (.A0(\shift_storage.storage [517]),
    .A1(\shift_storage.storage [516]),
    .S(net329),
    .X(_04362_));
 sg13g2_and2_1 _10629_ (.A(net330),
    .B(_04362_),
    .X(_01166_));
 sg13g2_mux2_1 _10630_ (.A0(\shift_storage.storage [518]),
    .A1(\shift_storage.storage [517]),
    .S(_04358_),
    .X(_04363_));
 sg13g2_and2_1 _10631_ (.A(net330),
    .B(_04363_),
    .X(_01167_));
 sg13g2_mux2_1 _10632_ (.A0(\shift_storage.storage [519]),
    .A1(\shift_storage.storage [518]),
    .S(net329),
    .X(_04364_));
 sg13g2_and2_1 _10633_ (.A(net330),
    .B(_04364_),
    .X(_01168_));
 sg13g2_buf_1 _10634_ (.A(net407),
    .X(_04365_));
 sg13g2_mux2_1 _10635_ (.A0(\shift_storage.storage [51]),
    .A1(\shift_storage.storage [50]),
    .S(_04358_),
    .X(_04366_));
 sg13g2_and2_1 _10636_ (.A(net328),
    .B(_04366_),
    .X(_01169_));
 sg13g2_mux2_1 _10637_ (.A0(\shift_storage.storage [520]),
    .A1(\shift_storage.storage [519]),
    .S(net329),
    .X(_04367_));
 sg13g2_and2_1 _10638_ (.A(net328),
    .B(_04367_),
    .X(_01170_));
 sg13g2_mux2_1 _10639_ (.A0(\shift_storage.storage [521]),
    .A1(\shift_storage.storage [520]),
    .S(net329),
    .X(_04368_));
 sg13g2_and2_1 _10640_ (.A(net328),
    .B(_04368_),
    .X(_01171_));
 sg13g2_mux2_1 _10641_ (.A0(\shift_storage.storage [522]),
    .A1(\shift_storage.storage [521]),
    .S(net329),
    .X(_04369_));
 sg13g2_and2_1 _10642_ (.A(net328),
    .B(_04369_),
    .X(_01172_));
 sg13g2_buf_1 _10643_ (.A(net408),
    .X(_04370_));
 sg13g2_mux2_1 _10644_ (.A0(\shift_storage.storage [523]),
    .A1(\shift_storage.storage [522]),
    .S(net327),
    .X(_04371_));
 sg13g2_and2_1 _10645_ (.A(net328),
    .B(_04371_),
    .X(_01173_));
 sg13g2_mux2_1 _10646_ (.A0(\shift_storage.storage [524]),
    .A1(\shift_storage.storage [523]),
    .S(net327),
    .X(_04372_));
 sg13g2_and2_1 _10647_ (.A(net328),
    .B(_04372_),
    .X(_01174_));
 sg13g2_mux2_1 _10648_ (.A0(\shift_storage.storage [525]),
    .A1(\shift_storage.storage [524]),
    .S(net327),
    .X(_04373_));
 sg13g2_and2_1 _10649_ (.A(net328),
    .B(_04373_),
    .X(_01175_));
 sg13g2_mux2_1 _10650_ (.A0(\shift_storage.storage [526]),
    .A1(\shift_storage.storage [525]),
    .S(net327),
    .X(_04374_));
 sg13g2_and2_1 _10651_ (.A(net328),
    .B(_04374_),
    .X(_01176_));
 sg13g2_mux2_1 _10652_ (.A0(\shift_storage.storage [527]),
    .A1(\shift_storage.storage [526]),
    .S(net327),
    .X(_04375_));
 sg13g2_and2_1 _10653_ (.A(_04365_),
    .B(_04375_),
    .X(_01177_));
 sg13g2_mux2_1 _10654_ (.A0(\shift_storage.storage [528]),
    .A1(\shift_storage.storage [527]),
    .S(net327),
    .X(_04376_));
 sg13g2_and2_1 _10655_ (.A(_04365_),
    .B(_04376_),
    .X(_01178_));
 sg13g2_buf_1 _10656_ (.A(net407),
    .X(_04377_));
 sg13g2_mux2_1 _10657_ (.A0(\shift_storage.storage [529]),
    .A1(\shift_storage.storage [528]),
    .S(net327),
    .X(_04378_));
 sg13g2_and2_1 _10658_ (.A(net326),
    .B(_04378_),
    .X(_01179_));
 sg13g2_mux2_1 _10659_ (.A0(\shift_storage.storage [52]),
    .A1(\shift_storage.storage [51]),
    .S(net327),
    .X(_04379_));
 sg13g2_and2_1 _10660_ (.A(net326),
    .B(_04379_),
    .X(_01180_));
 sg13g2_mux2_1 _10661_ (.A0(\shift_storage.storage [530]),
    .A1(\shift_storage.storage [529]),
    .S(_04370_),
    .X(_04380_));
 sg13g2_and2_1 _10662_ (.A(net326),
    .B(_04380_),
    .X(_01181_));
 sg13g2_mux2_1 _10663_ (.A0(\shift_storage.storage [531]),
    .A1(\shift_storage.storage [530]),
    .S(_04370_),
    .X(_04381_));
 sg13g2_and2_1 _10664_ (.A(net326),
    .B(_04381_),
    .X(_01182_));
 sg13g2_buf_1 _10665_ (.A(net408),
    .X(_04382_));
 sg13g2_mux2_1 _10666_ (.A0(\shift_storage.storage [532]),
    .A1(\shift_storage.storage [531]),
    .S(net325),
    .X(_04383_));
 sg13g2_and2_1 _10667_ (.A(net326),
    .B(_04383_),
    .X(_01183_));
 sg13g2_mux2_1 _10668_ (.A0(\shift_storage.storage [533]),
    .A1(\shift_storage.storage [532]),
    .S(net325),
    .X(_04384_));
 sg13g2_and2_1 _10669_ (.A(net326),
    .B(_04384_),
    .X(_01184_));
 sg13g2_mux2_1 _10670_ (.A0(\shift_storage.storage [534]),
    .A1(\shift_storage.storage [533]),
    .S(net325),
    .X(_04385_));
 sg13g2_and2_1 _10671_ (.A(net326),
    .B(_04385_),
    .X(_01185_));
 sg13g2_mux2_1 _10672_ (.A0(\shift_storage.storage [535]),
    .A1(\shift_storage.storage [534]),
    .S(net325),
    .X(_04386_));
 sg13g2_and2_1 _10673_ (.A(net326),
    .B(_04386_),
    .X(_01186_));
 sg13g2_mux2_1 _10674_ (.A0(\shift_storage.storage [536]),
    .A1(\shift_storage.storage [535]),
    .S(net325),
    .X(_04387_));
 sg13g2_and2_1 _10675_ (.A(_04377_),
    .B(_04387_),
    .X(_01187_));
 sg13g2_mux2_1 _10676_ (.A0(\shift_storage.storage [537]),
    .A1(\shift_storage.storage [536]),
    .S(net325),
    .X(_04388_));
 sg13g2_and2_1 _10677_ (.A(_04377_),
    .B(_04388_),
    .X(_01188_));
 sg13g2_buf_1 _10678_ (.A(net407),
    .X(_04389_));
 sg13g2_mux2_1 _10679_ (.A0(\shift_storage.storage [538]),
    .A1(\shift_storage.storage [537]),
    .S(net325),
    .X(_04390_));
 sg13g2_and2_1 _10680_ (.A(net324),
    .B(_04390_),
    .X(_01189_));
 sg13g2_mux2_1 _10681_ (.A0(\shift_storage.storage [539]),
    .A1(\shift_storage.storage [538]),
    .S(_04382_),
    .X(_04391_));
 sg13g2_and2_1 _10682_ (.A(net324),
    .B(_04391_),
    .X(_01190_));
 sg13g2_mux2_1 _10683_ (.A0(\shift_storage.storage [53]),
    .A1(\shift_storage.storage [52]),
    .S(net325),
    .X(_04392_));
 sg13g2_and2_1 _10684_ (.A(net324),
    .B(_04392_),
    .X(_01191_));
 sg13g2_mux2_1 _10685_ (.A0(\shift_storage.storage [540]),
    .A1(\shift_storage.storage [539]),
    .S(_04382_),
    .X(_04393_));
 sg13g2_and2_1 _10686_ (.A(net324),
    .B(_04393_),
    .X(_01192_));
 sg13g2_buf_1 _10687_ (.A(_03058_),
    .X(_04394_));
 sg13g2_buf_1 _10688_ (.A(net406),
    .X(_04395_));
 sg13g2_mux2_1 _10689_ (.A0(\shift_storage.storage [541]),
    .A1(\shift_storage.storage [540]),
    .S(net323),
    .X(_04396_));
 sg13g2_and2_1 _10690_ (.A(_04389_),
    .B(_04396_),
    .X(_01193_));
 sg13g2_mux2_1 _10691_ (.A0(\shift_storage.storage [542]),
    .A1(\shift_storage.storage [541]),
    .S(net323),
    .X(_04397_));
 sg13g2_and2_1 _10692_ (.A(_04389_),
    .B(_04397_),
    .X(_01194_));
 sg13g2_mux2_1 _10693_ (.A0(\shift_storage.storage [543]),
    .A1(\shift_storage.storage [542]),
    .S(_04395_),
    .X(_04398_));
 sg13g2_and2_1 _10694_ (.A(net324),
    .B(_04398_),
    .X(_01195_));
 sg13g2_mux2_1 _10695_ (.A0(\shift_storage.storage [544]),
    .A1(\shift_storage.storage [543]),
    .S(net323),
    .X(_04399_));
 sg13g2_and2_1 _10696_ (.A(net324),
    .B(_04399_),
    .X(_01196_));
 sg13g2_mux2_1 _10697_ (.A0(\shift_storage.storage [545]),
    .A1(\shift_storage.storage [544]),
    .S(net323),
    .X(_04400_));
 sg13g2_and2_1 _10698_ (.A(net324),
    .B(_04400_),
    .X(_01197_));
 sg13g2_mux2_1 _10699_ (.A0(\shift_storage.storage [546]),
    .A1(\shift_storage.storage [545]),
    .S(net323),
    .X(_04401_));
 sg13g2_and2_1 _10700_ (.A(net324),
    .B(_04401_),
    .X(_01198_));
 sg13g2_buf_1 _10701_ (.A(net494),
    .X(_04402_));
 sg13g2_buf_1 _10702_ (.A(net405),
    .X(_04403_));
 sg13g2_mux2_1 _10703_ (.A0(\shift_storage.storage [547]),
    .A1(\shift_storage.storage [546]),
    .S(net323),
    .X(_04404_));
 sg13g2_and2_1 _10704_ (.A(net322),
    .B(_04404_),
    .X(_01199_));
 sg13g2_mux2_1 _10705_ (.A0(\shift_storage.storage [548]),
    .A1(\shift_storage.storage [547]),
    .S(net323),
    .X(_04405_));
 sg13g2_and2_1 _10706_ (.A(net322),
    .B(_04405_),
    .X(_01200_));
 sg13g2_mux2_1 _10707_ (.A0(\shift_storage.storage [549]),
    .A1(\shift_storage.storage [548]),
    .S(net323),
    .X(_04406_));
 sg13g2_and2_1 _10708_ (.A(_04403_),
    .B(_04406_),
    .X(_01201_));
 sg13g2_mux2_1 _10709_ (.A0(\shift_storage.storage [54]),
    .A1(\shift_storage.storage [53]),
    .S(_04395_),
    .X(_04407_));
 sg13g2_and2_1 _10710_ (.A(_04403_),
    .B(_04407_),
    .X(_01202_));
 sg13g2_buf_1 _10711_ (.A(net406),
    .X(_04408_));
 sg13g2_mux2_1 _10712_ (.A0(\shift_storage.storage [550]),
    .A1(\shift_storage.storage [549]),
    .S(net321),
    .X(_04409_));
 sg13g2_and2_1 _10713_ (.A(net322),
    .B(_04409_),
    .X(_01203_));
 sg13g2_mux2_1 _10714_ (.A0(\shift_storage.storage [551]),
    .A1(\shift_storage.storage [550]),
    .S(net321),
    .X(_04410_));
 sg13g2_and2_1 _10715_ (.A(net322),
    .B(_04410_),
    .X(_01204_));
 sg13g2_mux2_1 _10716_ (.A0(\shift_storage.storage [552]),
    .A1(\shift_storage.storage [551]),
    .S(net321),
    .X(_04411_));
 sg13g2_and2_1 _10717_ (.A(net322),
    .B(_04411_),
    .X(_01205_));
 sg13g2_mux2_1 _10718_ (.A0(\shift_storage.storage [553]),
    .A1(\shift_storage.storage [552]),
    .S(net321),
    .X(_04412_));
 sg13g2_and2_1 _10719_ (.A(net322),
    .B(_04412_),
    .X(_01206_));
 sg13g2_mux2_1 _10720_ (.A0(\shift_storage.storage [554]),
    .A1(\shift_storage.storage [553]),
    .S(_04408_),
    .X(_04413_));
 sg13g2_and2_1 _10721_ (.A(net322),
    .B(_04413_),
    .X(_01207_));
 sg13g2_mux2_1 _10722_ (.A0(\shift_storage.storage [555]),
    .A1(\shift_storage.storage [554]),
    .S(_04408_),
    .X(_04414_));
 sg13g2_and2_1 _10723_ (.A(net322),
    .B(_04414_),
    .X(_01208_));
 sg13g2_buf_1 _10724_ (.A(net405),
    .X(_04415_));
 sg13g2_mux2_1 _10725_ (.A0(\shift_storage.storage [556]),
    .A1(\shift_storage.storage [555]),
    .S(net321),
    .X(_04416_));
 sg13g2_and2_1 _10726_ (.A(net320),
    .B(_04416_),
    .X(_01209_));
 sg13g2_mux2_1 _10727_ (.A0(\shift_storage.storage [557]),
    .A1(\shift_storage.storage [556]),
    .S(net321),
    .X(_04417_));
 sg13g2_and2_1 _10728_ (.A(net320),
    .B(_04417_),
    .X(_01210_));
 sg13g2_mux2_1 _10729_ (.A0(\shift_storage.storage [558]),
    .A1(\shift_storage.storage [557]),
    .S(net321),
    .X(_04418_));
 sg13g2_and2_1 _10730_ (.A(net320),
    .B(_04418_),
    .X(_01211_));
 sg13g2_mux2_1 _10731_ (.A0(\shift_storage.storage [559]),
    .A1(\shift_storage.storage [558]),
    .S(net321),
    .X(_04419_));
 sg13g2_and2_1 _10732_ (.A(net320),
    .B(_04419_),
    .X(_01212_));
 sg13g2_buf_1 _10733_ (.A(net406),
    .X(_04420_));
 sg13g2_mux2_1 _10734_ (.A0(\shift_storage.storage [55]),
    .A1(\shift_storage.storage [54]),
    .S(net319),
    .X(_04421_));
 sg13g2_and2_1 _10735_ (.A(net320),
    .B(_04421_),
    .X(_01213_));
 sg13g2_mux2_1 _10736_ (.A0(\shift_storage.storage [560]),
    .A1(\shift_storage.storage [559]),
    .S(net319),
    .X(_04422_));
 sg13g2_and2_1 _10737_ (.A(net320),
    .B(_04422_),
    .X(_01214_));
 sg13g2_mux2_1 _10738_ (.A0(\shift_storage.storage [561]),
    .A1(\shift_storage.storage [560]),
    .S(net319),
    .X(_04423_));
 sg13g2_and2_1 _10739_ (.A(net320),
    .B(_04423_),
    .X(_01215_));
 sg13g2_mux2_1 _10740_ (.A0(\shift_storage.storage [562]),
    .A1(\shift_storage.storage [561]),
    .S(net319),
    .X(_04424_));
 sg13g2_and2_1 _10741_ (.A(net320),
    .B(_04424_),
    .X(_01216_));
 sg13g2_mux2_1 _10742_ (.A0(\shift_storage.storage [563]),
    .A1(\shift_storage.storage [562]),
    .S(_04420_),
    .X(_04425_));
 sg13g2_and2_1 _10743_ (.A(_04415_),
    .B(_04425_),
    .X(_01217_));
 sg13g2_mux2_1 _10744_ (.A0(\shift_storage.storage [564]),
    .A1(\shift_storage.storage [563]),
    .S(_04420_),
    .X(_04426_));
 sg13g2_and2_1 _10745_ (.A(_04415_),
    .B(_04426_),
    .X(_01218_));
 sg13g2_buf_1 _10746_ (.A(_04402_),
    .X(_04427_));
 sg13g2_mux2_1 _10747_ (.A0(\shift_storage.storage [565]),
    .A1(\shift_storage.storage [564]),
    .S(net319),
    .X(_04428_));
 sg13g2_and2_1 _10748_ (.A(net318),
    .B(_04428_),
    .X(_01219_));
 sg13g2_mux2_1 _10749_ (.A0(\shift_storage.storage [566]),
    .A1(\shift_storage.storage [565]),
    .S(net319),
    .X(_04429_));
 sg13g2_and2_1 _10750_ (.A(net318),
    .B(_04429_),
    .X(_01220_));
 sg13g2_mux2_1 _10751_ (.A0(\shift_storage.storage [567]),
    .A1(\shift_storage.storage [566]),
    .S(net319),
    .X(_04430_));
 sg13g2_and2_1 _10752_ (.A(_04427_),
    .B(_04430_),
    .X(_01221_));
 sg13g2_mux2_1 _10753_ (.A0(\shift_storage.storage [568]),
    .A1(\shift_storage.storage [567]),
    .S(net319),
    .X(_04431_));
 sg13g2_and2_1 _10754_ (.A(_04427_),
    .B(_04431_),
    .X(_01222_));
 sg13g2_buf_1 _10755_ (.A(net406),
    .X(_04432_));
 sg13g2_mux2_1 _10756_ (.A0(\shift_storage.storage [569]),
    .A1(\shift_storage.storage [568]),
    .S(net317),
    .X(_04433_));
 sg13g2_and2_1 _10757_ (.A(net318),
    .B(_04433_),
    .X(_01223_));
 sg13g2_mux2_1 _10758_ (.A0(\shift_storage.storage [56]),
    .A1(\shift_storage.storage [55]),
    .S(net317),
    .X(_04434_));
 sg13g2_and2_1 _10759_ (.A(net318),
    .B(_04434_),
    .X(_01224_));
 sg13g2_mux2_1 _10760_ (.A0(\shift_storage.storage [570]),
    .A1(\shift_storage.storage [569]),
    .S(net317),
    .X(_04435_));
 sg13g2_and2_1 _10761_ (.A(net318),
    .B(_04435_),
    .X(_01225_));
 sg13g2_mux2_1 _10762_ (.A0(\shift_storage.storage [571]),
    .A1(\shift_storage.storage [570]),
    .S(net317),
    .X(_04436_));
 sg13g2_and2_1 _10763_ (.A(net318),
    .B(_04436_),
    .X(_01226_));
 sg13g2_mux2_1 _10764_ (.A0(\shift_storage.storage [572]),
    .A1(\shift_storage.storage [571]),
    .S(net317),
    .X(_04437_));
 sg13g2_and2_1 _10765_ (.A(net318),
    .B(_04437_),
    .X(_01227_));
 sg13g2_mux2_1 _10766_ (.A0(\shift_storage.storage [573]),
    .A1(\shift_storage.storage [572]),
    .S(net317),
    .X(_04438_));
 sg13g2_and2_1 _10767_ (.A(net318),
    .B(_04438_),
    .X(_01228_));
 sg13g2_buf_1 _10768_ (.A(net405),
    .X(_04439_));
 sg13g2_mux2_1 _10769_ (.A0(\shift_storage.storage [574]),
    .A1(\shift_storage.storage [573]),
    .S(net317),
    .X(_04440_));
 sg13g2_and2_1 _10770_ (.A(net316),
    .B(_04440_),
    .X(_01229_));
 sg13g2_mux2_1 _10771_ (.A0(\shift_storage.storage [575]),
    .A1(\shift_storage.storage [574]),
    .S(net317),
    .X(_04441_));
 sg13g2_and2_1 _10772_ (.A(net316),
    .B(_04441_),
    .X(_01230_));
 sg13g2_mux2_1 _10773_ (.A0(\shift_storage.storage [576]),
    .A1(\shift_storage.storage [575]),
    .S(_04432_),
    .X(_04442_));
 sg13g2_and2_1 _10774_ (.A(net316),
    .B(_04442_),
    .X(_01231_));
 sg13g2_mux2_1 _10775_ (.A0(\shift_storage.storage [577]),
    .A1(\shift_storage.storage [576]),
    .S(_04432_),
    .X(_04443_));
 sg13g2_and2_1 _10776_ (.A(net316),
    .B(_04443_),
    .X(_01232_));
 sg13g2_buf_1 _10777_ (.A(_04394_),
    .X(_04444_));
 sg13g2_mux2_1 _10778_ (.A0(\shift_storage.storage [578]),
    .A1(\shift_storage.storage [577]),
    .S(net315),
    .X(_04445_));
 sg13g2_and2_1 _10779_ (.A(net316),
    .B(_04445_),
    .X(_01233_));
 sg13g2_mux2_1 _10780_ (.A0(\shift_storage.storage [579]),
    .A1(\shift_storage.storage [578]),
    .S(net315),
    .X(_04446_));
 sg13g2_and2_1 _10781_ (.A(net316),
    .B(_04446_),
    .X(_01234_));
 sg13g2_mux2_1 _10782_ (.A0(\shift_storage.storage [57]),
    .A1(\shift_storage.storage [56]),
    .S(net315),
    .X(_04447_));
 sg13g2_and2_1 _10783_ (.A(net316),
    .B(_04447_),
    .X(_01235_));
 sg13g2_mux2_1 _10784_ (.A0(\shift_storage.storage [580]),
    .A1(\shift_storage.storage [579]),
    .S(net315),
    .X(_04448_));
 sg13g2_and2_1 _10785_ (.A(net316),
    .B(_04448_),
    .X(_01236_));
 sg13g2_mux2_1 _10786_ (.A0(\shift_storage.storage [581]),
    .A1(\shift_storage.storage [580]),
    .S(net315),
    .X(_04449_));
 sg13g2_and2_1 _10787_ (.A(_04439_),
    .B(_04449_),
    .X(_01237_));
 sg13g2_mux2_1 _10788_ (.A0(\shift_storage.storage [582]),
    .A1(\shift_storage.storage [581]),
    .S(net315),
    .X(_04450_));
 sg13g2_and2_1 _10789_ (.A(_04439_),
    .B(_04450_),
    .X(_01238_));
 sg13g2_buf_1 _10790_ (.A(_04402_),
    .X(_04451_));
 sg13g2_mux2_1 _10791_ (.A0(\shift_storage.storage [583]),
    .A1(\shift_storage.storage [582]),
    .S(net315),
    .X(_04452_));
 sg13g2_and2_1 _10792_ (.A(net314),
    .B(_04452_),
    .X(_01239_));
 sg13g2_mux2_1 _10793_ (.A0(\shift_storage.storage [584]),
    .A1(\shift_storage.storage [583]),
    .S(net315),
    .X(_04453_));
 sg13g2_and2_1 _10794_ (.A(net314),
    .B(_04453_),
    .X(_01240_));
 sg13g2_mux2_1 _10795_ (.A0(\shift_storage.storage [585]),
    .A1(\shift_storage.storage [584]),
    .S(_04444_),
    .X(_04454_));
 sg13g2_and2_1 _10796_ (.A(net314),
    .B(_04454_),
    .X(_01241_));
 sg13g2_mux2_1 _10797_ (.A0(\shift_storage.storage [586]),
    .A1(\shift_storage.storage [585]),
    .S(_04444_),
    .X(_04455_));
 sg13g2_and2_1 _10798_ (.A(net314),
    .B(_04455_),
    .X(_01242_));
 sg13g2_buf_1 _10799_ (.A(_04394_),
    .X(_04456_));
 sg13g2_mux2_1 _10800_ (.A0(\shift_storage.storage [587]),
    .A1(\shift_storage.storage [586]),
    .S(net313),
    .X(_04457_));
 sg13g2_and2_1 _10801_ (.A(net314),
    .B(_04457_),
    .X(_01243_));
 sg13g2_mux2_1 _10802_ (.A0(\shift_storage.storage [588]),
    .A1(\shift_storage.storage [587]),
    .S(net313),
    .X(_04458_));
 sg13g2_and2_1 _10803_ (.A(net314),
    .B(_04458_),
    .X(_01244_));
 sg13g2_mux2_1 _10804_ (.A0(\shift_storage.storage [589]),
    .A1(\shift_storage.storage [588]),
    .S(net313),
    .X(_04459_));
 sg13g2_and2_1 _10805_ (.A(net314),
    .B(_04459_),
    .X(_01245_));
 sg13g2_mux2_1 _10806_ (.A0(\shift_storage.storage [58]),
    .A1(\shift_storage.storage [57]),
    .S(net313),
    .X(_04460_));
 sg13g2_and2_1 _10807_ (.A(net314),
    .B(_04460_),
    .X(_01246_));
 sg13g2_mux2_1 _10808_ (.A0(\shift_storage.storage [590]),
    .A1(\shift_storage.storage [589]),
    .S(net313),
    .X(_04461_));
 sg13g2_and2_1 _10809_ (.A(_04451_),
    .B(_04461_),
    .X(_01247_));
 sg13g2_mux2_1 _10810_ (.A0(\shift_storage.storage [591]),
    .A1(\shift_storage.storage [590]),
    .S(net313),
    .X(_04462_));
 sg13g2_and2_1 _10811_ (.A(_04451_),
    .B(_04462_),
    .X(_01248_));
 sg13g2_buf_1 _10812_ (.A(net405),
    .X(_04463_));
 sg13g2_mux2_1 _10813_ (.A0(\shift_storage.storage [592]),
    .A1(\shift_storage.storage [591]),
    .S(_04456_),
    .X(_04464_));
 sg13g2_and2_1 _10814_ (.A(net312),
    .B(_04464_),
    .X(_01249_));
 sg13g2_mux2_1 _10815_ (.A0(\shift_storage.storage [593]),
    .A1(\shift_storage.storage [592]),
    .S(_04456_),
    .X(_04465_));
 sg13g2_and2_1 _10816_ (.A(net312),
    .B(_04465_),
    .X(_01250_));
 sg13g2_mux2_1 _10817_ (.A0(\shift_storage.storage [594]),
    .A1(\shift_storage.storage [593]),
    .S(net313),
    .X(_04466_));
 sg13g2_and2_1 _10818_ (.A(net312),
    .B(_04466_),
    .X(_01251_));
 sg13g2_mux2_1 _10819_ (.A0(\shift_storage.storage [595]),
    .A1(\shift_storage.storage [594]),
    .S(net313),
    .X(_04467_));
 sg13g2_and2_1 _10820_ (.A(net312),
    .B(_04467_),
    .X(_01252_));
 sg13g2_buf_1 _10821_ (.A(net406),
    .X(_04468_));
 sg13g2_mux2_1 _10822_ (.A0(\shift_storage.storage [596]),
    .A1(\shift_storage.storage [595]),
    .S(net311),
    .X(_04469_));
 sg13g2_and2_1 _10823_ (.A(net312),
    .B(_04469_),
    .X(_01253_));
 sg13g2_mux2_1 _10824_ (.A0(\shift_storage.storage [597]),
    .A1(\shift_storage.storage [596]),
    .S(net311),
    .X(_04470_));
 sg13g2_and2_1 _10825_ (.A(net312),
    .B(_04470_),
    .X(_01254_));
 sg13g2_mux2_1 _10826_ (.A0(\shift_storage.storage [598]),
    .A1(\shift_storage.storage [597]),
    .S(net311),
    .X(_04471_));
 sg13g2_and2_1 _10827_ (.A(net312),
    .B(_04471_),
    .X(_01255_));
 sg13g2_mux2_1 _10828_ (.A0(\shift_storage.storage [599]),
    .A1(\shift_storage.storage [598]),
    .S(net311),
    .X(_04472_));
 sg13g2_and2_1 _10829_ (.A(_04463_),
    .B(_04472_),
    .X(_01256_));
 sg13g2_mux2_1 _10830_ (.A0(\shift_storage.storage [59]),
    .A1(\shift_storage.storage [58]),
    .S(net311),
    .X(_04473_));
 sg13g2_and2_1 _10831_ (.A(net312),
    .B(_04473_),
    .X(_01257_));
 sg13g2_mux2_1 _10832_ (.A0(\shift_storage.storage [5]),
    .A1(\shift_storage.storage [4]),
    .S(net311),
    .X(_04474_));
 sg13g2_and2_1 _10833_ (.A(_04463_),
    .B(_04474_),
    .X(_01258_));
 sg13g2_buf_1 _10834_ (.A(net405),
    .X(_04475_));
 sg13g2_mux2_1 _10835_ (.A0(\shift_storage.storage [600]),
    .A1(\shift_storage.storage [599]),
    .S(net311),
    .X(_04476_));
 sg13g2_and2_1 _10836_ (.A(net310),
    .B(_04476_),
    .X(_01259_));
 sg13g2_mux2_1 _10837_ (.A0(\shift_storage.storage [601]),
    .A1(\shift_storage.storage [600]),
    .S(net311),
    .X(_04477_));
 sg13g2_and2_1 _10838_ (.A(net310),
    .B(_04477_),
    .X(_01260_));
 sg13g2_mux2_1 _10839_ (.A0(\shift_storage.storage [602]),
    .A1(\shift_storage.storage [601]),
    .S(_04468_),
    .X(_04478_));
 sg13g2_and2_1 _10840_ (.A(_04475_),
    .B(_04478_),
    .X(_01261_));
 sg13g2_mux2_1 _10841_ (.A0(\shift_storage.storage [603]),
    .A1(\shift_storage.storage [602]),
    .S(_04468_),
    .X(_04479_));
 sg13g2_and2_1 _10842_ (.A(_04475_),
    .B(_04479_),
    .X(_01262_));
 sg13g2_buf_1 _10843_ (.A(net406),
    .X(_04480_));
 sg13g2_mux2_1 _10844_ (.A0(\shift_storage.storage [604]),
    .A1(\shift_storage.storage [603]),
    .S(net309),
    .X(_04481_));
 sg13g2_and2_1 _10845_ (.A(net310),
    .B(_04481_),
    .X(_01263_));
 sg13g2_mux2_1 _10846_ (.A0(\shift_storage.storage [605]),
    .A1(\shift_storage.storage [604]),
    .S(net309),
    .X(_04482_));
 sg13g2_and2_1 _10847_ (.A(net310),
    .B(_04482_),
    .X(_01264_));
 sg13g2_mux2_1 _10848_ (.A0(\shift_storage.storage [606]),
    .A1(\shift_storage.storage [605]),
    .S(net309),
    .X(_04483_));
 sg13g2_and2_1 _10849_ (.A(net310),
    .B(_04483_),
    .X(_01265_));
 sg13g2_mux2_1 _10850_ (.A0(\shift_storage.storage [607]),
    .A1(\shift_storage.storage [606]),
    .S(net309),
    .X(_04484_));
 sg13g2_and2_1 _10851_ (.A(net310),
    .B(_04484_),
    .X(_01266_));
 sg13g2_mux2_1 _10852_ (.A0(\shift_storage.storage [608]),
    .A1(\shift_storage.storage [607]),
    .S(net309),
    .X(_04485_));
 sg13g2_and2_1 _10853_ (.A(net310),
    .B(_04485_),
    .X(_01267_));
 sg13g2_mux2_1 _10854_ (.A0(\shift_storage.storage [609]),
    .A1(\shift_storage.storage [608]),
    .S(_04480_),
    .X(_04486_));
 sg13g2_and2_1 _10855_ (.A(net310),
    .B(_04486_),
    .X(_01268_));
 sg13g2_buf_1 _10856_ (.A(net405),
    .X(_04487_));
 sg13g2_mux2_1 _10857_ (.A0(\shift_storage.storage [60]),
    .A1(\shift_storage.storage [59]),
    .S(_04480_),
    .X(_04488_));
 sg13g2_and2_1 _10858_ (.A(net308),
    .B(_04488_),
    .X(_01269_));
 sg13g2_mux2_1 _10859_ (.A0(\shift_storage.storage [610]),
    .A1(\shift_storage.storage [609]),
    .S(net309),
    .X(_04489_));
 sg13g2_and2_1 _10860_ (.A(net308),
    .B(_04489_),
    .X(_01270_));
 sg13g2_mux2_1 _10861_ (.A0(\shift_storage.storage [611]),
    .A1(\shift_storage.storage [610]),
    .S(net309),
    .X(_04490_));
 sg13g2_and2_1 _10862_ (.A(net308),
    .B(_04490_),
    .X(_01271_));
 sg13g2_mux2_1 _10863_ (.A0(\shift_storage.storage [612]),
    .A1(\shift_storage.storage [611]),
    .S(net309),
    .X(_04491_));
 sg13g2_and2_1 _10864_ (.A(net308),
    .B(_04491_),
    .X(_01272_));
 sg13g2_buf_1 _10865_ (.A(net406),
    .X(_04492_));
 sg13g2_mux2_1 _10866_ (.A0(\shift_storage.storage [613]),
    .A1(\shift_storage.storage [612]),
    .S(net307),
    .X(_04493_));
 sg13g2_and2_1 _10867_ (.A(net308),
    .B(_04493_),
    .X(_01273_));
 sg13g2_mux2_1 _10868_ (.A0(\shift_storage.storage [614]),
    .A1(\shift_storage.storage [613]),
    .S(net307),
    .X(_04494_));
 sg13g2_and2_1 _10869_ (.A(net308),
    .B(_04494_),
    .X(_01274_));
 sg13g2_mux2_1 _10870_ (.A0(\shift_storage.storage [615]),
    .A1(\shift_storage.storage [614]),
    .S(net307),
    .X(_04495_));
 sg13g2_and2_1 _10871_ (.A(net308),
    .B(_04495_),
    .X(_01275_));
 sg13g2_mux2_1 _10872_ (.A0(\shift_storage.storage [616]),
    .A1(\shift_storage.storage [615]),
    .S(net307),
    .X(_04496_));
 sg13g2_and2_1 _10873_ (.A(net308),
    .B(_04496_),
    .X(_01276_));
 sg13g2_mux2_1 _10874_ (.A0(\shift_storage.storage [617]),
    .A1(\shift_storage.storage [616]),
    .S(net307),
    .X(_04497_));
 sg13g2_and2_1 _10875_ (.A(_04487_),
    .B(_04497_),
    .X(_01277_));
 sg13g2_mux2_1 _10876_ (.A0(\shift_storage.storage [618]),
    .A1(\shift_storage.storage [617]),
    .S(net307),
    .X(_04498_));
 sg13g2_and2_1 _10877_ (.A(_04487_),
    .B(_04498_),
    .X(_01278_));
 sg13g2_buf_1 _10878_ (.A(net405),
    .X(_04499_));
 sg13g2_mux2_1 _10879_ (.A0(\shift_storage.storage [619]),
    .A1(\shift_storage.storage [618]),
    .S(net307),
    .X(_04500_));
 sg13g2_and2_1 _10880_ (.A(net306),
    .B(_04500_),
    .X(_01279_));
 sg13g2_mux2_1 _10881_ (.A0(\shift_storage.storage [61]),
    .A1(\shift_storage.storage [60]),
    .S(net307),
    .X(_04501_));
 sg13g2_and2_1 _10882_ (.A(net306),
    .B(_04501_),
    .X(_01280_));
 sg13g2_mux2_1 _10883_ (.A0(\shift_storage.storage [620]),
    .A1(\shift_storage.storage [619]),
    .S(_04492_),
    .X(_04502_));
 sg13g2_and2_1 _10884_ (.A(net306),
    .B(_04502_),
    .X(_01281_));
 sg13g2_mux2_1 _10885_ (.A0(\shift_storage.storage [621]),
    .A1(\shift_storage.storage [620]),
    .S(_04492_),
    .X(_04503_));
 sg13g2_and2_1 _10886_ (.A(_04499_),
    .B(_04503_),
    .X(_01282_));
 sg13g2_buf_1 _10887_ (.A(net406),
    .X(_04504_));
 sg13g2_mux2_1 _10888_ (.A0(\shift_storage.storage [622]),
    .A1(\shift_storage.storage [621]),
    .S(net305),
    .X(_04505_));
 sg13g2_and2_1 _10889_ (.A(_04499_),
    .B(_04505_),
    .X(_01283_));
 sg13g2_mux2_1 _10890_ (.A0(\shift_storage.storage [623]),
    .A1(\shift_storage.storage [622]),
    .S(_04504_),
    .X(_04506_));
 sg13g2_and2_1 _10891_ (.A(net306),
    .B(_04506_),
    .X(_01284_));
 sg13g2_mux2_1 _10892_ (.A0(\shift_storage.storage [624]),
    .A1(\shift_storage.storage [623]),
    .S(net305),
    .X(_04507_));
 sg13g2_and2_1 _10893_ (.A(net306),
    .B(_04507_),
    .X(_01285_));
 sg13g2_mux2_1 _10894_ (.A0(\shift_storage.storage [625]),
    .A1(\shift_storage.storage [624]),
    .S(net305),
    .X(_04508_));
 sg13g2_and2_1 _10895_ (.A(net306),
    .B(_04508_),
    .X(_01286_));
 sg13g2_mux2_1 _10896_ (.A0(\shift_storage.storage [626]),
    .A1(\shift_storage.storage [625]),
    .S(net305),
    .X(_04509_));
 sg13g2_and2_1 _10897_ (.A(net306),
    .B(_04509_),
    .X(_01287_));
 sg13g2_mux2_1 _10898_ (.A0(\shift_storage.storage [627]),
    .A1(\shift_storage.storage [626]),
    .S(net305),
    .X(_04510_));
 sg13g2_and2_1 _10899_ (.A(net306),
    .B(_04510_),
    .X(_01288_));
 sg13g2_buf_1 _10900_ (.A(net405),
    .X(_04511_));
 sg13g2_mux2_1 _10901_ (.A0(\shift_storage.storage [628]),
    .A1(\shift_storage.storage [627]),
    .S(net305),
    .X(_04512_));
 sg13g2_and2_1 _10902_ (.A(net304),
    .B(_04512_),
    .X(_01289_));
 sg13g2_mux2_1 _10903_ (.A0(\shift_storage.storage [629]),
    .A1(\shift_storage.storage [628]),
    .S(net305),
    .X(_04513_));
 sg13g2_and2_1 _10904_ (.A(net304),
    .B(_04513_),
    .X(_01290_));
 sg13g2_mux2_1 _10905_ (.A0(\shift_storage.storage [62]),
    .A1(\shift_storage.storage [61]),
    .S(_04504_),
    .X(_04514_));
 sg13g2_and2_1 _10906_ (.A(net304),
    .B(_04514_),
    .X(_01291_));
 sg13g2_mux2_1 _10907_ (.A0(\shift_storage.storage [630]),
    .A1(\shift_storage.storage [629]),
    .S(net305),
    .X(_04515_));
 sg13g2_and2_1 _10908_ (.A(net304),
    .B(_04515_),
    .X(_01292_));
 sg13g2_buf_1 _10909_ (.A(_03058_),
    .X(_04516_));
 sg13g2_buf_1 _10910_ (.A(net404),
    .X(_04517_));
 sg13g2_mux2_1 _10911_ (.A0(\shift_storage.storage [631]),
    .A1(\shift_storage.storage [630]),
    .S(net303),
    .X(_04518_));
 sg13g2_and2_1 _10912_ (.A(net304),
    .B(_04518_),
    .X(_01293_));
 sg13g2_mux2_1 _10913_ (.A0(\shift_storage.storage [632]),
    .A1(\shift_storage.storage [631]),
    .S(net303),
    .X(_04519_));
 sg13g2_and2_1 _10914_ (.A(net304),
    .B(_04519_),
    .X(_01294_));
 sg13g2_mux2_1 _10915_ (.A0(\shift_storage.storage [633]),
    .A1(\shift_storage.storage [632]),
    .S(net303),
    .X(_04520_));
 sg13g2_and2_1 _10916_ (.A(net304),
    .B(_04520_),
    .X(_01295_));
 sg13g2_mux2_1 _10917_ (.A0(\shift_storage.storage [634]),
    .A1(\shift_storage.storage [633]),
    .S(net303),
    .X(_04521_));
 sg13g2_and2_1 _10918_ (.A(net304),
    .B(_04521_),
    .X(_01296_));
 sg13g2_mux2_1 _10919_ (.A0(\shift_storage.storage [635]),
    .A1(\shift_storage.storage [634]),
    .S(net303),
    .X(_04522_));
 sg13g2_and2_1 _10920_ (.A(_04511_),
    .B(_04522_),
    .X(_01297_));
 sg13g2_mux2_1 _10921_ (.A0(\shift_storage.storage [636]),
    .A1(\shift_storage.storage [635]),
    .S(net303),
    .X(_04523_));
 sg13g2_and2_1 _10922_ (.A(_04511_),
    .B(_04523_),
    .X(_01298_));
 sg13g2_buf_1 _10923_ (.A(net494),
    .X(_04524_));
 sg13g2_buf_1 _10924_ (.A(net403),
    .X(_04525_));
 sg13g2_mux2_1 _10925_ (.A0(\shift_storage.storage [637]),
    .A1(\shift_storage.storage [636]),
    .S(_04517_),
    .X(_04526_));
 sg13g2_and2_1 _10926_ (.A(net302),
    .B(_04526_),
    .X(_01299_));
 sg13g2_mux2_1 _10927_ (.A0(\shift_storage.storage [638]),
    .A1(\shift_storage.storage [637]),
    .S(net303),
    .X(_04527_));
 sg13g2_and2_1 _10928_ (.A(net302),
    .B(_04527_),
    .X(_01300_));
 sg13g2_mux2_1 _10929_ (.A0(\shift_storage.storage [639]),
    .A1(\shift_storage.storage [638]),
    .S(net303),
    .X(_04528_));
 sg13g2_and2_1 _10930_ (.A(net302),
    .B(_04528_),
    .X(_01301_));
 sg13g2_mux2_1 _10931_ (.A0(\shift_storage.storage [63]),
    .A1(\shift_storage.storage [62]),
    .S(_04517_),
    .X(_04529_));
 sg13g2_and2_1 _10932_ (.A(net302),
    .B(_04529_),
    .X(_01302_));
 sg13g2_buf_1 _10933_ (.A(net404),
    .X(_04530_));
 sg13g2_mux2_1 _10934_ (.A0(\shift_storage.storage [640]),
    .A1(\shift_storage.storage [639]),
    .S(net301),
    .X(_04531_));
 sg13g2_and2_1 _10935_ (.A(net302),
    .B(_04531_),
    .X(_01303_));
 sg13g2_mux2_1 _10936_ (.A0(\shift_storage.storage [641]),
    .A1(\shift_storage.storage [640]),
    .S(net301),
    .X(_04532_));
 sg13g2_and2_1 _10937_ (.A(net302),
    .B(_04532_),
    .X(_01304_));
 sg13g2_mux2_1 _10938_ (.A0(\shift_storage.storage [642]),
    .A1(\shift_storage.storage [641]),
    .S(net301),
    .X(_04533_));
 sg13g2_and2_1 _10939_ (.A(net302),
    .B(_04533_),
    .X(_01305_));
 sg13g2_mux2_1 _10940_ (.A0(\shift_storage.storage [643]),
    .A1(\shift_storage.storage [642]),
    .S(net301),
    .X(_04534_));
 sg13g2_and2_1 _10941_ (.A(net302),
    .B(_04534_),
    .X(_01306_));
 sg13g2_mux2_1 _10942_ (.A0(\shift_storage.storage [644]),
    .A1(\shift_storage.storage [643]),
    .S(net301),
    .X(_04535_));
 sg13g2_and2_1 _10943_ (.A(_04525_),
    .B(_04535_),
    .X(_01307_));
 sg13g2_mux2_1 _10944_ (.A0(\shift_storage.storage [645]),
    .A1(\shift_storage.storage [644]),
    .S(net301),
    .X(_04536_));
 sg13g2_and2_1 _10945_ (.A(_04525_),
    .B(_04536_),
    .X(_01308_));
 sg13g2_buf_1 _10946_ (.A(net403),
    .X(_04537_));
 sg13g2_mux2_1 _10947_ (.A0(\shift_storage.storage [646]),
    .A1(\shift_storage.storage [645]),
    .S(_04530_),
    .X(_04538_));
 sg13g2_and2_1 _10948_ (.A(net300),
    .B(_04538_),
    .X(_01309_));
 sg13g2_mux2_1 _10949_ (.A0(\shift_storage.storage [647]),
    .A1(\shift_storage.storage [646]),
    .S(_04530_),
    .X(_04539_));
 sg13g2_and2_1 _10950_ (.A(net300),
    .B(_04539_),
    .X(_01310_));
 sg13g2_mux2_1 _10951_ (.A0(\shift_storage.storage [648]),
    .A1(\shift_storage.storage [647]),
    .S(net301),
    .X(_04540_));
 sg13g2_and2_1 _10952_ (.A(net300),
    .B(_04540_),
    .X(_01311_));
 sg13g2_mux2_1 _10953_ (.A0(\shift_storage.storage [649]),
    .A1(\shift_storage.storage [648]),
    .S(net301),
    .X(_04541_));
 sg13g2_and2_1 _10954_ (.A(net300),
    .B(_04541_),
    .X(_01312_));
 sg13g2_buf_1 _10955_ (.A(net404),
    .X(_04542_));
 sg13g2_mux2_1 _10956_ (.A0(\shift_storage.storage [64]),
    .A1(\shift_storage.storage [63]),
    .S(net299),
    .X(_04543_));
 sg13g2_and2_1 _10957_ (.A(_04537_),
    .B(_04543_),
    .X(_01313_));
 sg13g2_mux2_1 _10958_ (.A0(\shift_storage.storage [650]),
    .A1(\shift_storage.storage [649]),
    .S(net299),
    .X(_04544_));
 sg13g2_and2_1 _10959_ (.A(net300),
    .B(_04544_),
    .X(_01314_));
 sg13g2_mux2_1 _10960_ (.A0(\shift_storage.storage [651]),
    .A1(\shift_storage.storage [650]),
    .S(net299),
    .X(_04545_));
 sg13g2_and2_1 _10961_ (.A(net300),
    .B(_04545_),
    .X(_01315_));
 sg13g2_mux2_1 _10962_ (.A0(\shift_storage.storage [652]),
    .A1(\shift_storage.storage [651]),
    .S(net299),
    .X(_04546_));
 sg13g2_and2_1 _10963_ (.A(net300),
    .B(_04546_),
    .X(_01316_));
 sg13g2_mux2_1 _10964_ (.A0(\shift_storage.storage [653]),
    .A1(\shift_storage.storage [652]),
    .S(_04542_),
    .X(_04547_));
 sg13g2_and2_1 _10965_ (.A(net300),
    .B(_04547_),
    .X(_01317_));
 sg13g2_mux2_1 _10966_ (.A0(\shift_storage.storage [654]),
    .A1(\shift_storage.storage [653]),
    .S(_04542_),
    .X(_04548_));
 sg13g2_and2_1 _10967_ (.A(_04537_),
    .B(_04548_),
    .X(_01318_));
 sg13g2_buf_1 _10968_ (.A(net403),
    .X(_04549_));
 sg13g2_mux2_1 _10969_ (.A0(\shift_storage.storage [655]),
    .A1(\shift_storage.storage [654]),
    .S(net299),
    .X(_04550_));
 sg13g2_and2_1 _10970_ (.A(net298),
    .B(_04550_),
    .X(_01319_));
 sg13g2_mux2_1 _10971_ (.A0(\shift_storage.storage [656]),
    .A1(\shift_storage.storage [655]),
    .S(net299),
    .X(_04551_));
 sg13g2_and2_1 _10972_ (.A(net298),
    .B(_04551_),
    .X(_01320_));
 sg13g2_mux2_1 _10973_ (.A0(\shift_storage.storage [657]),
    .A1(\shift_storage.storage [656]),
    .S(net299),
    .X(_04552_));
 sg13g2_and2_1 _10974_ (.A(net298),
    .B(_04552_),
    .X(_01321_));
 sg13g2_mux2_1 _10975_ (.A0(\shift_storage.storage [658]),
    .A1(\shift_storage.storage [657]),
    .S(net299),
    .X(_04553_));
 sg13g2_and2_1 _10976_ (.A(_04549_),
    .B(_04553_),
    .X(_01322_));
 sg13g2_buf_1 _10977_ (.A(net404),
    .X(_04554_));
 sg13g2_mux2_1 _10978_ (.A0(\shift_storage.storage [659]),
    .A1(\shift_storage.storage [658]),
    .S(_04554_),
    .X(_04555_));
 sg13g2_and2_1 _10979_ (.A(net298),
    .B(_04555_),
    .X(_01323_));
 sg13g2_mux2_1 _10980_ (.A0(\shift_storage.storage [65]),
    .A1(\shift_storage.storage [64]),
    .S(_04554_),
    .X(_04556_));
 sg13g2_and2_1 _10981_ (.A(_04549_),
    .B(_04556_),
    .X(_01324_));
 sg13g2_mux2_1 _10982_ (.A0(\shift_storage.storage [660]),
    .A1(\shift_storage.storage [659]),
    .S(net297),
    .X(_04557_));
 sg13g2_and2_1 _10983_ (.A(net298),
    .B(_04557_),
    .X(_01325_));
 sg13g2_mux2_1 _10984_ (.A0(\shift_storage.storage [661]),
    .A1(\shift_storage.storage [660]),
    .S(net297),
    .X(_04558_));
 sg13g2_and2_1 _10985_ (.A(net298),
    .B(_04558_),
    .X(_01326_));
 sg13g2_mux2_1 _10986_ (.A0(\shift_storage.storage [662]),
    .A1(\shift_storage.storage [661]),
    .S(net297),
    .X(_04559_));
 sg13g2_and2_1 _10987_ (.A(net298),
    .B(_04559_),
    .X(_01327_));
 sg13g2_mux2_1 _10988_ (.A0(\shift_storage.storage [663]),
    .A1(\shift_storage.storage [662]),
    .S(net297),
    .X(_04560_));
 sg13g2_and2_1 _10989_ (.A(net298),
    .B(_04560_),
    .X(_01328_));
 sg13g2_buf_1 _10990_ (.A(net403),
    .X(_04561_));
 sg13g2_mux2_1 _10991_ (.A0(\shift_storage.storage [664]),
    .A1(\shift_storage.storage [663]),
    .S(net297),
    .X(_04562_));
 sg13g2_and2_1 _10992_ (.A(net296),
    .B(_04562_),
    .X(_01329_));
 sg13g2_mux2_1 _10993_ (.A0(\shift_storage.storage [665]),
    .A1(\shift_storage.storage [664]),
    .S(net297),
    .X(_04563_));
 sg13g2_and2_1 _10994_ (.A(net296),
    .B(_04563_),
    .X(_01330_));
 sg13g2_mux2_1 _10995_ (.A0(\shift_storage.storage [666]),
    .A1(\shift_storage.storage [665]),
    .S(net297),
    .X(_04564_));
 sg13g2_and2_1 _10996_ (.A(net296),
    .B(_04564_),
    .X(_01331_));
 sg13g2_mux2_1 _10997_ (.A0(\shift_storage.storage [667]),
    .A1(\shift_storage.storage [666]),
    .S(net297),
    .X(_04565_));
 sg13g2_and2_1 _10998_ (.A(net296),
    .B(_04565_),
    .X(_01332_));
 sg13g2_buf_1 _10999_ (.A(net404),
    .X(_04566_));
 sg13g2_mux2_1 _11000_ (.A0(\shift_storage.storage [668]),
    .A1(\shift_storage.storage [667]),
    .S(net295),
    .X(_04567_));
 sg13g2_and2_1 _11001_ (.A(net296),
    .B(_04567_),
    .X(_01333_));
 sg13g2_mux2_1 _11002_ (.A0(\shift_storage.storage [669]),
    .A1(\shift_storage.storage [668]),
    .S(_04566_),
    .X(_04568_));
 sg13g2_and2_1 _11003_ (.A(_04561_),
    .B(_04568_),
    .X(_01334_));
 sg13g2_mux2_1 _11004_ (.A0(\shift_storage.storage [66]),
    .A1(\shift_storage.storage [65]),
    .S(_04566_),
    .X(_04569_));
 sg13g2_and2_1 _11005_ (.A(_04561_),
    .B(_04569_),
    .X(_01335_));
 sg13g2_mux2_1 _11006_ (.A0(\shift_storage.storage [670]),
    .A1(\shift_storage.storage [669]),
    .S(net295),
    .X(_04570_));
 sg13g2_and2_1 _11007_ (.A(net296),
    .B(_04570_),
    .X(_01336_));
 sg13g2_mux2_1 _11008_ (.A0(\shift_storage.storage [671]),
    .A1(\shift_storage.storage [670]),
    .S(net295),
    .X(_04571_));
 sg13g2_and2_1 _11009_ (.A(net296),
    .B(_04571_),
    .X(_01337_));
 sg13g2_mux2_1 _11010_ (.A0(\shift_storage.storage [672]),
    .A1(\shift_storage.storage [671]),
    .S(net295),
    .X(_04572_));
 sg13g2_and2_1 _11011_ (.A(net296),
    .B(_04572_),
    .X(_01338_));
 sg13g2_buf_1 _11012_ (.A(net403),
    .X(_04573_));
 sg13g2_mux2_1 _11013_ (.A0(\shift_storage.storage [673]),
    .A1(\shift_storage.storage [672]),
    .S(net295),
    .X(_04574_));
 sg13g2_and2_1 _11014_ (.A(net294),
    .B(_04574_),
    .X(_01339_));
 sg13g2_mux2_1 _11015_ (.A0(\shift_storage.storage [674]),
    .A1(\shift_storage.storage [673]),
    .S(net295),
    .X(_04575_));
 sg13g2_and2_1 _11016_ (.A(net294),
    .B(_04575_),
    .X(_01340_));
 sg13g2_mux2_1 _11017_ (.A0(\shift_storage.storage [675]),
    .A1(\shift_storage.storage [674]),
    .S(net295),
    .X(_04576_));
 sg13g2_and2_1 _11018_ (.A(net294),
    .B(_04576_),
    .X(_01341_));
 sg13g2_mux2_1 _11019_ (.A0(\shift_storage.storage [676]),
    .A1(\shift_storage.storage [675]),
    .S(net295),
    .X(_04577_));
 sg13g2_and2_1 _11020_ (.A(net294),
    .B(_04577_),
    .X(_01342_));
 sg13g2_buf_1 _11021_ (.A(net404),
    .X(_04578_));
 sg13g2_mux2_1 _11022_ (.A0(\shift_storage.storage [677]),
    .A1(\shift_storage.storage [676]),
    .S(net293),
    .X(_04579_));
 sg13g2_and2_1 _11023_ (.A(net294),
    .B(_04579_),
    .X(_01343_));
 sg13g2_mux2_1 _11024_ (.A0(\shift_storage.storage [678]),
    .A1(\shift_storage.storage [677]),
    .S(net293),
    .X(_04580_));
 sg13g2_and2_1 _11025_ (.A(net294),
    .B(_04580_),
    .X(_01344_));
 sg13g2_mux2_1 _11026_ (.A0(\shift_storage.storage [679]),
    .A1(\shift_storage.storage [678]),
    .S(net293),
    .X(_04581_));
 sg13g2_and2_1 _11027_ (.A(net294),
    .B(_04581_),
    .X(_01345_));
 sg13g2_mux2_1 _11028_ (.A0(\shift_storage.storage [67]),
    .A1(\shift_storage.storage [66]),
    .S(net293),
    .X(_04582_));
 sg13g2_and2_1 _11029_ (.A(net294),
    .B(_04582_),
    .X(_01346_));
 sg13g2_mux2_1 _11030_ (.A0(\shift_storage.storage [680]),
    .A1(\shift_storage.storage [679]),
    .S(net293),
    .X(_04583_));
 sg13g2_and2_1 _11031_ (.A(_04573_),
    .B(_04583_),
    .X(_01347_));
 sg13g2_mux2_1 _11032_ (.A0(\shift_storage.storage [681]),
    .A1(\shift_storage.storage [680]),
    .S(net293),
    .X(_04584_));
 sg13g2_and2_1 _11033_ (.A(_04573_),
    .B(_04584_),
    .X(_01348_));
 sg13g2_buf_1 _11034_ (.A(net403),
    .X(_04585_));
 sg13g2_mux2_1 _11035_ (.A0(\shift_storage.storage [682]),
    .A1(\shift_storage.storage [681]),
    .S(net293),
    .X(_04586_));
 sg13g2_and2_1 _11036_ (.A(net292),
    .B(_04586_),
    .X(_01349_));
 sg13g2_mux2_1 _11037_ (.A0(\shift_storage.storage [683]),
    .A1(\shift_storage.storage [682]),
    .S(net293),
    .X(_04587_));
 sg13g2_and2_1 _11038_ (.A(net292),
    .B(_04587_),
    .X(_01350_));
 sg13g2_mux2_1 _11039_ (.A0(\shift_storage.storage [684]),
    .A1(\shift_storage.storage [683]),
    .S(_04578_),
    .X(_04588_));
 sg13g2_and2_1 _11040_ (.A(net292),
    .B(_04588_),
    .X(_01351_));
 sg13g2_mux2_1 _11041_ (.A0(\shift_storage.storage [685]),
    .A1(\shift_storage.storage [684]),
    .S(_04578_),
    .X(_04589_));
 sg13g2_and2_1 _11042_ (.A(net292),
    .B(_04589_),
    .X(_01352_));
 sg13g2_buf_1 _11043_ (.A(net404),
    .X(_04590_));
 sg13g2_mux2_1 _11044_ (.A0(\shift_storage.storage [686]),
    .A1(\shift_storage.storage [685]),
    .S(net291),
    .X(_04591_));
 sg13g2_and2_1 _11045_ (.A(net292),
    .B(_04591_),
    .X(_01353_));
 sg13g2_mux2_1 _11046_ (.A0(\shift_storage.storage [687]),
    .A1(\shift_storage.storage [686]),
    .S(net291),
    .X(_04592_));
 sg13g2_and2_1 _11047_ (.A(net292),
    .B(_04592_),
    .X(_01354_));
 sg13g2_mux2_1 _11048_ (.A0(\shift_storage.storage [688]),
    .A1(\shift_storage.storage [687]),
    .S(net291),
    .X(_04593_));
 sg13g2_and2_1 _11049_ (.A(net292),
    .B(_04593_),
    .X(_01355_));
 sg13g2_mux2_1 _11050_ (.A0(\shift_storage.storage [689]),
    .A1(\shift_storage.storage [688]),
    .S(net291),
    .X(_04594_));
 sg13g2_and2_1 _11051_ (.A(_04585_),
    .B(_04594_),
    .X(_01356_));
 sg13g2_mux2_1 _11052_ (.A0(\shift_storage.storage [68]),
    .A1(\shift_storage.storage [67]),
    .S(net291),
    .X(_04595_));
 sg13g2_and2_1 _11053_ (.A(net292),
    .B(_04595_),
    .X(_01357_));
 sg13g2_mux2_1 _11054_ (.A0(\shift_storage.storage [690]),
    .A1(\shift_storage.storage [689]),
    .S(net291),
    .X(_04596_));
 sg13g2_and2_1 _11055_ (.A(_04585_),
    .B(_04596_),
    .X(_01358_));
 sg13g2_buf_1 _11056_ (.A(net403),
    .X(_04597_));
 sg13g2_mux2_1 _11057_ (.A0(\shift_storage.storage [691]),
    .A1(\shift_storage.storage [690]),
    .S(net291),
    .X(_04598_));
 sg13g2_and2_1 _11058_ (.A(net290),
    .B(_04598_),
    .X(_01359_));
 sg13g2_mux2_1 _11059_ (.A0(\shift_storage.storage [692]),
    .A1(\shift_storage.storage [691]),
    .S(net291),
    .X(_04599_));
 sg13g2_and2_1 _11060_ (.A(net290),
    .B(_04599_),
    .X(_01360_));
 sg13g2_mux2_1 _11061_ (.A0(\shift_storage.storage [693]),
    .A1(\shift_storage.storage [692]),
    .S(_04590_),
    .X(_04600_));
 sg13g2_and2_1 _11062_ (.A(net290),
    .B(_04600_),
    .X(_01361_));
 sg13g2_mux2_1 _11063_ (.A0(\shift_storage.storage [694]),
    .A1(\shift_storage.storage [693]),
    .S(_04590_),
    .X(_04601_));
 sg13g2_and2_1 _11064_ (.A(net290),
    .B(_04601_),
    .X(_01362_));
 sg13g2_buf_1 _11065_ (.A(_04516_),
    .X(_04602_));
 sg13g2_mux2_1 _11066_ (.A0(\shift_storage.storage [695]),
    .A1(\shift_storage.storage [694]),
    .S(net289),
    .X(_04603_));
 sg13g2_and2_1 _11067_ (.A(net290),
    .B(_04603_),
    .X(_01363_));
 sg13g2_mux2_1 _11068_ (.A0(\shift_storage.storage [696]),
    .A1(\shift_storage.storage [695]),
    .S(net289),
    .X(_04604_));
 sg13g2_and2_1 _11069_ (.A(net290),
    .B(_04604_),
    .X(_01364_));
 sg13g2_mux2_1 _11070_ (.A0(\shift_storage.storage [697]),
    .A1(\shift_storage.storage [696]),
    .S(net289),
    .X(_04605_));
 sg13g2_and2_1 _11071_ (.A(net290),
    .B(_04605_),
    .X(_01365_));
 sg13g2_mux2_1 _11072_ (.A0(\shift_storage.storage [698]),
    .A1(\shift_storage.storage [697]),
    .S(net289),
    .X(_04606_));
 sg13g2_and2_1 _11073_ (.A(net290),
    .B(_04606_),
    .X(_01366_));
 sg13g2_mux2_1 _11074_ (.A0(\shift_storage.storage [699]),
    .A1(\shift_storage.storage [698]),
    .S(net289),
    .X(_04607_));
 sg13g2_and2_1 _11075_ (.A(_04597_),
    .B(_04607_),
    .X(_01367_));
 sg13g2_mux2_1 _11076_ (.A0(\shift_storage.storage [69]),
    .A1(\shift_storage.storage [68]),
    .S(net289),
    .X(_04608_));
 sg13g2_and2_1 _11077_ (.A(_04597_),
    .B(_04608_),
    .X(_01368_));
 sg13g2_buf_1 _11078_ (.A(net403),
    .X(_04609_));
 sg13g2_mux2_1 _11079_ (.A0(\shift_storage.storage [6]),
    .A1(\shift_storage.storage [5]),
    .S(net289),
    .X(_04610_));
 sg13g2_and2_1 _11080_ (.A(net288),
    .B(_04610_),
    .X(_01369_));
 sg13g2_mux2_1 _11081_ (.A0(\shift_storage.storage [700]),
    .A1(\shift_storage.storage [699]),
    .S(net289),
    .X(_04611_));
 sg13g2_and2_1 _11082_ (.A(net288),
    .B(_04611_),
    .X(_01370_));
 sg13g2_mux2_1 _11083_ (.A0(\shift_storage.storage [701]),
    .A1(\shift_storage.storage [700]),
    .S(_04602_),
    .X(_04612_));
 sg13g2_and2_1 _11084_ (.A(_04609_),
    .B(_04612_),
    .X(_01371_));
 sg13g2_mux2_1 _11085_ (.A0(\shift_storage.storage [702]),
    .A1(\shift_storage.storage [701]),
    .S(_04602_),
    .X(_04613_));
 sg13g2_and2_1 _11086_ (.A(_04609_),
    .B(_04613_),
    .X(_01372_));
 sg13g2_buf_1 _11087_ (.A(_04516_),
    .X(_04614_));
 sg13g2_mux2_1 _11088_ (.A0(\shift_storage.storage [703]),
    .A1(\shift_storage.storage [702]),
    .S(net287),
    .X(_04615_));
 sg13g2_and2_1 _11089_ (.A(net288),
    .B(_04615_),
    .X(_01373_));
 sg13g2_mux2_1 _11090_ (.A0(\shift_storage.storage [704]),
    .A1(\shift_storage.storage [703]),
    .S(net287),
    .X(_04616_));
 sg13g2_and2_1 _11091_ (.A(net288),
    .B(_04616_),
    .X(_01374_));
 sg13g2_mux2_1 _11092_ (.A0(\shift_storage.storage [705]),
    .A1(\shift_storage.storage [704]),
    .S(_04614_),
    .X(_04617_));
 sg13g2_and2_1 _11093_ (.A(net288),
    .B(_04617_),
    .X(_01375_));
 sg13g2_mux2_1 _11094_ (.A0(\shift_storage.storage [706]),
    .A1(\shift_storage.storage [705]),
    .S(net287),
    .X(_04618_));
 sg13g2_and2_1 _11095_ (.A(net288),
    .B(_04618_),
    .X(_01376_));
 sg13g2_mux2_1 _11096_ (.A0(\shift_storage.storage [707]),
    .A1(\shift_storage.storage [706]),
    .S(net287),
    .X(_04619_));
 sg13g2_and2_1 _11097_ (.A(net288),
    .B(_04619_),
    .X(_01377_));
 sg13g2_mux2_1 _11098_ (.A0(\shift_storage.storage [708]),
    .A1(\shift_storage.storage [707]),
    .S(net287),
    .X(_04620_));
 sg13g2_and2_1 _11099_ (.A(net288),
    .B(_04620_),
    .X(_01378_));
 sg13g2_buf_1 _11100_ (.A(_04524_),
    .X(_04621_));
 sg13g2_mux2_1 _11101_ (.A0(\shift_storage.storage [709]),
    .A1(\shift_storage.storage [708]),
    .S(net287),
    .X(_04622_));
 sg13g2_and2_1 _11102_ (.A(net286),
    .B(_04622_),
    .X(_01379_));
 sg13g2_mux2_1 _11103_ (.A0(\shift_storage.storage [70]),
    .A1(\shift_storage.storage [69]),
    .S(net287),
    .X(_04623_));
 sg13g2_and2_1 _11104_ (.A(net286),
    .B(_04623_),
    .X(_01380_));
 sg13g2_mux2_1 _11105_ (.A0(\shift_storage.storage [710]),
    .A1(\shift_storage.storage [709]),
    .S(net287),
    .X(_04624_));
 sg13g2_and2_1 _11106_ (.A(_04621_),
    .B(_04624_),
    .X(_01381_));
 sg13g2_mux2_1 _11107_ (.A0(\shift_storage.storage [711]),
    .A1(\shift_storage.storage [710]),
    .S(_04614_),
    .X(_04625_));
 sg13g2_and2_1 _11108_ (.A(_04621_),
    .B(_04625_),
    .X(_01382_));
 sg13g2_buf_1 _11109_ (.A(net404),
    .X(_04626_));
 sg13g2_mux2_1 _11110_ (.A0(\shift_storage.storage [712]),
    .A1(\shift_storage.storage [711]),
    .S(net285),
    .X(_04627_));
 sg13g2_and2_1 _11111_ (.A(net286),
    .B(_04627_),
    .X(_01383_));
 sg13g2_mux2_1 _11112_ (.A0(\shift_storage.storage [713]),
    .A1(\shift_storage.storage [712]),
    .S(net285),
    .X(_04628_));
 sg13g2_and2_1 _11113_ (.A(net286),
    .B(_04628_),
    .X(_01384_));
 sg13g2_mux2_1 _11114_ (.A0(\shift_storage.storage [714]),
    .A1(\shift_storage.storage [713]),
    .S(net285),
    .X(_04629_));
 sg13g2_and2_1 _11115_ (.A(net286),
    .B(_04629_),
    .X(_01385_));
 sg13g2_mux2_1 _11116_ (.A0(\shift_storage.storage [715]),
    .A1(\shift_storage.storage [714]),
    .S(net285),
    .X(_04630_));
 sg13g2_and2_1 _11117_ (.A(net286),
    .B(_04630_),
    .X(_01386_));
 sg13g2_mux2_1 _11118_ (.A0(\shift_storage.storage [716]),
    .A1(\shift_storage.storage [715]),
    .S(_04626_),
    .X(_04631_));
 sg13g2_and2_1 _11119_ (.A(net286),
    .B(_04631_),
    .X(_01387_));
 sg13g2_mux2_1 _11120_ (.A0(\shift_storage.storage [717]),
    .A1(\shift_storage.storage [716]),
    .S(_04626_),
    .X(_04632_));
 sg13g2_and2_1 _11121_ (.A(net286),
    .B(_04632_),
    .X(_01388_));
 sg13g2_buf_1 _11122_ (.A(_04524_),
    .X(_04633_));
 sg13g2_mux2_1 _11123_ (.A0(\shift_storage.storage [718]),
    .A1(\shift_storage.storage [717]),
    .S(net285),
    .X(_04634_));
 sg13g2_and2_1 _11124_ (.A(net284),
    .B(_04634_),
    .X(_01389_));
 sg13g2_mux2_1 _11125_ (.A0(\shift_storage.storage [719]),
    .A1(\shift_storage.storage [718]),
    .S(net285),
    .X(_04635_));
 sg13g2_and2_1 _11126_ (.A(net284),
    .B(_04635_),
    .X(_01390_));
 sg13g2_mux2_1 _11127_ (.A0(\shift_storage.storage [71]),
    .A1(\shift_storage.storage [70]),
    .S(net285),
    .X(_04636_));
 sg13g2_and2_1 _11128_ (.A(_04633_),
    .B(_04636_),
    .X(_01391_));
 sg13g2_mux2_1 _11129_ (.A0(\shift_storage.storage [720]),
    .A1(\shift_storage.storage [719]),
    .S(net285),
    .X(_04637_));
 sg13g2_and2_1 _11130_ (.A(_04633_),
    .B(_04637_),
    .X(_01392_));
 sg13g2_buf_1 _11131_ (.A(_03058_),
    .X(_04638_));
 sg13g2_buf_1 _11132_ (.A(net402),
    .X(_04639_));
 sg13g2_mux2_1 _11133_ (.A0(\shift_storage.storage [721]),
    .A1(\shift_storage.storage [720]),
    .S(net283),
    .X(_04640_));
 sg13g2_and2_1 _11134_ (.A(net284),
    .B(_04640_),
    .X(_01393_));
 sg13g2_mux2_1 _11135_ (.A0(\shift_storage.storage [722]),
    .A1(\shift_storage.storage [721]),
    .S(net283),
    .X(_04641_));
 sg13g2_and2_1 _11136_ (.A(net284),
    .B(_04641_),
    .X(_01394_));
 sg13g2_mux2_1 _11137_ (.A0(\shift_storage.storage [723]),
    .A1(\shift_storage.storage [722]),
    .S(net283),
    .X(_04642_));
 sg13g2_and2_1 _11138_ (.A(net284),
    .B(_04642_),
    .X(_01395_));
 sg13g2_mux2_1 _11139_ (.A0(\shift_storage.storage [724]),
    .A1(\shift_storage.storage [723]),
    .S(net283),
    .X(_04643_));
 sg13g2_and2_1 _11140_ (.A(net284),
    .B(_04643_),
    .X(_01396_));
 sg13g2_mux2_1 _11141_ (.A0(\shift_storage.storage [725]),
    .A1(\shift_storage.storage [724]),
    .S(net283),
    .X(_04644_));
 sg13g2_and2_1 _11142_ (.A(net284),
    .B(_04644_),
    .X(_01397_));
 sg13g2_mux2_1 _11143_ (.A0(\shift_storage.storage [726]),
    .A1(\shift_storage.storage [725]),
    .S(net283),
    .X(_04645_));
 sg13g2_and2_1 _11144_ (.A(net284),
    .B(_04645_),
    .X(_01398_));
 sg13g2_buf_1 _11145_ (.A(net494),
    .X(_04646_));
 sg13g2_buf_1 _11146_ (.A(net401),
    .X(_04647_));
 sg13g2_mux2_1 _11147_ (.A0(\shift_storage.storage [727]),
    .A1(\shift_storage.storage [726]),
    .S(net283),
    .X(_04648_));
 sg13g2_and2_1 _11148_ (.A(net282),
    .B(_04648_),
    .X(_01399_));
 sg13g2_mux2_1 _11149_ (.A0(\shift_storage.storage [728]),
    .A1(\shift_storage.storage [727]),
    .S(net283),
    .X(_04649_));
 sg13g2_and2_1 _11150_ (.A(net282),
    .B(_04649_),
    .X(_01400_));
 sg13g2_mux2_1 _11151_ (.A0(\shift_storage.storage [729]),
    .A1(\shift_storage.storage [728]),
    .S(_04639_),
    .X(_04650_));
 sg13g2_and2_1 _11152_ (.A(net282),
    .B(_04650_),
    .X(_01401_));
 sg13g2_mux2_1 _11153_ (.A0(\shift_storage.storage [72]),
    .A1(\shift_storage.storage [71]),
    .S(_04639_),
    .X(_04651_));
 sg13g2_and2_1 _11154_ (.A(net282),
    .B(_04651_),
    .X(_01402_));
 sg13g2_buf_1 _11155_ (.A(net402),
    .X(_04652_));
 sg13g2_mux2_1 _11156_ (.A0(\shift_storage.storage [730]),
    .A1(\shift_storage.storage [729]),
    .S(net281),
    .X(_04653_));
 sg13g2_and2_1 _11157_ (.A(net282),
    .B(_04653_),
    .X(_01403_));
 sg13g2_mux2_1 _11158_ (.A0(\shift_storage.storage [731]),
    .A1(\shift_storage.storage [730]),
    .S(net281),
    .X(_04654_));
 sg13g2_and2_1 _11159_ (.A(net282),
    .B(_04654_),
    .X(_01404_));
 sg13g2_mux2_1 _11160_ (.A0(\shift_storage.storage [732]),
    .A1(\shift_storage.storage [731]),
    .S(net281),
    .X(_04655_));
 sg13g2_and2_1 _11161_ (.A(net282),
    .B(_04655_),
    .X(_01405_));
 sg13g2_mux2_1 _11162_ (.A0(\shift_storage.storage [733]),
    .A1(\shift_storage.storage [732]),
    .S(net281),
    .X(_04656_));
 sg13g2_and2_1 _11163_ (.A(net282),
    .B(_04656_),
    .X(_01406_));
 sg13g2_mux2_1 _11164_ (.A0(\shift_storage.storage [734]),
    .A1(\shift_storage.storage [733]),
    .S(net281),
    .X(_04657_));
 sg13g2_and2_1 _11165_ (.A(_04647_),
    .B(_04657_),
    .X(_01407_));
 sg13g2_mux2_1 _11166_ (.A0(\shift_storage.storage [735]),
    .A1(\shift_storage.storage [734]),
    .S(net281),
    .X(_04658_));
 sg13g2_and2_1 _11167_ (.A(_04647_),
    .B(_04658_),
    .X(_01408_));
 sg13g2_buf_1 _11168_ (.A(net401),
    .X(_04659_));
 sg13g2_mux2_1 _11169_ (.A0(\shift_storage.storage [736]),
    .A1(\shift_storage.storage [735]),
    .S(net281),
    .X(_04660_));
 sg13g2_and2_1 _11170_ (.A(net280),
    .B(_04660_),
    .X(_01409_));
 sg13g2_mux2_1 _11171_ (.A0(\shift_storage.storage [737]),
    .A1(\shift_storage.storage [736]),
    .S(net281),
    .X(_04661_));
 sg13g2_and2_1 _11172_ (.A(net280),
    .B(_04661_),
    .X(_01410_));
 sg13g2_mux2_1 _11173_ (.A0(\shift_storage.storage [738]),
    .A1(\shift_storage.storage [737]),
    .S(_04652_),
    .X(_04662_));
 sg13g2_and2_1 _11174_ (.A(net280),
    .B(_04662_),
    .X(_01411_));
 sg13g2_mux2_1 _11175_ (.A0(\shift_storage.storage [739]),
    .A1(\shift_storage.storage [738]),
    .S(_04652_),
    .X(_04663_));
 sg13g2_and2_1 _11176_ (.A(_04659_),
    .B(_04663_),
    .X(_01412_));
 sg13g2_buf_1 _11177_ (.A(net402),
    .X(_04664_));
 sg13g2_mux2_1 _11178_ (.A0(\shift_storage.storage [73]),
    .A1(\shift_storage.storage [72]),
    .S(net279),
    .X(_04665_));
 sg13g2_and2_1 _11179_ (.A(_04659_),
    .B(_04665_),
    .X(_01413_));
 sg13g2_mux2_1 _11180_ (.A0(\shift_storage.storage [740]),
    .A1(\shift_storage.storage [739]),
    .S(net279),
    .X(_04666_));
 sg13g2_and2_1 _11181_ (.A(net280),
    .B(_04666_),
    .X(_01414_));
 sg13g2_mux2_1 _11182_ (.A0(\shift_storage.storage [741]),
    .A1(\shift_storage.storage [740]),
    .S(net279),
    .X(_04667_));
 sg13g2_and2_1 _11183_ (.A(net280),
    .B(_04667_),
    .X(_01415_));
 sg13g2_mux2_1 _11184_ (.A0(\shift_storage.storage [742]),
    .A1(\shift_storage.storage [741]),
    .S(net279),
    .X(_04668_));
 sg13g2_and2_1 _11185_ (.A(net280),
    .B(_04668_),
    .X(_01416_));
 sg13g2_mux2_1 _11186_ (.A0(\shift_storage.storage [743]),
    .A1(\shift_storage.storage [742]),
    .S(net279),
    .X(_04669_));
 sg13g2_and2_1 _11187_ (.A(net280),
    .B(_04669_),
    .X(_01417_));
 sg13g2_mux2_1 _11188_ (.A0(\shift_storage.storage [744]),
    .A1(\shift_storage.storage [743]),
    .S(net279),
    .X(_04670_));
 sg13g2_and2_1 _11189_ (.A(net280),
    .B(_04670_),
    .X(_01418_));
 sg13g2_buf_1 _11190_ (.A(net401),
    .X(_04671_));
 sg13g2_mux2_1 _11191_ (.A0(\shift_storage.storage [745]),
    .A1(\shift_storage.storage [744]),
    .S(net279),
    .X(_04672_));
 sg13g2_and2_1 _11192_ (.A(net278),
    .B(_04672_),
    .X(_01419_));
 sg13g2_mux2_1 _11193_ (.A0(\shift_storage.storage [746]),
    .A1(\shift_storage.storage [745]),
    .S(net279),
    .X(_04673_));
 sg13g2_and2_1 _11194_ (.A(net278),
    .B(_04673_),
    .X(_01420_));
 sg13g2_mux2_1 _11195_ (.A0(\shift_storage.storage [747]),
    .A1(\shift_storage.storage [746]),
    .S(_04664_),
    .X(_04674_));
 sg13g2_and2_1 _11196_ (.A(net278),
    .B(_04674_),
    .X(_01421_));
 sg13g2_mux2_1 _11197_ (.A0(\shift_storage.storage [748]),
    .A1(\shift_storage.storage [747]),
    .S(_04664_),
    .X(_04675_));
 sg13g2_and2_1 _11198_ (.A(net278),
    .B(_04675_),
    .X(_01422_));
 sg13g2_buf_1 _11199_ (.A(net402),
    .X(_04676_));
 sg13g2_mux2_1 _11200_ (.A0(\shift_storage.storage [749]),
    .A1(\shift_storage.storage [748]),
    .S(net277),
    .X(_04677_));
 sg13g2_and2_1 _11201_ (.A(net278),
    .B(_04677_),
    .X(_01423_));
 sg13g2_mux2_1 _11202_ (.A0(\shift_storage.storage [74]),
    .A1(\shift_storage.storage [73]),
    .S(net277),
    .X(_04678_));
 sg13g2_and2_1 _11203_ (.A(net278),
    .B(_04678_),
    .X(_01424_));
 sg13g2_mux2_1 _11204_ (.A0(\shift_storage.storage [750]),
    .A1(\shift_storage.storage [749]),
    .S(net277),
    .X(_04679_));
 sg13g2_and2_1 _11205_ (.A(net278),
    .B(_04679_),
    .X(_01425_));
 sg13g2_mux2_1 _11206_ (.A0(\shift_storage.storage [751]),
    .A1(\shift_storage.storage [750]),
    .S(net277),
    .X(_04680_));
 sg13g2_and2_1 _11207_ (.A(net278),
    .B(_04680_),
    .X(_01426_));
 sg13g2_mux2_1 _11208_ (.A0(\shift_storage.storage [752]),
    .A1(\shift_storage.storage [751]),
    .S(net277),
    .X(_04681_));
 sg13g2_and2_1 _11209_ (.A(_04671_),
    .B(_04681_),
    .X(_01427_));
 sg13g2_mux2_1 _11210_ (.A0(\shift_storage.storage [753]),
    .A1(\shift_storage.storage [752]),
    .S(net277),
    .X(_04682_));
 sg13g2_and2_1 _11211_ (.A(_04671_),
    .B(_04682_),
    .X(_01428_));
 sg13g2_buf_1 _11212_ (.A(net401),
    .X(_04683_));
 sg13g2_mux2_1 _11213_ (.A0(\shift_storage.storage [754]),
    .A1(\shift_storage.storage [753]),
    .S(net277),
    .X(_04684_));
 sg13g2_and2_1 _11214_ (.A(net276),
    .B(_04684_),
    .X(_01429_));
 sg13g2_mux2_1 _11215_ (.A0(\shift_storage.storage [755]),
    .A1(\shift_storage.storage [754]),
    .S(net277),
    .X(_04685_));
 sg13g2_and2_1 _11216_ (.A(net276),
    .B(_04685_),
    .X(_01430_));
 sg13g2_mux2_1 _11217_ (.A0(\shift_storage.storage [756]),
    .A1(\shift_storage.storage [755]),
    .S(_04676_),
    .X(_04686_));
 sg13g2_and2_1 _11218_ (.A(net276),
    .B(_04686_),
    .X(_01431_));
 sg13g2_mux2_1 _11219_ (.A0(\shift_storage.storage [757]),
    .A1(\shift_storage.storage [756]),
    .S(_04676_),
    .X(_04687_));
 sg13g2_and2_1 _11220_ (.A(net276),
    .B(_04687_),
    .X(_01432_));
 sg13g2_buf_1 _11221_ (.A(net402),
    .X(_04688_));
 sg13g2_mux2_1 _11222_ (.A0(\shift_storage.storage [758]),
    .A1(\shift_storage.storage [757]),
    .S(net275),
    .X(_04689_));
 sg13g2_and2_1 _11223_ (.A(_04683_),
    .B(_04689_),
    .X(_01433_));
 sg13g2_mux2_1 _11224_ (.A0(\shift_storage.storage [759]),
    .A1(\shift_storage.storage [758]),
    .S(net275),
    .X(_04690_));
 sg13g2_and2_1 _11225_ (.A(net276),
    .B(_04690_),
    .X(_01434_));
 sg13g2_mux2_1 _11226_ (.A0(\shift_storage.storage [75]),
    .A1(\shift_storage.storage [74]),
    .S(net275),
    .X(_04691_));
 sg13g2_and2_1 _11227_ (.A(net276),
    .B(_04691_),
    .X(_01435_));
 sg13g2_mux2_1 _11228_ (.A0(\shift_storage.storage [760]),
    .A1(\shift_storage.storage [759]),
    .S(net275),
    .X(_04692_));
 sg13g2_and2_1 _11229_ (.A(net276),
    .B(_04692_),
    .X(_01436_));
 sg13g2_mux2_1 _11230_ (.A0(\shift_storage.storage [761]),
    .A1(\shift_storage.storage [760]),
    .S(net275),
    .X(_04693_));
 sg13g2_and2_1 _11231_ (.A(net276),
    .B(_04693_),
    .X(_01437_));
 sg13g2_mux2_1 _11232_ (.A0(\shift_storage.storage [762]),
    .A1(\shift_storage.storage [761]),
    .S(net275),
    .X(_04694_));
 sg13g2_and2_1 _11233_ (.A(_04683_),
    .B(_04694_),
    .X(_01438_));
 sg13g2_buf_1 _11234_ (.A(net401),
    .X(_04695_));
 sg13g2_mux2_1 _11235_ (.A0(\shift_storage.storage [763]),
    .A1(\shift_storage.storage [762]),
    .S(net275),
    .X(_04696_));
 sg13g2_and2_1 _11236_ (.A(net274),
    .B(_04696_),
    .X(_01439_));
 sg13g2_mux2_1 _11237_ (.A0(\shift_storage.storage [764]),
    .A1(\shift_storage.storage [763]),
    .S(net275),
    .X(_04697_));
 sg13g2_and2_1 _11238_ (.A(net274),
    .B(_04697_),
    .X(_01440_));
 sg13g2_mux2_1 _11239_ (.A0(\shift_storage.storage [765]),
    .A1(\shift_storage.storage [764]),
    .S(_04688_),
    .X(_04698_));
 sg13g2_and2_1 _11240_ (.A(net274),
    .B(_04698_),
    .X(_01441_));
 sg13g2_mux2_1 _11241_ (.A0(\shift_storage.storage [766]),
    .A1(\shift_storage.storage [765]),
    .S(_04688_),
    .X(_04699_));
 sg13g2_and2_1 _11242_ (.A(net274),
    .B(_04699_),
    .X(_01442_));
 sg13g2_buf_1 _11243_ (.A(net402),
    .X(_04700_));
 sg13g2_mux2_1 _11244_ (.A0(\shift_storage.storage [767]),
    .A1(\shift_storage.storage [766]),
    .S(net273),
    .X(_04701_));
 sg13g2_and2_1 _11245_ (.A(net274),
    .B(_04701_),
    .X(_01443_));
 sg13g2_mux2_1 _11246_ (.A0(\shift_storage.storage [768]),
    .A1(\shift_storage.storage [767]),
    .S(net273),
    .X(_04702_));
 sg13g2_and2_1 _11247_ (.A(_04695_),
    .B(_04702_),
    .X(_01444_));
 sg13g2_mux2_1 _11248_ (.A0(\shift_storage.storage [769]),
    .A1(\shift_storage.storage [768]),
    .S(net273),
    .X(_04703_));
 sg13g2_and2_1 _11249_ (.A(_04695_),
    .B(_04703_),
    .X(_01445_));
 sg13g2_mux2_1 _11250_ (.A0(\shift_storage.storage [76]),
    .A1(\shift_storage.storage [75]),
    .S(net273),
    .X(_04704_));
 sg13g2_and2_1 _11251_ (.A(net274),
    .B(_04704_),
    .X(_01446_));
 sg13g2_mux2_1 _11252_ (.A0(\shift_storage.storage [770]),
    .A1(\shift_storage.storage [769]),
    .S(_04700_),
    .X(_04705_));
 sg13g2_and2_1 _11253_ (.A(net274),
    .B(_04705_),
    .X(_01447_));
 sg13g2_mux2_1 _11254_ (.A0(\shift_storage.storage [771]),
    .A1(\shift_storage.storage [770]),
    .S(_04700_),
    .X(_04706_));
 sg13g2_and2_1 _11255_ (.A(net274),
    .B(_04706_),
    .X(_01448_));
 sg13g2_buf_1 _11256_ (.A(net401),
    .X(_04707_));
 sg13g2_mux2_1 _11257_ (.A0(\shift_storage.storage [772]),
    .A1(\shift_storage.storage [771]),
    .S(net273),
    .X(_04708_));
 sg13g2_and2_1 _11258_ (.A(net272),
    .B(_04708_),
    .X(_01449_));
 sg13g2_mux2_1 _11259_ (.A0(\shift_storage.storage [773]),
    .A1(\shift_storage.storage [772]),
    .S(net273),
    .X(_04709_));
 sg13g2_and2_1 _11260_ (.A(net272),
    .B(_04709_),
    .X(_01450_));
 sg13g2_mux2_1 _11261_ (.A0(\shift_storage.storage [774]),
    .A1(\shift_storage.storage [773]),
    .S(net273),
    .X(_04710_));
 sg13g2_and2_1 _11262_ (.A(net272),
    .B(_04710_),
    .X(_01451_));
 sg13g2_mux2_1 _11263_ (.A0(\shift_storage.storage [775]),
    .A1(\shift_storage.storage [774]),
    .S(net273),
    .X(_04711_));
 sg13g2_and2_1 _11264_ (.A(_04707_),
    .B(_04711_),
    .X(_01452_));
 sg13g2_buf_1 _11265_ (.A(net402),
    .X(_04712_));
 sg13g2_mux2_1 _11266_ (.A0(\shift_storage.storage [776]),
    .A1(\shift_storage.storage [775]),
    .S(net271),
    .X(_04713_));
 sg13g2_and2_1 _11267_ (.A(net272),
    .B(_04713_),
    .X(_01453_));
 sg13g2_mux2_1 _11268_ (.A0(\shift_storage.storage [777]),
    .A1(\shift_storage.storage [776]),
    .S(net271),
    .X(_04714_));
 sg13g2_and2_1 _11269_ (.A(net272),
    .B(_04714_),
    .X(_01454_));
 sg13g2_mux2_1 _11270_ (.A0(\shift_storage.storage [778]),
    .A1(\shift_storage.storage [777]),
    .S(net271),
    .X(_04715_));
 sg13g2_and2_1 _11271_ (.A(net272),
    .B(_04715_),
    .X(_01455_));
 sg13g2_mux2_1 _11272_ (.A0(\shift_storage.storage [779]),
    .A1(\shift_storage.storage [778]),
    .S(net271),
    .X(_04716_));
 sg13g2_and2_1 _11273_ (.A(net272),
    .B(_04716_),
    .X(_01456_));
 sg13g2_mux2_1 _11274_ (.A0(\shift_storage.storage [77]),
    .A1(\shift_storage.storage [76]),
    .S(net271),
    .X(_04717_));
 sg13g2_and2_1 _11275_ (.A(_04707_),
    .B(_04717_),
    .X(_01457_));
 sg13g2_mux2_1 _11276_ (.A0(\shift_storage.storage [780]),
    .A1(\shift_storage.storage [779]),
    .S(net271),
    .X(_04718_));
 sg13g2_and2_1 _11277_ (.A(net272),
    .B(_04718_),
    .X(_01458_));
 sg13g2_buf_1 _11278_ (.A(net401),
    .X(_04719_));
 sg13g2_mux2_1 _11279_ (.A0(\shift_storage.storage [781]),
    .A1(\shift_storage.storage [780]),
    .S(net271),
    .X(_04720_));
 sg13g2_and2_1 _11280_ (.A(net270),
    .B(_04720_),
    .X(_01459_));
 sg13g2_mux2_1 _11281_ (.A0(\shift_storage.storage [782]),
    .A1(\shift_storage.storage [781]),
    .S(net271),
    .X(_04721_));
 sg13g2_and2_1 _11282_ (.A(net270),
    .B(_04721_),
    .X(_01460_));
 sg13g2_mux2_1 _11283_ (.A0(\shift_storage.storage [783]),
    .A1(\shift_storage.storage [782]),
    .S(_04712_),
    .X(_04722_));
 sg13g2_and2_1 _11284_ (.A(net270),
    .B(_04722_),
    .X(_01461_));
 sg13g2_mux2_1 _11285_ (.A0(\shift_storage.storage [784]),
    .A1(\shift_storage.storage [783]),
    .S(_04712_),
    .X(_04723_));
 sg13g2_and2_1 _11286_ (.A(net270),
    .B(_04723_),
    .X(_01462_));
 sg13g2_buf_1 _11287_ (.A(net402),
    .X(_04724_));
 sg13g2_mux2_1 _11288_ (.A0(\shift_storage.storage [785]),
    .A1(\shift_storage.storage [784]),
    .S(net269),
    .X(_04725_));
 sg13g2_and2_1 _11289_ (.A(net270),
    .B(_04725_),
    .X(_01463_));
 sg13g2_mux2_1 _11290_ (.A0(\shift_storage.storage [786]),
    .A1(\shift_storage.storage [785]),
    .S(net269),
    .X(_04726_));
 sg13g2_and2_1 _11291_ (.A(_04719_),
    .B(_04726_),
    .X(_01464_));
 sg13g2_mux2_1 _11292_ (.A0(\shift_storage.storage [787]),
    .A1(\shift_storage.storage [786]),
    .S(net269),
    .X(_04727_));
 sg13g2_and2_1 _11293_ (.A(net270),
    .B(_04727_),
    .X(_01465_));
 sg13g2_mux2_1 _11294_ (.A0(\shift_storage.storage [788]),
    .A1(\shift_storage.storage [787]),
    .S(net269),
    .X(_04728_));
 sg13g2_and2_1 _11295_ (.A(net270),
    .B(_04728_),
    .X(_01466_));
 sg13g2_mux2_1 _11296_ (.A0(\shift_storage.storage [789]),
    .A1(\shift_storage.storage [788]),
    .S(net269),
    .X(_04729_));
 sg13g2_and2_1 _11297_ (.A(net270),
    .B(_04729_),
    .X(_01467_));
 sg13g2_mux2_1 _11298_ (.A0(\shift_storage.storage [78]),
    .A1(\shift_storage.storage [77]),
    .S(net269),
    .X(_04730_));
 sg13g2_and2_1 _11299_ (.A(_04719_),
    .B(_04730_),
    .X(_01468_));
 sg13g2_buf_1 _11300_ (.A(net401),
    .X(_04731_));
 sg13g2_mux2_1 _11301_ (.A0(\shift_storage.storage [790]),
    .A1(\shift_storage.storage [789]),
    .S(net269),
    .X(_04732_));
 sg13g2_and2_1 _11302_ (.A(net268),
    .B(_04732_),
    .X(_01469_));
 sg13g2_mux2_1 _11303_ (.A0(\shift_storage.storage [791]),
    .A1(\shift_storage.storage [790]),
    .S(net269),
    .X(_04733_));
 sg13g2_and2_1 _11304_ (.A(net268),
    .B(_04733_),
    .X(_01470_));
 sg13g2_mux2_1 _11305_ (.A0(\shift_storage.storage [792]),
    .A1(\shift_storage.storage [791]),
    .S(_04724_),
    .X(_04734_));
 sg13g2_and2_1 _11306_ (.A(net268),
    .B(_04734_),
    .X(_01471_));
 sg13g2_mux2_1 _11307_ (.A0(\shift_storage.storage [793]),
    .A1(\shift_storage.storage [792]),
    .S(_04724_),
    .X(_04735_));
 sg13g2_and2_1 _11308_ (.A(net268),
    .B(_04735_),
    .X(_01472_));
 sg13g2_buf_1 _11309_ (.A(_04638_),
    .X(_04736_));
 sg13g2_mux2_1 _11310_ (.A0(\shift_storage.storage [794]),
    .A1(\shift_storage.storage [793]),
    .S(net267),
    .X(_04737_));
 sg13g2_and2_1 _11311_ (.A(net268),
    .B(_04737_),
    .X(_01473_));
 sg13g2_mux2_1 _11312_ (.A0(\shift_storage.storage [795]),
    .A1(\shift_storage.storage [794]),
    .S(net267),
    .X(_04738_));
 sg13g2_and2_1 _11313_ (.A(net268),
    .B(_04738_),
    .X(_01474_));
 sg13g2_mux2_1 _11314_ (.A0(\shift_storage.storage [796]),
    .A1(\shift_storage.storage [795]),
    .S(net267),
    .X(_04739_));
 sg13g2_and2_1 _11315_ (.A(net268),
    .B(_04739_),
    .X(_01475_));
 sg13g2_mux2_1 _11316_ (.A0(\shift_storage.storage [797]),
    .A1(\shift_storage.storage [796]),
    .S(net267),
    .X(_04740_));
 sg13g2_and2_1 _11317_ (.A(net268),
    .B(_04740_),
    .X(_01476_));
 sg13g2_mux2_1 _11318_ (.A0(\shift_storage.storage [798]),
    .A1(\shift_storage.storage [797]),
    .S(net267),
    .X(_04741_));
 sg13g2_and2_1 _11319_ (.A(_04731_),
    .B(_04741_),
    .X(_01477_));
 sg13g2_mux2_1 _11320_ (.A0(\shift_storage.storage [799]),
    .A1(\shift_storage.storage [798]),
    .S(net267),
    .X(_04742_));
 sg13g2_and2_1 _11321_ (.A(_04731_),
    .B(_04742_),
    .X(_01478_));
 sg13g2_buf_1 _11322_ (.A(_04646_),
    .X(_04743_));
 sg13g2_mux2_1 _11323_ (.A0(\shift_storage.storage [79]),
    .A1(\shift_storage.storage [78]),
    .S(net267),
    .X(_04744_));
 sg13g2_and2_1 _11324_ (.A(net266),
    .B(_04744_),
    .X(_01479_));
 sg13g2_mux2_1 _11325_ (.A0(\shift_storage.storage [7]),
    .A1(\shift_storage.storage [6]),
    .S(net267),
    .X(_04745_));
 sg13g2_and2_1 _11326_ (.A(net266),
    .B(_04745_),
    .X(_01480_));
 sg13g2_mux2_1 _11327_ (.A0(\shift_storage.storage [800]),
    .A1(\shift_storage.storage [799]),
    .S(_04736_),
    .X(_04746_));
 sg13g2_and2_1 _11328_ (.A(net266),
    .B(_04746_),
    .X(_01481_));
 sg13g2_mux2_1 _11329_ (.A0(\shift_storage.storage [801]),
    .A1(\shift_storage.storage [800]),
    .S(_04736_),
    .X(_04747_));
 sg13g2_and2_1 _11330_ (.A(net266),
    .B(_04747_),
    .X(_01482_));
 sg13g2_buf_1 _11331_ (.A(_04638_),
    .X(_04748_));
 sg13g2_mux2_1 _11332_ (.A0(\shift_storage.storage [802]),
    .A1(\shift_storage.storage [801]),
    .S(net265),
    .X(_04749_));
 sg13g2_and2_1 _11333_ (.A(net266),
    .B(_04749_),
    .X(_01483_));
 sg13g2_mux2_1 _11334_ (.A0(\shift_storage.storage [803]),
    .A1(\shift_storage.storage [802]),
    .S(net265),
    .X(_04750_));
 sg13g2_and2_1 _11335_ (.A(_04743_),
    .B(_04750_),
    .X(_01484_));
 sg13g2_mux2_1 _11336_ (.A0(\shift_storage.storage [804]),
    .A1(\shift_storage.storage [803]),
    .S(net265),
    .X(_04751_));
 sg13g2_and2_1 _11337_ (.A(_04743_),
    .B(_04751_),
    .X(_01485_));
 sg13g2_mux2_1 _11338_ (.A0(\shift_storage.storage [805]),
    .A1(\shift_storage.storage [804]),
    .S(net265),
    .X(_04752_));
 sg13g2_and2_1 _11339_ (.A(net266),
    .B(_04752_),
    .X(_01486_));
 sg13g2_mux2_1 _11340_ (.A0(\shift_storage.storage [806]),
    .A1(\shift_storage.storage [805]),
    .S(net265),
    .X(_04753_));
 sg13g2_and2_1 _11341_ (.A(net266),
    .B(_04753_),
    .X(_01487_));
 sg13g2_mux2_1 _11342_ (.A0(\shift_storage.storage [807]),
    .A1(\shift_storage.storage [806]),
    .S(net265),
    .X(_04754_));
 sg13g2_and2_1 _11343_ (.A(net266),
    .B(_04754_),
    .X(_01488_));
 sg13g2_buf_1 _11344_ (.A(_04646_),
    .X(_04755_));
 sg13g2_mux2_1 _11345_ (.A0(\shift_storage.storage [808]),
    .A1(\shift_storage.storage [807]),
    .S(net265),
    .X(_04756_));
 sg13g2_and2_1 _11346_ (.A(net264),
    .B(_04756_),
    .X(_01489_));
 sg13g2_mux2_1 _11347_ (.A0(\shift_storage.storage [809]),
    .A1(\shift_storage.storage [808]),
    .S(_04748_),
    .X(_04757_));
 sg13g2_and2_1 _11348_ (.A(net264),
    .B(_04757_),
    .X(_01490_));
 sg13g2_mux2_1 _11349_ (.A0(\shift_storage.storage [80]),
    .A1(\shift_storage.storage [79]),
    .S(_04748_),
    .X(_04758_));
 sg13g2_and2_1 _11350_ (.A(net264),
    .B(_04758_),
    .X(_01491_));
 sg13g2_mux2_1 _11351_ (.A0(\shift_storage.storage [810]),
    .A1(\shift_storage.storage [809]),
    .S(net265),
    .X(_04759_));
 sg13g2_and2_1 _11352_ (.A(net264),
    .B(_04759_),
    .X(_01492_));
 sg13g2_buf_1 _11353_ (.A(_03058_),
    .X(_04760_));
 sg13g2_buf_1 _11354_ (.A(net400),
    .X(_04761_));
 sg13g2_mux2_1 _11355_ (.A0(\shift_storage.storage [811]),
    .A1(\shift_storage.storage [810]),
    .S(net263),
    .X(_04762_));
 sg13g2_and2_1 _11356_ (.A(net264),
    .B(_04762_),
    .X(_01493_));
 sg13g2_mux2_1 _11357_ (.A0(\shift_storage.storage [812]),
    .A1(\shift_storage.storage [811]),
    .S(net263),
    .X(_04763_));
 sg13g2_and2_1 _11358_ (.A(net264),
    .B(_04763_),
    .X(_01494_));
 sg13g2_mux2_1 _11359_ (.A0(\shift_storage.storage [813]),
    .A1(\shift_storage.storage [812]),
    .S(net263),
    .X(_04764_));
 sg13g2_and2_1 _11360_ (.A(net264),
    .B(_04764_),
    .X(_01495_));
 sg13g2_mux2_1 _11361_ (.A0(\shift_storage.storage [814]),
    .A1(\shift_storage.storage [813]),
    .S(net263),
    .X(_04765_));
 sg13g2_and2_1 _11362_ (.A(net264),
    .B(_04765_),
    .X(_01496_));
 sg13g2_mux2_1 _11363_ (.A0(\shift_storage.storage [815]),
    .A1(\shift_storage.storage [814]),
    .S(net263),
    .X(_04766_));
 sg13g2_and2_1 _11364_ (.A(_04755_),
    .B(_04766_),
    .X(_01497_));
 sg13g2_mux2_1 _11365_ (.A0(\shift_storage.storage [816]),
    .A1(\shift_storage.storage [815]),
    .S(net263),
    .X(_04767_));
 sg13g2_and2_1 _11366_ (.A(_04755_),
    .B(_04767_),
    .X(_01498_));
 sg13g2_buf_1 _11367_ (.A(net494),
    .X(_04768_));
 sg13g2_buf_1 _11368_ (.A(net399),
    .X(_04769_));
 sg13g2_mux2_1 _11369_ (.A0(\shift_storage.storage [817]),
    .A1(\shift_storage.storage [816]),
    .S(net263),
    .X(_04770_));
 sg13g2_and2_1 _11370_ (.A(net262),
    .B(_04770_),
    .X(_01499_));
 sg13g2_mux2_1 _11371_ (.A0(\shift_storage.storage [818]),
    .A1(\shift_storage.storage [817]),
    .S(net263),
    .X(_04771_));
 sg13g2_and2_1 _11372_ (.A(net262),
    .B(_04771_),
    .X(_01500_));
 sg13g2_mux2_1 _11373_ (.A0(\shift_storage.storage [819]),
    .A1(\shift_storage.storage [818]),
    .S(_04761_),
    .X(_04772_));
 sg13g2_and2_1 _11374_ (.A(_04769_),
    .B(_04772_),
    .X(_01501_));
 sg13g2_mux2_1 _11375_ (.A0(\shift_storage.storage [81]),
    .A1(\shift_storage.storage [80]),
    .S(_04761_),
    .X(_04773_));
 sg13g2_and2_1 _11376_ (.A(_04769_),
    .B(_04773_),
    .X(_01502_));
 sg13g2_buf_1 _11377_ (.A(net400),
    .X(_04774_));
 sg13g2_mux2_1 _11378_ (.A0(\shift_storage.storage [820]),
    .A1(\shift_storage.storage [819]),
    .S(net261),
    .X(_04775_));
 sg13g2_and2_1 _11379_ (.A(net262),
    .B(_04775_),
    .X(_01503_));
 sg13g2_mux2_1 _11380_ (.A0(\shift_storage.storage [821]),
    .A1(\shift_storage.storage [820]),
    .S(net261),
    .X(_04776_));
 sg13g2_and2_1 _11381_ (.A(net262),
    .B(_04776_),
    .X(_01504_));
 sg13g2_mux2_1 _11382_ (.A0(\shift_storage.storage [822]),
    .A1(\shift_storage.storage [821]),
    .S(net261),
    .X(_04777_));
 sg13g2_and2_1 _11383_ (.A(net262),
    .B(_04777_),
    .X(_01505_));
 sg13g2_mux2_1 _11384_ (.A0(\shift_storage.storage [823]),
    .A1(\shift_storage.storage [822]),
    .S(_04774_),
    .X(_04778_));
 sg13g2_and2_1 _11385_ (.A(net262),
    .B(_04778_),
    .X(_01506_));
 sg13g2_mux2_1 _11386_ (.A0(\shift_storage.storage [824]),
    .A1(\shift_storage.storage [823]),
    .S(_04774_),
    .X(_04779_));
 sg13g2_and2_1 _11387_ (.A(net262),
    .B(_04779_),
    .X(_01507_));
 sg13g2_mux2_1 _11388_ (.A0(\shift_storage.storage [825]),
    .A1(\shift_storage.storage [824]),
    .S(net261),
    .X(_04780_));
 sg13g2_and2_1 _11389_ (.A(net262),
    .B(_04780_),
    .X(_01508_));
 sg13g2_buf_1 _11390_ (.A(net399),
    .X(_04781_));
 sg13g2_mux2_1 _11391_ (.A0(\shift_storage.storage [826]),
    .A1(\shift_storage.storage [825]),
    .S(net261),
    .X(_04782_));
 sg13g2_and2_1 _11392_ (.A(net260),
    .B(_04782_),
    .X(_01509_));
 sg13g2_mux2_1 _11393_ (.A0(\shift_storage.storage [827]),
    .A1(\shift_storage.storage [826]),
    .S(net261),
    .X(_04783_));
 sg13g2_and2_1 _11394_ (.A(net260),
    .B(_04783_),
    .X(_01510_));
 sg13g2_mux2_1 _11395_ (.A0(\shift_storage.storage [828]),
    .A1(\shift_storage.storage [827]),
    .S(net261),
    .X(_04784_));
 sg13g2_and2_1 _11396_ (.A(net260),
    .B(_04784_),
    .X(_01511_));
 sg13g2_mux2_1 _11397_ (.A0(\shift_storage.storage [829]),
    .A1(\shift_storage.storage [828]),
    .S(net261),
    .X(_04785_));
 sg13g2_and2_1 _11398_ (.A(net260),
    .B(_04785_),
    .X(_01512_));
 sg13g2_buf_1 _11399_ (.A(net400),
    .X(_04786_));
 sg13g2_mux2_1 _11400_ (.A0(\shift_storage.storage [82]),
    .A1(\shift_storage.storage [81]),
    .S(net259),
    .X(_04787_));
 sg13g2_and2_1 _11401_ (.A(net260),
    .B(_04787_),
    .X(_01513_));
 sg13g2_mux2_1 _11402_ (.A0(\shift_storage.storage [830]),
    .A1(\shift_storage.storage [829]),
    .S(net259),
    .X(_04788_));
 sg13g2_and2_1 _11403_ (.A(net260),
    .B(_04788_),
    .X(_01514_));
 sg13g2_mux2_1 _11404_ (.A0(\shift_storage.storage [831]),
    .A1(\shift_storage.storage [830]),
    .S(net259),
    .X(_04789_));
 sg13g2_and2_1 _11405_ (.A(net260),
    .B(_04789_),
    .X(_01515_));
 sg13g2_mux2_1 _11406_ (.A0(\shift_storage.storage [832]),
    .A1(\shift_storage.storage [831]),
    .S(net259),
    .X(_04790_));
 sg13g2_and2_1 _11407_ (.A(net260),
    .B(_04790_),
    .X(_01516_));
 sg13g2_mux2_1 _11408_ (.A0(\shift_storage.storage [833]),
    .A1(\shift_storage.storage [832]),
    .S(net259),
    .X(_04791_));
 sg13g2_and2_1 _11409_ (.A(_04781_),
    .B(_04791_),
    .X(_01517_));
 sg13g2_mux2_1 _11410_ (.A0(\shift_storage.storage [834]),
    .A1(\shift_storage.storage [833]),
    .S(net259),
    .X(_04792_));
 sg13g2_and2_1 _11411_ (.A(_04781_),
    .B(_04792_),
    .X(_01518_));
 sg13g2_buf_1 _11412_ (.A(net399),
    .X(_04793_));
 sg13g2_mux2_1 _11413_ (.A0(\shift_storage.storage [835]),
    .A1(\shift_storage.storage [834]),
    .S(_04786_),
    .X(_04794_));
 sg13g2_and2_1 _11414_ (.A(net258),
    .B(_04794_),
    .X(_01519_));
 sg13g2_mux2_1 _11415_ (.A0(\shift_storage.storage [836]),
    .A1(\shift_storage.storage [835]),
    .S(_04786_),
    .X(_04795_));
 sg13g2_and2_1 _11416_ (.A(net258),
    .B(_04795_),
    .X(_01520_));
 sg13g2_mux2_1 _11417_ (.A0(\shift_storage.storage [837]),
    .A1(\shift_storage.storage [836]),
    .S(net259),
    .X(_04796_));
 sg13g2_and2_1 _11418_ (.A(_04793_),
    .B(_04796_),
    .X(_01521_));
 sg13g2_mux2_1 _11419_ (.A0(\shift_storage.storage [838]),
    .A1(\shift_storage.storage [837]),
    .S(net259),
    .X(_04797_));
 sg13g2_and2_1 _11420_ (.A(net258),
    .B(_04797_),
    .X(_01522_));
 sg13g2_buf_1 _11421_ (.A(net400),
    .X(_04798_));
 sg13g2_mux2_1 _11422_ (.A0(\shift_storage.storage [839]),
    .A1(\shift_storage.storage [838]),
    .S(net257),
    .X(_04799_));
 sg13g2_and2_1 _11423_ (.A(net258),
    .B(_04799_),
    .X(_01523_));
 sg13g2_mux2_1 _11424_ (.A0(\shift_storage.storage [83]),
    .A1(\shift_storage.storage [82]),
    .S(_04798_),
    .X(_04800_));
 sg13g2_and2_1 _11425_ (.A(_04793_),
    .B(_04800_),
    .X(_01524_));
 sg13g2_mux2_1 _11426_ (.A0(\shift_storage.storage [840]),
    .A1(\shift_storage.storage [839]),
    .S(net257),
    .X(_04801_));
 sg13g2_and2_1 _11427_ (.A(net258),
    .B(_04801_),
    .X(_01525_));
 sg13g2_mux2_1 _11428_ (.A0(\shift_storage.storage [841]),
    .A1(\shift_storage.storage [840]),
    .S(net257),
    .X(_04802_));
 sg13g2_and2_1 _11429_ (.A(net258),
    .B(_04802_),
    .X(_01526_));
 sg13g2_mux2_1 _11430_ (.A0(\shift_storage.storage [842]),
    .A1(\shift_storage.storage [841]),
    .S(net257),
    .X(_04803_));
 sg13g2_and2_1 _11431_ (.A(net258),
    .B(_04803_),
    .X(_01527_));
 sg13g2_mux2_1 _11432_ (.A0(\shift_storage.storage [843]),
    .A1(\shift_storage.storage [842]),
    .S(net257),
    .X(_04804_));
 sg13g2_and2_1 _11433_ (.A(net258),
    .B(_04804_),
    .X(_01528_));
 sg13g2_buf_1 _11434_ (.A(net399),
    .X(_04805_));
 sg13g2_mux2_1 _11435_ (.A0(\shift_storage.storage [844]),
    .A1(\shift_storage.storage [843]),
    .S(net257),
    .X(_04806_));
 sg13g2_and2_1 _11436_ (.A(net256),
    .B(_04806_),
    .X(_01529_));
 sg13g2_mux2_1 _11437_ (.A0(\shift_storage.storage [845]),
    .A1(\shift_storage.storage [844]),
    .S(net257),
    .X(_04807_));
 sg13g2_and2_1 _11438_ (.A(net256),
    .B(_04807_),
    .X(_01530_));
 sg13g2_mux2_1 _11439_ (.A0(\shift_storage.storage [846]),
    .A1(\shift_storage.storage [845]),
    .S(net257),
    .X(_04808_));
 sg13g2_and2_1 _11440_ (.A(net256),
    .B(_04808_),
    .X(_01531_));
 sg13g2_mux2_1 _11441_ (.A0(\shift_storage.storage [847]),
    .A1(\shift_storage.storage [846]),
    .S(_04798_),
    .X(_04809_));
 sg13g2_and2_1 _11442_ (.A(net256),
    .B(_04809_),
    .X(_01532_));
 sg13g2_buf_1 _11443_ (.A(net400),
    .X(_04810_));
 sg13g2_mux2_1 _11444_ (.A0(\shift_storage.storage [848]),
    .A1(\shift_storage.storage [847]),
    .S(net255),
    .X(_04811_));
 sg13g2_and2_1 _11445_ (.A(net256),
    .B(_04811_),
    .X(_01533_));
 sg13g2_mux2_1 _11446_ (.A0(\shift_storage.storage [849]),
    .A1(\shift_storage.storage [848]),
    .S(net255),
    .X(_04812_));
 sg13g2_and2_1 _11447_ (.A(net256),
    .B(_04812_),
    .X(_01534_));
 sg13g2_mux2_1 _11448_ (.A0(\shift_storage.storage [84]),
    .A1(\shift_storage.storage [83]),
    .S(net255),
    .X(_04813_));
 sg13g2_and2_1 _11449_ (.A(net256),
    .B(_04813_),
    .X(_01535_));
 sg13g2_mux2_1 _11450_ (.A0(\shift_storage.storage [850]),
    .A1(\shift_storage.storage [849]),
    .S(net255),
    .X(_04814_));
 sg13g2_and2_1 _11451_ (.A(net256),
    .B(_04814_),
    .X(_01536_));
 sg13g2_mux2_1 _11452_ (.A0(\shift_storage.storage [851]),
    .A1(\shift_storage.storage [850]),
    .S(net255),
    .X(_04815_));
 sg13g2_and2_1 _11453_ (.A(_04805_),
    .B(_04815_),
    .X(_01537_));
 sg13g2_mux2_1 _11454_ (.A0(\shift_storage.storage [852]),
    .A1(\shift_storage.storage [851]),
    .S(net255),
    .X(_04816_));
 sg13g2_and2_1 _11455_ (.A(_04805_),
    .B(_04816_),
    .X(_01538_));
 sg13g2_buf_1 _11456_ (.A(net399),
    .X(_04817_));
 sg13g2_mux2_1 _11457_ (.A0(\shift_storage.storage [853]),
    .A1(\shift_storage.storage [852]),
    .S(net255),
    .X(_04818_));
 sg13g2_and2_1 _11458_ (.A(net254),
    .B(_04818_),
    .X(_01539_));
 sg13g2_mux2_1 _11459_ (.A0(\shift_storage.storage [854]),
    .A1(\shift_storage.storage [853]),
    .S(net255),
    .X(_04819_));
 sg13g2_and2_1 _11460_ (.A(net254),
    .B(_04819_),
    .X(_01540_));
 sg13g2_mux2_1 _11461_ (.A0(\shift_storage.storage [855]),
    .A1(\shift_storage.storage [854]),
    .S(_04810_),
    .X(_04820_));
 sg13g2_and2_1 _11462_ (.A(net254),
    .B(_04820_),
    .X(_01541_));
 sg13g2_mux2_1 _11463_ (.A0(\shift_storage.storage [856]),
    .A1(\shift_storage.storage [855]),
    .S(_04810_),
    .X(_04821_));
 sg13g2_and2_1 _11464_ (.A(net254),
    .B(_04821_),
    .X(_01542_));
 sg13g2_buf_1 _11465_ (.A(net400),
    .X(_04822_));
 sg13g2_mux2_1 _11466_ (.A0(\shift_storage.storage [857]),
    .A1(\shift_storage.storage [856]),
    .S(net253),
    .X(_04823_));
 sg13g2_and2_1 _11467_ (.A(net254),
    .B(_04823_),
    .X(_01543_));
 sg13g2_mux2_1 _11468_ (.A0(\shift_storage.storage [858]),
    .A1(\shift_storage.storage [857]),
    .S(net253),
    .X(_04824_));
 sg13g2_and2_1 _11469_ (.A(_04817_),
    .B(_04824_),
    .X(_01544_));
 sg13g2_mux2_1 _11470_ (.A0(\shift_storage.storage [859]),
    .A1(\shift_storage.storage [858]),
    .S(net253),
    .X(_04825_));
 sg13g2_and2_1 _11471_ (.A(_04817_),
    .B(_04825_),
    .X(_01545_));
 sg13g2_mux2_1 _11472_ (.A0(\shift_storage.storage [85]),
    .A1(\shift_storage.storage [84]),
    .S(net253),
    .X(_04826_));
 sg13g2_and2_1 _11473_ (.A(net254),
    .B(_04826_),
    .X(_01546_));
 sg13g2_mux2_1 _11474_ (.A0(\shift_storage.storage [860]),
    .A1(\shift_storage.storage [859]),
    .S(net253),
    .X(_04827_));
 sg13g2_and2_1 _11475_ (.A(net254),
    .B(_04827_),
    .X(_01547_));
 sg13g2_mux2_1 _11476_ (.A0(\shift_storage.storage [861]),
    .A1(\shift_storage.storage [860]),
    .S(net253),
    .X(_04828_));
 sg13g2_and2_1 _11477_ (.A(net254),
    .B(_04828_),
    .X(_01548_));
 sg13g2_buf_1 _11478_ (.A(_04768_),
    .X(_04829_));
 sg13g2_mux2_1 _11479_ (.A0(\shift_storage.storage [862]),
    .A1(\shift_storage.storage [861]),
    .S(net253),
    .X(_04830_));
 sg13g2_and2_1 _11480_ (.A(net252),
    .B(_04830_),
    .X(_01549_));
 sg13g2_mux2_1 _11481_ (.A0(\shift_storage.storage [863]),
    .A1(\shift_storage.storage [862]),
    .S(net253),
    .X(_04831_));
 sg13g2_and2_1 _11482_ (.A(net252),
    .B(_04831_),
    .X(_01550_));
 sg13g2_mux2_1 _11483_ (.A0(\shift_storage.storage [864]),
    .A1(\shift_storage.storage [863]),
    .S(_04822_),
    .X(_04832_));
 sg13g2_and2_1 _11484_ (.A(net252),
    .B(_04832_),
    .X(_01551_));
 sg13g2_mux2_1 _11485_ (.A0(\shift_storage.storage [865]),
    .A1(\shift_storage.storage [864]),
    .S(_04822_),
    .X(_04833_));
 sg13g2_and2_1 _11486_ (.A(net252),
    .B(_04833_),
    .X(_01552_));
 sg13g2_buf_1 _11487_ (.A(_04760_),
    .X(_04834_));
 sg13g2_mux2_1 _11488_ (.A0(\shift_storage.storage [866]),
    .A1(\shift_storage.storage [865]),
    .S(net251),
    .X(_04835_));
 sg13g2_and2_1 _11489_ (.A(net252),
    .B(_04835_),
    .X(_01553_));
 sg13g2_mux2_1 _11490_ (.A0(\shift_storage.storage [867]),
    .A1(\shift_storage.storage [866]),
    .S(net251),
    .X(_04836_));
 sg13g2_and2_1 _11491_ (.A(_04829_),
    .B(_04836_),
    .X(_01554_));
 sg13g2_mux2_1 _11492_ (.A0(\shift_storage.storage [868]),
    .A1(\shift_storage.storage [867]),
    .S(_04834_),
    .X(_04837_));
 sg13g2_and2_1 _11493_ (.A(_04829_),
    .B(_04837_),
    .X(_01555_));
 sg13g2_mux2_1 _11494_ (.A0(\shift_storage.storage [869]),
    .A1(\shift_storage.storage [868]),
    .S(_04834_),
    .X(_04838_));
 sg13g2_and2_1 _11495_ (.A(net252),
    .B(_04838_),
    .X(_01556_));
 sg13g2_mux2_1 _11496_ (.A0(\shift_storage.storage [86]),
    .A1(\shift_storage.storage [85]),
    .S(net251),
    .X(_04839_));
 sg13g2_and2_1 _11497_ (.A(net252),
    .B(_04839_),
    .X(_01557_));
 sg13g2_mux2_1 _11498_ (.A0(\shift_storage.storage [870]),
    .A1(\shift_storage.storage [869]),
    .S(net251),
    .X(_04840_));
 sg13g2_and2_1 _11499_ (.A(net252),
    .B(_04840_),
    .X(_01558_));
 sg13g2_buf_1 _11500_ (.A(_04768_),
    .X(_04841_));
 sg13g2_mux2_1 _11501_ (.A0(\shift_storage.storage [871]),
    .A1(\shift_storage.storage [870]),
    .S(net251),
    .X(_04842_));
 sg13g2_and2_1 _11502_ (.A(net250),
    .B(_04842_),
    .X(_01559_));
 sg13g2_mux2_1 _11503_ (.A0(\shift_storage.storage [872]),
    .A1(\shift_storage.storage [871]),
    .S(net251),
    .X(_04843_));
 sg13g2_and2_1 _11504_ (.A(net250),
    .B(_04843_),
    .X(_01560_));
 sg13g2_mux2_1 _11505_ (.A0(\shift_storage.storage [873]),
    .A1(\shift_storage.storage [872]),
    .S(net251),
    .X(_04844_));
 sg13g2_and2_1 _11506_ (.A(net250),
    .B(_04844_),
    .X(_01561_));
 sg13g2_mux2_1 _11507_ (.A0(\shift_storage.storage [874]),
    .A1(\shift_storage.storage [873]),
    .S(net251),
    .X(_04845_));
 sg13g2_and2_1 _11508_ (.A(net250),
    .B(_04845_),
    .X(_01562_));
 sg13g2_buf_1 _11509_ (.A(_04760_),
    .X(_04846_));
 sg13g2_mux2_1 _11510_ (.A0(\shift_storage.storage [875]),
    .A1(\shift_storage.storage [874]),
    .S(net249),
    .X(_04847_));
 sg13g2_and2_1 _11511_ (.A(_04841_),
    .B(_04847_),
    .X(_01563_));
 sg13g2_mux2_1 _11512_ (.A0(\shift_storage.storage [876]),
    .A1(\shift_storage.storage [875]),
    .S(_04846_),
    .X(_04848_));
 sg13g2_and2_1 _11513_ (.A(net250),
    .B(_04848_),
    .X(_01564_));
 sg13g2_mux2_1 _11514_ (.A0(\shift_storage.storage [877]),
    .A1(\shift_storage.storage [876]),
    .S(net249),
    .X(_04849_));
 sg13g2_and2_1 _11515_ (.A(net250),
    .B(_04849_),
    .X(_01565_));
 sg13g2_mux2_1 _11516_ (.A0(\shift_storage.storage [878]),
    .A1(\shift_storage.storage [877]),
    .S(net249),
    .X(_04850_));
 sg13g2_and2_1 _11517_ (.A(net250),
    .B(_04850_),
    .X(_01566_));
 sg13g2_mux2_1 _11518_ (.A0(\shift_storage.storage [879]),
    .A1(\shift_storage.storage [878]),
    .S(net249),
    .X(_04851_));
 sg13g2_and2_1 _11519_ (.A(net250),
    .B(_04851_),
    .X(_01567_));
 sg13g2_mux2_1 _11520_ (.A0(\shift_storage.storage [87]),
    .A1(\shift_storage.storage [86]),
    .S(_04846_),
    .X(_04852_));
 sg13g2_and2_1 _11521_ (.A(_04841_),
    .B(_04852_),
    .X(_01568_));
 sg13g2_buf_1 _11522_ (.A(net399),
    .X(_04853_));
 sg13g2_mux2_1 _11523_ (.A0(\shift_storage.storage [880]),
    .A1(\shift_storage.storage [879]),
    .S(net249),
    .X(_04854_));
 sg13g2_and2_1 _11524_ (.A(net248),
    .B(_04854_),
    .X(_01569_));
 sg13g2_mux2_1 _11525_ (.A0(\shift_storage.storage [881]),
    .A1(\shift_storage.storage [880]),
    .S(net249),
    .X(_04855_));
 sg13g2_and2_1 _11526_ (.A(net248),
    .B(_04855_),
    .X(_01570_));
 sg13g2_mux2_1 _11527_ (.A0(\shift_storage.storage [882]),
    .A1(\shift_storage.storage [881]),
    .S(net249),
    .X(_04856_));
 sg13g2_and2_1 _11528_ (.A(net248),
    .B(_04856_),
    .X(_01571_));
 sg13g2_mux2_1 _11529_ (.A0(\shift_storage.storage [883]),
    .A1(\shift_storage.storage [882]),
    .S(net249),
    .X(_04857_));
 sg13g2_and2_1 _11530_ (.A(net248),
    .B(_04857_),
    .X(_01572_));
 sg13g2_buf_1 _11531_ (.A(net400),
    .X(_04858_));
 sg13g2_mux2_1 _11532_ (.A0(\shift_storage.storage [884]),
    .A1(\shift_storage.storage [883]),
    .S(net247),
    .X(_04859_));
 sg13g2_and2_1 _11533_ (.A(net248),
    .B(_04859_),
    .X(_01573_));
 sg13g2_mux2_1 _11534_ (.A0(\shift_storage.storage [885]),
    .A1(\shift_storage.storage [884]),
    .S(net247),
    .X(_04860_));
 sg13g2_and2_1 _11535_ (.A(net248),
    .B(_04860_),
    .X(_01574_));
 sg13g2_mux2_1 _11536_ (.A0(\shift_storage.storage [886]),
    .A1(\shift_storage.storage [885]),
    .S(net247),
    .X(_04861_));
 sg13g2_and2_1 _11537_ (.A(net248),
    .B(_04861_),
    .X(_01575_));
 sg13g2_mux2_1 _11538_ (.A0(\shift_storage.storage [887]),
    .A1(\shift_storage.storage [886]),
    .S(net247),
    .X(_04862_));
 sg13g2_and2_1 _11539_ (.A(net248),
    .B(_04862_),
    .X(_01576_));
 sg13g2_mux2_1 _11540_ (.A0(\shift_storage.storage [888]),
    .A1(\shift_storage.storage [887]),
    .S(net247),
    .X(_04863_));
 sg13g2_and2_1 _11541_ (.A(_04853_),
    .B(_04863_),
    .X(_01577_));
 sg13g2_mux2_1 _11542_ (.A0(\shift_storage.storage [889]),
    .A1(\shift_storage.storage [888]),
    .S(net247),
    .X(_04864_));
 sg13g2_and2_1 _11543_ (.A(_04853_),
    .B(_04864_),
    .X(_01578_));
 sg13g2_buf_1 _11544_ (.A(net399),
    .X(_04865_));
 sg13g2_mux2_1 _11545_ (.A0(\shift_storage.storage [88]),
    .A1(\shift_storage.storage [87]),
    .S(net247),
    .X(_04866_));
 sg13g2_and2_1 _11546_ (.A(net246),
    .B(_04866_),
    .X(_01579_));
 sg13g2_mux2_1 _11547_ (.A0(\shift_storage.storage [890]),
    .A1(\shift_storage.storage [889]),
    .S(net247),
    .X(_04867_));
 sg13g2_and2_1 _11548_ (.A(net246),
    .B(_04867_),
    .X(_01580_));
 sg13g2_mux2_1 _11549_ (.A0(\shift_storage.storage [891]),
    .A1(\shift_storage.storage [890]),
    .S(_04858_),
    .X(_04868_));
 sg13g2_and2_1 _11550_ (.A(_04865_),
    .B(_04868_),
    .X(_01581_));
 sg13g2_mux2_1 _11551_ (.A0(\shift_storage.storage [892]),
    .A1(\shift_storage.storage [891]),
    .S(_04858_),
    .X(_04869_));
 sg13g2_and2_1 _11552_ (.A(_04865_),
    .B(_04869_),
    .X(_01582_));
 sg13g2_buf_1 _11553_ (.A(net400),
    .X(_04870_));
 sg13g2_mux2_1 _11554_ (.A0(\shift_storage.storage [893]),
    .A1(\shift_storage.storage [892]),
    .S(net245),
    .X(_04871_));
 sg13g2_and2_1 _11555_ (.A(net246),
    .B(_04871_),
    .X(_01583_));
 sg13g2_mux2_1 _11556_ (.A0(\shift_storage.storage [894]),
    .A1(\shift_storage.storage [893]),
    .S(net245),
    .X(_04872_));
 sg13g2_and2_1 _11557_ (.A(net246),
    .B(_04872_),
    .X(_01584_));
 sg13g2_mux2_1 _11558_ (.A0(\shift_storage.storage [895]),
    .A1(\shift_storage.storage [894]),
    .S(net245),
    .X(_04873_));
 sg13g2_and2_1 _11559_ (.A(net246),
    .B(_04873_),
    .X(_01585_));
 sg13g2_mux2_1 _11560_ (.A0(\shift_storage.storage [896]),
    .A1(\shift_storage.storage [895]),
    .S(net245),
    .X(_04874_));
 sg13g2_and2_1 _11561_ (.A(net246),
    .B(_04874_),
    .X(_01586_));
 sg13g2_mux2_1 _11562_ (.A0(\shift_storage.storage [897]),
    .A1(\shift_storage.storage [896]),
    .S(net245),
    .X(_04875_));
 sg13g2_and2_1 _11563_ (.A(net246),
    .B(_04875_),
    .X(_01587_));
 sg13g2_mux2_1 _11564_ (.A0(\shift_storage.storage [898]),
    .A1(\shift_storage.storage [897]),
    .S(net245),
    .X(_04876_));
 sg13g2_and2_1 _11565_ (.A(net246),
    .B(_04876_),
    .X(_01588_));
 sg13g2_buf_1 _11566_ (.A(net399),
    .X(_04877_));
 sg13g2_mux2_1 _11567_ (.A0(\shift_storage.storage [899]),
    .A1(\shift_storage.storage [898]),
    .S(net245),
    .X(_04878_));
 sg13g2_and2_1 _11568_ (.A(net244),
    .B(_04878_),
    .X(_01589_));
 sg13g2_mux2_1 _11569_ (.A0(\shift_storage.storage [89]),
    .A1(\shift_storage.storage [88]),
    .S(net245),
    .X(_04879_));
 sg13g2_and2_1 _11570_ (.A(net244),
    .B(_04879_),
    .X(_01590_));
 sg13g2_mux2_1 _11571_ (.A0(\shift_storage.storage [8]),
    .A1(\shift_storage.storage [7]),
    .S(_04870_),
    .X(_04880_));
 sg13g2_and2_1 _11572_ (.A(net244),
    .B(_04880_),
    .X(_01591_));
 sg13g2_mux2_1 _11573_ (.A0(\shift_storage.storage [900]),
    .A1(\shift_storage.storage [899]),
    .S(_04870_),
    .X(_04881_));
 sg13g2_and2_1 _11574_ (.A(_04877_),
    .B(_04881_),
    .X(_01592_));
 sg13g2_buf_1 _11575_ (.A(_03058_),
    .X(_04882_));
 sg13g2_buf_1 _11576_ (.A(net398),
    .X(_04883_));
 sg13g2_mux2_1 _11577_ (.A0(\shift_storage.storage [901]),
    .A1(\shift_storage.storage [900]),
    .S(net243),
    .X(_04884_));
 sg13g2_and2_1 _11578_ (.A(net244),
    .B(_04884_),
    .X(_01593_));
 sg13g2_mux2_1 _11579_ (.A0(\shift_storage.storage [902]),
    .A1(\shift_storage.storage [901]),
    .S(net243),
    .X(_04885_));
 sg13g2_and2_1 _11580_ (.A(net244),
    .B(_04885_),
    .X(_01594_));
 sg13g2_mux2_1 _11581_ (.A0(\shift_storage.storage [903]),
    .A1(\shift_storage.storage [902]),
    .S(net243),
    .X(_04886_));
 sg13g2_and2_1 _11582_ (.A(net244),
    .B(_04886_),
    .X(_01595_));
 sg13g2_mux2_1 _11583_ (.A0(\shift_storage.storage [904]),
    .A1(\shift_storage.storage [903]),
    .S(net243),
    .X(_04887_));
 sg13g2_and2_1 _11584_ (.A(net244),
    .B(_04887_),
    .X(_01596_));
 sg13g2_mux2_1 _11585_ (.A0(\shift_storage.storage [905]),
    .A1(\shift_storage.storage [904]),
    .S(net243),
    .X(_04888_));
 sg13g2_and2_1 _11586_ (.A(net244),
    .B(_04888_),
    .X(_01597_));
 sg13g2_mux2_1 _11587_ (.A0(\shift_storage.storage [906]),
    .A1(\shift_storage.storage [905]),
    .S(net243),
    .X(_04889_));
 sg13g2_and2_1 _11588_ (.A(_04877_),
    .B(_04889_),
    .X(_01598_));
 sg13g2_buf_1 _11589_ (.A(net494),
    .X(_04890_));
 sg13g2_buf_1 _11590_ (.A(net397),
    .X(_04891_));
 sg13g2_mux2_1 _11591_ (.A0(\shift_storage.storage [907]),
    .A1(\shift_storage.storage [906]),
    .S(net243),
    .X(_04892_));
 sg13g2_and2_1 _11592_ (.A(net242),
    .B(_04892_),
    .X(_01599_));
 sg13g2_mux2_1 _11593_ (.A0(\shift_storage.storage [908]),
    .A1(\shift_storage.storage [907]),
    .S(net243),
    .X(_04893_));
 sg13g2_and2_1 _11594_ (.A(net242),
    .B(_04893_),
    .X(_01600_));
 sg13g2_mux2_1 _11595_ (.A0(\shift_storage.storage [909]),
    .A1(\shift_storage.storage [908]),
    .S(_04883_),
    .X(_04894_));
 sg13g2_and2_1 _11596_ (.A(net242),
    .B(_04894_),
    .X(_01601_));
 sg13g2_mux2_1 _11597_ (.A0(\shift_storage.storage [90]),
    .A1(\shift_storage.storage [89]),
    .S(_04883_),
    .X(_04895_));
 sg13g2_and2_1 _11598_ (.A(net242),
    .B(_04895_),
    .X(_01602_));
 sg13g2_buf_1 _11599_ (.A(net398),
    .X(_04896_));
 sg13g2_mux2_1 _11600_ (.A0(\shift_storage.storage [910]),
    .A1(\shift_storage.storage [909]),
    .S(net241),
    .X(_04897_));
 sg13g2_and2_1 _11601_ (.A(net242),
    .B(_04897_),
    .X(_01603_));
 sg13g2_mux2_1 _11602_ (.A0(\shift_storage.storage [911]),
    .A1(\shift_storage.storage [910]),
    .S(net241),
    .X(_04898_));
 sg13g2_and2_1 _11603_ (.A(net242),
    .B(_04898_),
    .X(_01604_));
 sg13g2_mux2_1 _11604_ (.A0(\shift_storage.storage [912]),
    .A1(\shift_storage.storage [911]),
    .S(net241),
    .X(_04899_));
 sg13g2_and2_1 _11605_ (.A(net242),
    .B(_04899_),
    .X(_01605_));
 sg13g2_mux2_1 _11606_ (.A0(\shift_storage.storage [913]),
    .A1(\shift_storage.storage [912]),
    .S(net241),
    .X(_04900_));
 sg13g2_and2_1 _11607_ (.A(net242),
    .B(_04900_),
    .X(_01606_));
 sg13g2_mux2_1 _11608_ (.A0(\shift_storage.storage [914]),
    .A1(\shift_storage.storage [913]),
    .S(_04896_),
    .X(_04901_));
 sg13g2_and2_1 _11609_ (.A(_04891_),
    .B(_04901_),
    .X(_01607_));
 sg13g2_mux2_1 _11610_ (.A0(\shift_storage.storage [915]),
    .A1(\shift_storage.storage [914]),
    .S(_04896_),
    .X(_04902_));
 sg13g2_and2_1 _11611_ (.A(_04891_),
    .B(_04902_),
    .X(_01608_));
 sg13g2_buf_1 _11612_ (.A(net397),
    .X(_04903_));
 sg13g2_mux2_1 _11613_ (.A0(\shift_storage.storage [916]),
    .A1(\shift_storage.storage [915]),
    .S(net241),
    .X(_04904_));
 sg13g2_and2_1 _11614_ (.A(net240),
    .B(_04904_),
    .X(_01609_));
 sg13g2_mux2_1 _11615_ (.A0(\shift_storage.storage [917]),
    .A1(\shift_storage.storage [916]),
    .S(net241),
    .X(_04905_));
 sg13g2_and2_1 _11616_ (.A(net240),
    .B(_04905_),
    .X(_01610_));
 sg13g2_mux2_1 _11617_ (.A0(\shift_storage.storage [918]),
    .A1(\shift_storage.storage [917]),
    .S(net241),
    .X(_04906_));
 sg13g2_and2_1 _11618_ (.A(net240),
    .B(_04906_),
    .X(_01611_));
 sg13g2_mux2_1 _11619_ (.A0(\shift_storage.storage [919]),
    .A1(\shift_storage.storage [918]),
    .S(net241),
    .X(_04907_));
 sg13g2_and2_1 _11620_ (.A(_04903_),
    .B(_04907_),
    .X(_01612_));
 sg13g2_buf_1 _11621_ (.A(net398),
    .X(_04908_));
 sg13g2_mux2_1 _11622_ (.A0(\shift_storage.storage [91]),
    .A1(\shift_storage.storage [90]),
    .S(net239),
    .X(_04909_));
 sg13g2_and2_1 _11623_ (.A(_04903_),
    .B(_04909_),
    .X(_01613_));
 sg13g2_mux2_1 _11624_ (.A0(\shift_storage.storage [920]),
    .A1(\shift_storage.storage [919]),
    .S(net239),
    .X(_04910_));
 sg13g2_and2_1 _11625_ (.A(net240),
    .B(_04910_),
    .X(_01614_));
 sg13g2_mux2_1 _11626_ (.A0(\shift_storage.storage [921]),
    .A1(\shift_storage.storage [920]),
    .S(net239),
    .X(_04911_));
 sg13g2_and2_1 _11627_ (.A(net240),
    .B(_04911_),
    .X(_01615_));
 sg13g2_mux2_1 _11628_ (.A0(\shift_storage.storage [922]),
    .A1(\shift_storage.storage [921]),
    .S(net239),
    .X(_04912_));
 sg13g2_and2_1 _11629_ (.A(net240),
    .B(_04912_),
    .X(_01616_));
 sg13g2_mux2_1 _11630_ (.A0(\shift_storage.storage [923]),
    .A1(\shift_storage.storage [922]),
    .S(_04908_),
    .X(_04913_));
 sg13g2_and2_1 _11631_ (.A(net240),
    .B(_04913_),
    .X(_01617_));
 sg13g2_mux2_1 _11632_ (.A0(\shift_storage.storage [924]),
    .A1(\shift_storage.storage [923]),
    .S(_04908_),
    .X(_04914_));
 sg13g2_and2_1 _11633_ (.A(net240),
    .B(_04914_),
    .X(_01618_));
 sg13g2_buf_1 _11634_ (.A(net397),
    .X(_04915_));
 sg13g2_mux2_1 _11635_ (.A0(\shift_storage.storage [925]),
    .A1(\shift_storage.storage [924]),
    .S(net239),
    .X(_04916_));
 sg13g2_and2_1 _11636_ (.A(net238),
    .B(_04916_),
    .X(_01619_));
 sg13g2_mux2_1 _11637_ (.A0(\shift_storage.storage [926]),
    .A1(\shift_storage.storage [925]),
    .S(net239),
    .X(_04917_));
 sg13g2_and2_1 _11638_ (.A(net238),
    .B(_04917_),
    .X(_01620_));
 sg13g2_mux2_1 _11639_ (.A0(\shift_storage.storage [927]),
    .A1(\shift_storage.storage [926]),
    .S(net239),
    .X(_04918_));
 sg13g2_and2_1 _11640_ (.A(net238),
    .B(_04918_),
    .X(_01621_));
 sg13g2_mux2_1 _11641_ (.A0(\shift_storage.storage [928]),
    .A1(\shift_storage.storage [927]),
    .S(net239),
    .X(_04919_));
 sg13g2_and2_1 _11642_ (.A(net238),
    .B(_04919_),
    .X(_01622_));
 sg13g2_buf_1 _11643_ (.A(net398),
    .X(_04920_));
 sg13g2_mux2_1 _11644_ (.A0(\shift_storage.storage [929]),
    .A1(\shift_storage.storage [928]),
    .S(net237),
    .X(_04921_));
 sg13g2_and2_1 _11645_ (.A(net238),
    .B(_04921_),
    .X(_01623_));
 sg13g2_mux2_1 _11646_ (.A0(\shift_storage.storage [92]),
    .A1(\shift_storage.storage [91]),
    .S(net237),
    .X(_04922_));
 sg13g2_and2_1 _11647_ (.A(net238),
    .B(_04922_),
    .X(_01624_));
 sg13g2_mux2_1 _11648_ (.A0(\shift_storage.storage [930]),
    .A1(\shift_storage.storage [929]),
    .S(net237),
    .X(_04923_));
 sg13g2_and2_1 _11649_ (.A(net238),
    .B(_04923_),
    .X(_01625_));
 sg13g2_mux2_1 _11650_ (.A0(\shift_storage.storage [931]),
    .A1(\shift_storage.storage [930]),
    .S(net237),
    .X(_04924_));
 sg13g2_and2_1 _11651_ (.A(net238),
    .B(_04924_),
    .X(_01626_));
 sg13g2_mux2_1 _11652_ (.A0(\shift_storage.storage [932]),
    .A1(\shift_storage.storage [931]),
    .S(net237),
    .X(_04925_));
 sg13g2_and2_1 _11653_ (.A(_04915_),
    .B(_04925_),
    .X(_01627_));
 sg13g2_mux2_1 _11654_ (.A0(\shift_storage.storage [933]),
    .A1(\shift_storage.storage [932]),
    .S(net237),
    .X(_04926_));
 sg13g2_and2_1 _11655_ (.A(_04915_),
    .B(_04926_),
    .X(_01628_));
 sg13g2_buf_1 _11656_ (.A(net397),
    .X(_04927_));
 sg13g2_mux2_1 _11657_ (.A0(\shift_storage.storage [934]),
    .A1(\shift_storage.storage [933]),
    .S(net237),
    .X(_04928_));
 sg13g2_and2_1 _11658_ (.A(net236),
    .B(_04928_),
    .X(_01629_));
 sg13g2_mux2_1 _11659_ (.A0(\shift_storage.storage [935]),
    .A1(\shift_storage.storage [934]),
    .S(net237),
    .X(_04929_));
 sg13g2_and2_1 _11660_ (.A(net236),
    .B(_04929_),
    .X(_01630_));
 sg13g2_mux2_1 _11661_ (.A0(\shift_storage.storage [936]),
    .A1(\shift_storage.storage [935]),
    .S(_04920_),
    .X(_04930_));
 sg13g2_and2_1 _11662_ (.A(net236),
    .B(_04930_),
    .X(_01631_));
 sg13g2_mux2_1 _11663_ (.A0(\shift_storage.storage [937]),
    .A1(\shift_storage.storage [936]),
    .S(_04920_),
    .X(_04931_));
 sg13g2_and2_1 _11664_ (.A(net236),
    .B(_04931_),
    .X(_01632_));
 sg13g2_buf_1 _11665_ (.A(net398),
    .X(_04932_));
 sg13g2_mux2_1 _11666_ (.A0(\shift_storage.storage [938]),
    .A1(\shift_storage.storage [937]),
    .S(net235),
    .X(_04933_));
 sg13g2_and2_1 _11667_ (.A(net236),
    .B(_04933_),
    .X(_01633_));
 sg13g2_mux2_1 _11668_ (.A0(\shift_storage.storage [939]),
    .A1(\shift_storage.storage [938]),
    .S(net235),
    .X(_04934_));
 sg13g2_and2_1 _11669_ (.A(net236),
    .B(_04934_),
    .X(_01634_));
 sg13g2_mux2_1 _11670_ (.A0(\shift_storage.storage [93]),
    .A1(\shift_storage.storage [92]),
    .S(_04932_),
    .X(_04935_));
 sg13g2_and2_1 _11671_ (.A(net236),
    .B(_04935_),
    .X(_01635_));
 sg13g2_mux2_1 _11672_ (.A0(\shift_storage.storage [940]),
    .A1(\shift_storage.storage [939]),
    .S(net235),
    .X(_04936_));
 sg13g2_and2_1 _11673_ (.A(net236),
    .B(_04936_),
    .X(_01636_));
 sg13g2_mux2_1 _11674_ (.A0(\shift_storage.storage [941]),
    .A1(\shift_storage.storage [940]),
    .S(net235),
    .X(_04937_));
 sg13g2_and2_1 _11675_ (.A(_04927_),
    .B(_04937_),
    .X(_01637_));
 sg13g2_mux2_1 _11676_ (.A0(\shift_storage.storage [942]),
    .A1(\shift_storage.storage [941]),
    .S(net235),
    .X(_04938_));
 sg13g2_and2_1 _11677_ (.A(_04927_),
    .B(_04938_),
    .X(_01638_));
 sg13g2_buf_1 _11678_ (.A(net397),
    .X(_04939_));
 sg13g2_mux2_1 _11679_ (.A0(\shift_storage.storage [943]),
    .A1(\shift_storage.storage [942]),
    .S(net235),
    .X(_04940_));
 sg13g2_and2_1 _11680_ (.A(net234),
    .B(_04940_),
    .X(_01639_));
 sg13g2_mux2_1 _11681_ (.A0(\shift_storage.storage [944]),
    .A1(\shift_storage.storage [943]),
    .S(net235),
    .X(_04941_));
 sg13g2_and2_1 _11682_ (.A(net234),
    .B(_04941_),
    .X(_01640_));
 sg13g2_mux2_1 _11683_ (.A0(\shift_storage.storage [945]),
    .A1(\shift_storage.storage [944]),
    .S(net235),
    .X(_04942_));
 sg13g2_and2_1 _11684_ (.A(net234),
    .B(_04942_),
    .X(_01641_));
 sg13g2_mux2_1 _11685_ (.A0(\shift_storage.storage [946]),
    .A1(\shift_storage.storage [945]),
    .S(_04932_),
    .X(_04943_));
 sg13g2_and2_1 _11686_ (.A(net234),
    .B(_04943_),
    .X(_01642_));
 sg13g2_buf_1 _11687_ (.A(net398),
    .X(_04944_));
 sg13g2_mux2_1 _11688_ (.A0(\shift_storage.storage [947]),
    .A1(\shift_storage.storage [946]),
    .S(net233),
    .X(_04945_));
 sg13g2_and2_1 _11689_ (.A(net234),
    .B(_04945_),
    .X(_01643_));
 sg13g2_mux2_1 _11690_ (.A0(\shift_storage.storage [948]),
    .A1(\shift_storage.storage [947]),
    .S(net233),
    .X(_04946_));
 sg13g2_and2_1 _11691_ (.A(_04939_),
    .B(_04946_),
    .X(_01644_));
 sg13g2_mux2_1 _11692_ (.A0(\shift_storage.storage [949]),
    .A1(\shift_storage.storage [948]),
    .S(net233),
    .X(_04947_));
 sg13g2_and2_1 _11693_ (.A(net234),
    .B(_04947_),
    .X(_01645_));
 sg13g2_mux2_1 _11694_ (.A0(\shift_storage.storage [94]),
    .A1(\shift_storage.storage [93]),
    .S(net233),
    .X(_04948_));
 sg13g2_and2_1 _11695_ (.A(_04939_),
    .B(_04948_),
    .X(_01646_));
 sg13g2_mux2_1 _11696_ (.A0(\shift_storage.storage [950]),
    .A1(\shift_storage.storage [949]),
    .S(net233),
    .X(_04949_));
 sg13g2_and2_1 _11697_ (.A(net234),
    .B(_04949_),
    .X(_01647_));
 sg13g2_mux2_1 _11698_ (.A0(\shift_storage.storage [951]),
    .A1(\shift_storage.storage [950]),
    .S(net233),
    .X(_04950_));
 sg13g2_and2_1 _11699_ (.A(net234),
    .B(_04950_),
    .X(_01648_));
 sg13g2_buf_1 _11700_ (.A(net397),
    .X(_04951_));
 sg13g2_mux2_1 _11701_ (.A0(\shift_storage.storage [952]),
    .A1(\shift_storage.storage [951]),
    .S(net233),
    .X(_04952_));
 sg13g2_and2_1 _11702_ (.A(net232),
    .B(_04952_),
    .X(_01649_));
 sg13g2_mux2_1 _11703_ (.A0(\shift_storage.storage [953]),
    .A1(\shift_storage.storage [952]),
    .S(net233),
    .X(_04953_));
 sg13g2_and2_1 _11704_ (.A(net232),
    .B(_04953_),
    .X(_01650_));
 sg13g2_mux2_1 _11705_ (.A0(\shift_storage.storage [954]),
    .A1(\shift_storage.storage [953]),
    .S(_04944_),
    .X(_04954_));
 sg13g2_and2_1 _11706_ (.A(net232),
    .B(_04954_),
    .X(_01651_));
 sg13g2_mux2_1 _11707_ (.A0(\shift_storage.storage [955]),
    .A1(\shift_storage.storage [954]),
    .S(_04944_),
    .X(_04955_));
 sg13g2_and2_1 _11708_ (.A(net232),
    .B(_04955_),
    .X(_01652_));
 sg13g2_buf_1 _11709_ (.A(net398),
    .X(_04956_));
 sg13g2_mux2_1 _11710_ (.A0(\shift_storage.storage [956]),
    .A1(\shift_storage.storage [955]),
    .S(net231),
    .X(_04957_));
 sg13g2_and2_1 _11711_ (.A(net232),
    .B(_04957_),
    .X(_01653_));
 sg13g2_mux2_1 _11712_ (.A0(\shift_storage.storage [957]),
    .A1(\shift_storage.storage [956]),
    .S(net231),
    .X(_04958_));
 sg13g2_and2_1 _11713_ (.A(net232),
    .B(_04958_),
    .X(_01654_));
 sg13g2_mux2_1 _11714_ (.A0(\shift_storage.storage [958]),
    .A1(\shift_storage.storage [957]),
    .S(net231),
    .X(_04959_));
 sg13g2_and2_1 _11715_ (.A(net232),
    .B(_04959_),
    .X(_01655_));
 sg13g2_mux2_1 _11716_ (.A0(\shift_storage.storage [959]),
    .A1(\shift_storage.storage [958]),
    .S(net231),
    .X(_04960_));
 sg13g2_and2_1 _11717_ (.A(_04951_),
    .B(_04960_),
    .X(_01656_));
 sg13g2_mux2_1 _11718_ (.A0(\shift_storage.storage [95]),
    .A1(\shift_storage.storage [94]),
    .S(net231),
    .X(_04961_));
 sg13g2_and2_1 _11719_ (.A(net232),
    .B(_04961_),
    .X(_01657_));
 sg13g2_mux2_1 _11720_ (.A0(\shift_storage.storage [960]),
    .A1(\shift_storage.storage [959]),
    .S(net231),
    .X(_04962_));
 sg13g2_and2_1 _11721_ (.A(_04951_),
    .B(_04962_),
    .X(_01658_));
 sg13g2_buf_1 _11722_ (.A(net397),
    .X(_04963_));
 sg13g2_mux2_1 _11723_ (.A0(\shift_storage.storage [961]),
    .A1(\shift_storage.storage [960]),
    .S(net231),
    .X(_04964_));
 sg13g2_and2_1 _11724_ (.A(net230),
    .B(_04964_),
    .X(_01659_));
 sg13g2_mux2_1 _11725_ (.A0(\shift_storage.storage [962]),
    .A1(\shift_storage.storage [961]),
    .S(net231),
    .X(_04965_));
 sg13g2_and2_1 _11726_ (.A(net230),
    .B(_04965_),
    .X(_01660_));
 sg13g2_mux2_1 _11727_ (.A0(\shift_storage.storage [963]),
    .A1(\shift_storage.storage [962]),
    .S(_04956_),
    .X(_04966_));
 sg13g2_and2_1 _11728_ (.A(net230),
    .B(_04966_),
    .X(_01661_));
 sg13g2_mux2_1 _11729_ (.A0(\shift_storage.storage [964]),
    .A1(\shift_storage.storage [963]),
    .S(_04956_),
    .X(_04967_));
 sg13g2_and2_1 _11730_ (.A(_04963_),
    .B(_04967_),
    .X(_01662_));
 sg13g2_buf_1 _11731_ (.A(net398),
    .X(_04968_));
 sg13g2_mux2_1 _11732_ (.A0(\shift_storage.storage [965]),
    .A1(\shift_storage.storage [964]),
    .S(net229),
    .X(_04969_));
 sg13g2_and2_1 _11733_ (.A(_04963_),
    .B(_04969_),
    .X(_01663_));
 sg13g2_mux2_1 _11734_ (.A0(\shift_storage.storage [966]),
    .A1(\shift_storage.storage [965]),
    .S(net229),
    .X(_04970_));
 sg13g2_and2_1 _11735_ (.A(net230),
    .B(_04970_),
    .X(_01664_));
 sg13g2_mux2_1 _11736_ (.A0(\shift_storage.storage [967]),
    .A1(\shift_storage.storage [966]),
    .S(_04968_),
    .X(_04971_));
 sg13g2_and2_1 _11737_ (.A(net230),
    .B(_04971_),
    .X(_01665_));
 sg13g2_mux2_1 _11738_ (.A0(\shift_storage.storage [968]),
    .A1(\shift_storage.storage [967]),
    .S(_04968_),
    .X(_04972_));
 sg13g2_and2_1 _11739_ (.A(net230),
    .B(_04972_),
    .X(_01666_));
 sg13g2_mux2_1 _11740_ (.A0(\shift_storage.storage [969]),
    .A1(\shift_storage.storage [968]),
    .S(net229),
    .X(_04973_));
 sg13g2_and2_1 _11741_ (.A(net230),
    .B(_04973_),
    .X(_01667_));
 sg13g2_mux2_1 _11742_ (.A0(\shift_storage.storage [96]),
    .A1(\shift_storage.storage [95]),
    .S(net229),
    .X(_04974_));
 sg13g2_and2_1 _11743_ (.A(net230),
    .B(_04974_),
    .X(_01668_));
 sg13g2_buf_1 _11744_ (.A(net397),
    .X(_04975_));
 sg13g2_mux2_1 _11745_ (.A0(\shift_storage.storage [970]),
    .A1(\shift_storage.storage [969]),
    .S(net229),
    .X(_04976_));
 sg13g2_and2_1 _11746_ (.A(net228),
    .B(_04976_),
    .X(_01669_));
 sg13g2_mux2_1 _11747_ (.A0(\shift_storage.storage [971]),
    .A1(\shift_storage.storage [970]),
    .S(net229),
    .X(_04977_));
 sg13g2_and2_1 _11748_ (.A(net228),
    .B(_04977_),
    .X(_01670_));
 sg13g2_mux2_1 _11749_ (.A0(\shift_storage.storage [972]),
    .A1(\shift_storage.storage [971]),
    .S(net229),
    .X(_04978_));
 sg13g2_and2_1 _11750_ (.A(net228),
    .B(_04978_),
    .X(_01671_));
 sg13g2_mux2_1 _11751_ (.A0(\shift_storage.storage [973]),
    .A1(\shift_storage.storage [972]),
    .S(net229),
    .X(_04979_));
 sg13g2_and2_1 _11752_ (.A(_04975_),
    .B(_04979_),
    .X(_01672_));
 sg13g2_buf_1 _11753_ (.A(_04882_),
    .X(_04980_));
 sg13g2_mux2_1 _11754_ (.A0(\shift_storage.storage [974]),
    .A1(\shift_storage.storage [973]),
    .S(net227),
    .X(_04981_));
 sg13g2_and2_1 _11755_ (.A(_04975_),
    .B(_04981_),
    .X(_01673_));
 sg13g2_mux2_1 _11756_ (.A0(\shift_storage.storage [975]),
    .A1(\shift_storage.storage [974]),
    .S(net227),
    .X(_04982_));
 sg13g2_and2_1 _11757_ (.A(net228),
    .B(_04982_),
    .X(_01674_));
 sg13g2_mux2_1 _11758_ (.A0(\shift_storage.storage [976]),
    .A1(\shift_storage.storage [975]),
    .S(net227),
    .X(_04983_));
 sg13g2_and2_1 _11759_ (.A(net228),
    .B(_04983_),
    .X(_01675_));
 sg13g2_mux2_1 _11760_ (.A0(\shift_storage.storage [977]),
    .A1(\shift_storage.storage [976]),
    .S(net227),
    .X(_04984_));
 sg13g2_and2_1 _11761_ (.A(net228),
    .B(_04984_),
    .X(_01676_));
 sg13g2_mux2_1 _11762_ (.A0(\shift_storage.storage [978]),
    .A1(\shift_storage.storage [977]),
    .S(net227),
    .X(_04985_));
 sg13g2_and2_1 _11763_ (.A(net228),
    .B(_04985_),
    .X(_01677_));
 sg13g2_mux2_1 _11764_ (.A0(\shift_storage.storage [979]),
    .A1(\shift_storage.storage [978]),
    .S(net227),
    .X(_04986_));
 sg13g2_and2_1 _11765_ (.A(net228),
    .B(_04986_),
    .X(_01678_));
 sg13g2_buf_1 _11766_ (.A(_04890_),
    .X(_04987_));
 sg13g2_mux2_1 _11767_ (.A0(\shift_storage.storage [97]),
    .A1(\shift_storage.storage [96]),
    .S(_04980_),
    .X(_04988_));
 sg13g2_and2_1 _11768_ (.A(net226),
    .B(_04988_),
    .X(_01679_));
 sg13g2_mux2_1 _11769_ (.A0(\shift_storage.storage [980]),
    .A1(\shift_storage.storage [979]),
    .S(net227),
    .X(_04989_));
 sg13g2_and2_1 _11770_ (.A(net226),
    .B(_04989_),
    .X(_01680_));
 sg13g2_mux2_1 _11771_ (.A0(\shift_storage.storage [981]),
    .A1(\shift_storage.storage [980]),
    .S(net227),
    .X(_04990_));
 sg13g2_and2_1 _11772_ (.A(net226),
    .B(_04990_),
    .X(_01681_));
 sg13g2_mux2_1 _11773_ (.A0(\shift_storage.storage [982]),
    .A1(\shift_storage.storage [981]),
    .S(_04980_),
    .X(_04991_));
 sg13g2_and2_1 _11774_ (.A(net226),
    .B(_04991_),
    .X(_01682_));
 sg13g2_buf_1 _11775_ (.A(_04882_),
    .X(_04992_));
 sg13g2_mux2_1 _11776_ (.A0(\shift_storage.storage [983]),
    .A1(\shift_storage.storage [982]),
    .S(net225),
    .X(_04993_));
 sg13g2_and2_1 _11777_ (.A(net226),
    .B(_04993_),
    .X(_01683_));
 sg13g2_mux2_1 _11778_ (.A0(\shift_storage.storage [984]),
    .A1(\shift_storage.storage [983]),
    .S(net225),
    .X(_04994_));
 sg13g2_and2_1 _11779_ (.A(net226),
    .B(_04994_),
    .X(_01684_));
 sg13g2_mux2_1 _11780_ (.A0(\shift_storage.storage [985]),
    .A1(\shift_storage.storage [984]),
    .S(net225),
    .X(_04995_));
 sg13g2_and2_1 _11781_ (.A(net226),
    .B(_04995_),
    .X(_01685_));
 sg13g2_mux2_1 _11782_ (.A0(\shift_storage.storage [986]),
    .A1(\shift_storage.storage [985]),
    .S(net225),
    .X(_04996_));
 sg13g2_and2_1 _11783_ (.A(net226),
    .B(_04996_),
    .X(_01686_));
 sg13g2_mux2_1 _11784_ (.A0(\shift_storage.storage [987]),
    .A1(\shift_storage.storage [986]),
    .S(net225),
    .X(_04997_));
 sg13g2_and2_1 _11785_ (.A(_04987_),
    .B(_04997_),
    .X(_01687_));
 sg13g2_mux2_1 _11786_ (.A0(\shift_storage.storage [988]),
    .A1(\shift_storage.storage [987]),
    .S(net225),
    .X(_04998_));
 sg13g2_and2_1 _11787_ (.A(_04987_),
    .B(_04998_),
    .X(_01688_));
 sg13g2_buf_1 _11788_ (.A(_04890_),
    .X(_04999_));
 sg13g2_mux2_1 _11789_ (.A0(\shift_storage.storage [989]),
    .A1(\shift_storage.storage [988]),
    .S(net225),
    .X(_05000_));
 sg13g2_and2_1 _11790_ (.A(net224),
    .B(_05000_),
    .X(_01689_));
 sg13g2_mux2_1 _11791_ (.A0(\shift_storage.storage [98]),
    .A1(\shift_storage.storage [97]),
    .S(net225),
    .X(_05001_));
 sg13g2_and2_1 _11792_ (.A(net224),
    .B(_05001_),
    .X(_01690_));
 sg13g2_mux2_1 _11793_ (.A0(\shift_storage.storage [990]),
    .A1(\shift_storage.storage [989]),
    .S(_04992_),
    .X(_05002_));
 sg13g2_and2_1 _11794_ (.A(net224),
    .B(_05002_),
    .X(_01691_));
 sg13g2_mux2_1 _11795_ (.A0(\shift_storage.storage [991]),
    .A1(\shift_storage.storage [990]),
    .S(_04992_),
    .X(_05003_));
 sg13g2_and2_1 _11796_ (.A(net224),
    .B(_05003_),
    .X(_01692_));
 sg13g2_buf_1 _11797_ (.A(net410),
    .X(_05004_));
 sg13g2_mux2_1 _11798_ (.A0(\shift_storage.storage [992]),
    .A1(\shift_storage.storage [991]),
    .S(net223),
    .X(_05005_));
 sg13g2_and2_1 _11799_ (.A(net224),
    .B(_05005_),
    .X(_01693_));
 sg13g2_mux2_1 _11800_ (.A0(\shift_storage.storage [993]),
    .A1(\shift_storage.storage [992]),
    .S(net223),
    .X(_05006_));
 sg13g2_and2_1 _11801_ (.A(net224),
    .B(_05006_),
    .X(_01694_));
 sg13g2_mux2_1 _11802_ (.A0(\shift_storage.storage [994]),
    .A1(\shift_storage.storage [993]),
    .S(net223),
    .X(_05007_));
 sg13g2_and2_1 _11803_ (.A(net224),
    .B(_05007_),
    .X(_01695_));
 sg13g2_mux2_1 _11804_ (.A0(\shift_storage.storage [995]),
    .A1(\shift_storage.storage [994]),
    .S(net223),
    .X(_05008_));
 sg13g2_and2_1 _11805_ (.A(net224),
    .B(_05008_),
    .X(_01696_));
 sg13g2_mux2_1 _11806_ (.A0(\shift_storage.storage [996]),
    .A1(\shift_storage.storage [995]),
    .S(net223),
    .X(_05009_));
 sg13g2_and2_1 _11807_ (.A(_04999_),
    .B(_05009_),
    .X(_01697_));
 sg13g2_mux2_1 _11808_ (.A0(\shift_storage.storage [997]),
    .A1(\shift_storage.storage [996]),
    .S(net223),
    .X(_05010_));
 sg13g2_and2_1 _11809_ (.A(_04999_),
    .B(_05010_),
    .X(_01698_));
 sg13g2_mux2_1 _11810_ (.A0(\shift_storage.storage [998]),
    .A1(\shift_storage.storage [997]),
    .S(net223),
    .X(_05011_));
 sg13g2_and2_1 _11811_ (.A(net412),
    .B(_05011_),
    .X(_01699_));
 sg13g2_mux2_1 _11812_ (.A0(\shift_storage.storage [999]),
    .A1(\shift_storage.storage [998]),
    .S(_05004_),
    .X(_05012_));
 sg13g2_and2_1 _11813_ (.A(net412),
    .B(_05012_),
    .X(_01700_));
 sg13g2_mux2_1 _11814_ (.A0(\shift_storage.storage [99]),
    .A1(\shift_storage.storage [98]),
    .S(net223),
    .X(_05013_));
 sg13g2_and2_1 _11815_ (.A(net412),
    .B(_05013_),
    .X(_01701_));
 sg13g2_mux2_1 _11816_ (.A0(\shift_storage.storage [9]),
    .A1(\shift_storage.storage [8]),
    .S(_05004_),
    .X(_05014_));
 sg13g2_and2_1 _11817_ (.A(net412),
    .B(_05014_),
    .X(_01702_));
 sg13g2_buf_1 _11818_ (.A(out_select_p2c_2),
    .X(_05015_));
 sg13g2_inv_1 _11819_ (.Y(_05016_),
    .A(net487));
 sg13g2_buf_1 _11820_ (.A(out_select_p2c_1),
    .X(_05017_));
 sg13g2_nand3_1 _11821_ (.B(\median_processor.median_processor.median_out [0]),
    .C(net493),
    .A(net486),
    .Y(_05018_));
 sg13g2_o21ai_1 _11822_ (.B1(_05018_),
    .Y(_05019_),
    .A1(net486),
    .A2(\median_processor.median_processor.median_out [0]));
 sg13g2_buf_1 _11823_ (.A(out_select_p2c_1),
    .X(_05020_));
 sg13g2_nand2_1 _11824_ (.Y(_05021_),
    .A(net485),
    .B(\median_processor.median_processor.median_out [0]));
 sg13g2_inv_2 _11825_ (.Y(_05022_),
    .A(out_select_p2c_1));
 sg13g2_nand2_1 _11826_ (.Y(_05023_),
    .A(_05022_),
    .B(data_in_p2c_1));
 sg13g2_nand3_1 _11827_ (.B(_05021_),
    .C(_05023_),
    .A(out_select_p2c_2),
    .Y(_05024_));
 sg13g2_o21ai_1 _11828_ (.B1(_05024_),
    .Y(_05025_),
    .A1(\median_processor.median_processor.median_out [0]),
    .A2(net493));
 sg13g2_a21oi_2 _11829_ (.B1(_05025_),
    .Y(data_out_c2p[0]),
    .A2(_05019_),
    .A1(_05016_));
 sg13g2_nor2b_2 _11830_ (.A(data_in_p2c_1),
    .B_N(\median_processor.median_processor.median_out [0]),
    .Y(_05026_));
 sg13g2_o21ai_1 _11831_ (.B1(net486),
    .Y(_05027_),
    .A1(net488),
    .A2(_05026_));
 sg13g2_xor2_1 _11832_ (.B(_05026_),
    .A(data_in_p2c_2),
    .X(_05028_));
 sg13g2_nor2_1 _11833_ (.A(_05022_),
    .B(\median_processor.median_processor.median_out [1]),
    .Y(_05029_));
 sg13g2_a22oi_1 _11834_ (.Y(_05030_),
    .B1(_05028_),
    .B2(_05029_),
    .A2(_05027_),
    .A1(\median_processor.median_processor.median_out [1]));
 sg13g2_and2_1 _11835_ (.A(\median_processor.median_processor.median_out [1]),
    .B(data_in_p2c_2),
    .X(_05031_));
 sg13g2_mux2_1 _11836_ (.A0(net488),
    .A1(\median_processor.median_processor.median_out [1]),
    .S(net485),
    .X(_05032_));
 sg13g2_a22oi_1 _11837_ (.Y(_05033_),
    .B1(_05032_),
    .B2(net487),
    .A2(_05031_),
    .A1(_05026_));
 sg13g2_o21ai_1 _11838_ (.B1(_05033_),
    .Y(net29),
    .A1(net487),
    .A2(_05030_));
 sg13g2_nand2b_1 _11839_ (.Y(_05034_),
    .B(data_in_p2c_2),
    .A_N(\median_processor.median_processor.median_out [1]));
 sg13g2_nor2b_1 _11840_ (.A(data_in_p2c_2),
    .B_N(\median_processor.median_processor.median_out [1]),
    .Y(_05035_));
 sg13g2_a21o_2 _11841_ (.A2(_05034_),
    .A1(_05026_),
    .B1(_05035_),
    .X(_05036_));
 sg13g2_o21ai_1 _11842_ (.B1(net486),
    .Y(_05037_),
    .A1(data_in_p2c_3),
    .A2(_05036_));
 sg13g2_nor2_1 _11843_ (.A(_05022_),
    .B(\median_processor.median_processor.median_out [2]),
    .Y(_05038_));
 sg13g2_xnor2_1 _11844_ (.Y(_05039_),
    .A(_02920_),
    .B(_05036_));
 sg13g2_a22oi_1 _11845_ (.Y(_05040_),
    .B1(_05038_),
    .B2(_05039_),
    .A2(_05037_),
    .A1(\median_processor.median_processor.median_out [2]));
 sg13g2_nand2_1 _11846_ (.Y(_05041_),
    .A(net485),
    .B(\median_processor.median_processor.median_out [2]));
 sg13g2_o21ai_1 _11847_ (.B1(_05041_),
    .Y(_05042_),
    .A1(net485),
    .A2(_02920_));
 sg13g2_and2_1 _11848_ (.A(\median_processor.median_processor.median_out [2]),
    .B(data_in_p2c_3),
    .X(_05043_));
 sg13g2_a22oi_1 _11849_ (.Y(_05044_),
    .B1(_05043_),
    .B2(_05036_),
    .A2(_05042_),
    .A1(out_select_p2c_2));
 sg13g2_o21ai_1 _11850_ (.B1(_05044_),
    .Y(net27),
    .A1(net487),
    .A2(_05040_));
 sg13g2_nor2_1 _11851_ (.A(_02920_),
    .B(_05036_),
    .Y(_05045_));
 sg13g2_a21oi_1 _11852_ (.A1(_02920_),
    .A2(_05036_),
    .Y(_05046_),
    .B1(\median_processor.median_processor.median_out [2]));
 sg13g2_or2_1 _11853_ (.X(_05047_),
    .B(_05046_),
    .A(_05045_));
 sg13g2_nor2_1 _11854_ (.A(\median_processor.median_processor.median_out [3]),
    .B(net492),
    .Y(_05048_));
 sg13g2_and2_1 _11855_ (.A(out_select_p2c_1),
    .B(\median_processor.median_processor.median_out [3]),
    .X(_05049_));
 sg13g2_a21oi_1 _11856_ (.A1(_05022_),
    .A2(net492),
    .Y(_05050_),
    .B1(_05049_));
 sg13g2_xnor2_1 _11857_ (.Y(_05051_),
    .A(data_in_p2c_4),
    .B(_05047_));
 sg13g2_nand2b_1 _11858_ (.Y(_05052_),
    .B(data_in_p2c_4),
    .A_N(_05047_));
 sg13g2_a21oi_1 _11859_ (.A1(net485),
    .A2(_05052_),
    .Y(_05053_),
    .B1(\median_processor.median_processor.median_out [3]));
 sg13g2_a21oi_1 _11860_ (.A1(_05049_),
    .A2(_05051_),
    .Y(_05054_),
    .B1(_05053_));
 sg13g2_nor2_1 _11861_ (.A(out_select_p2c_2),
    .B(_05054_),
    .Y(_05055_));
 sg13g2_a221oi_1 _11862_ (.B2(net487),
    .C1(_05055_),
    .B1(_05050_),
    .A1(_05047_),
    .Y(net13),
    .A2(_05048_));
 sg13g2_o21ai_1 _11863_ (.B1(data_in_p2c_4),
    .Y(_05056_),
    .A1(_05045_),
    .A2(_05046_));
 sg13g2_nor3_1 _11864_ (.A(data_in_p2c_4),
    .B(_05045_),
    .C(_05046_),
    .Y(_05057_));
 sg13g2_a21o_1 _11865_ (.A2(_05056_),
    .A1(\median_processor.median_processor.median_out [3]),
    .B1(_05057_),
    .X(_05058_));
 sg13g2_o21ai_1 _11866_ (.B1(net486),
    .Y(_05059_),
    .A1(net491),
    .A2(_05058_));
 sg13g2_xnor2_1 _11867_ (.Y(_05060_),
    .A(data_in_p2c_5),
    .B(_05058_));
 sg13g2_nor3_1 _11868_ (.A(_05022_),
    .B(\median_processor.median_processor.median_out [4]),
    .C(_05060_),
    .Y(_05061_));
 sg13g2_a21oi_1 _11869_ (.A1(\median_processor.median_processor.median_out [4]),
    .A2(_05059_),
    .Y(_05062_),
    .B1(_05061_));
 sg13g2_mux2_1 _11870_ (.A0(data_in_p2c_5),
    .A1(\median_processor.median_processor.median_out [4]),
    .S(out_select_p2c_1),
    .X(_05063_));
 sg13g2_and2_1 _11871_ (.A(\median_processor.median_processor.median_out [4]),
    .B(net491),
    .X(_05064_));
 sg13g2_a22oi_1 _11872_ (.Y(_05065_),
    .B1(_05064_),
    .B2(_05058_),
    .A2(_05063_),
    .A1(out_select_p2c_2));
 sg13g2_o21ai_1 _11873_ (.B1(_05065_),
    .Y(net12),
    .A1(net487),
    .A2(_05062_));
 sg13g2_nor2b_1 _11874_ (.A(data_in_p2c_5),
    .B_N(_05058_),
    .Y(_05066_));
 sg13g2_nand2b_1 _11875_ (.Y(_05067_),
    .B(data_in_p2c_5),
    .A_N(_05058_));
 sg13g2_o21ai_1 _11876_ (.B1(_05067_),
    .Y(_05068_),
    .A1(\median_processor.median_processor.median_out [4]),
    .A2(_05066_));
 sg13g2_nor2_1 _11877_ (.A(\median_processor.median_processor.median_out [5]),
    .B(net490),
    .Y(_05069_));
 sg13g2_and2_1 _11878_ (.A(net485),
    .B(\median_processor.median_processor.median_out [5]),
    .X(_05070_));
 sg13g2_a21oi_1 _11879_ (.A1(_05022_),
    .A2(net490),
    .Y(_05071_),
    .B1(_05070_));
 sg13g2_nand2b_1 _11880_ (.Y(_05072_),
    .B(data_in_p2c_6),
    .A_N(_05068_));
 sg13g2_a21o_1 _11881_ (.A2(_05072_),
    .A1(net485),
    .B1(\median_processor.median_processor.median_out [5]),
    .X(_05073_));
 sg13g2_nand2b_1 _11882_ (.Y(_05074_),
    .B(_05068_),
    .A_N(data_in_p2c_6));
 sg13g2_nand4_1 _11883_ (.B(\median_processor.median_processor.median_out [5]),
    .C(_05072_),
    .A(net486),
    .Y(_05075_),
    .D(_05074_));
 sg13g2_a21oi_1 _11884_ (.A1(_05073_),
    .A2(_05075_),
    .Y(_05076_),
    .B1(net487));
 sg13g2_a221oi_1 _11885_ (.B2(net487),
    .C1(_05076_),
    .B1(_05071_),
    .A1(_05068_),
    .Y(net11),
    .A2(_05069_));
 sg13g2_nand2_1 _11886_ (.Y(_05077_),
    .A(data_in_p2c_6),
    .B(_05068_));
 sg13g2_nor2_1 _11887_ (.A(data_in_p2c_6),
    .B(_05068_),
    .Y(_05078_));
 sg13g2_a21oi_2 _11888_ (.B1(_05078_),
    .Y(_05079_),
    .A2(_05077_),
    .A1(\median_processor.median_processor.median_out [5]));
 sg13g2_nor2_1 _11889_ (.A(\median_processor.median_processor.median_out [6]),
    .B(net495),
    .Y(_05080_));
 sg13g2_nor2_1 _11890_ (.A(net486),
    .B(_02929_),
    .Y(_05081_));
 sg13g2_a21oi_1 _11891_ (.A1(net486),
    .A2(\median_processor.median_processor.median_out [6]),
    .Y(_05082_),
    .B1(_05081_));
 sg13g2_o21ai_1 _11892_ (.B1(net485),
    .Y(_05083_),
    .A1(_02929_),
    .A2(_05079_));
 sg13g2_nand2b_1 _11893_ (.Y(_05084_),
    .B(_05083_),
    .A_N(\median_processor.median_processor.median_out [6]));
 sg13g2_xnor2_1 _11894_ (.Y(_05085_),
    .A(net495),
    .B(_05079_));
 sg13g2_nand3_1 _11895_ (.B(\median_processor.median_processor.median_out [6]),
    .C(_05085_),
    .A(_05017_),
    .Y(_05086_));
 sg13g2_a21oi_1 _11896_ (.A1(_05084_),
    .A2(_05086_),
    .Y(_05087_),
    .B1(out_select_p2c_2));
 sg13g2_a221oi_1 _11897_ (.B2(_05015_),
    .C1(_05087_),
    .B1(_05082_),
    .A1(_05079_),
    .Y(net8),
    .A2(_05080_));
 sg13g2_nand2_1 _11898_ (.Y(_05088_),
    .A(net495),
    .B(_05079_));
 sg13g2_nor2_1 _11899_ (.A(net495),
    .B(_05079_),
    .Y(_05089_));
 sg13g2_a21oi_1 _11900_ (.A1(\median_processor.median_processor.median_out [6]),
    .A2(_05088_),
    .Y(_05090_),
    .B1(_05089_));
 sg13g2_nor2_1 _11901_ (.A(\median_processor.median_processor.median_out [7]),
    .B(net489),
    .Y(_05091_));
 sg13g2_and2_1 _11902_ (.A(_05020_),
    .B(\median_processor.median_processor.median_out [7]),
    .X(_05092_));
 sg13g2_a21oi_1 _11903_ (.A1(_05022_),
    .A2(net489),
    .Y(_05093_),
    .B1(_05092_));
 sg13g2_nand2b_1 _11904_ (.Y(_05094_),
    .B(data_in_p2c_8),
    .A_N(_05090_));
 sg13g2_a21o_1 _11905_ (.A2(_05094_),
    .A1(_05020_),
    .B1(\median_processor.median_processor.median_out [7]),
    .X(_05095_));
 sg13g2_nand2b_1 _11906_ (.Y(_05096_),
    .B(_05090_),
    .A_N(data_in_p2c_8));
 sg13g2_nand4_1 _11907_ (.B(\median_processor.median_processor.median_out [7]),
    .C(_05094_),
    .A(_05017_),
    .Y(_05097_),
    .D(_05096_));
 sg13g2_a21oi_1 _11908_ (.A1(_05095_),
    .A2(_05097_),
    .Y(_05098_),
    .B1(out_select_p2c_2));
 sg13g2_a221oi_1 _11909_ (.B2(_05015_),
    .C1(_05098_),
    .B1(_05093_),
    .A1(_05090_),
    .Y(net3),
    .A2(_05091_));
 sg13g2_buf_4 clkbuf_leaf_0_clk_p2c (.X(clknet_leaf_0_clk_p2c),
    .A(clknet_5_0__leaf_clk_p2c));
 sg13g2_dfrbp_1 \median_processor.input_storage[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_181_clk_p2c),
    .RESET_B(net496),
    .D(_00000_),
    .Q_N(_06801_),
    .Q(\median_processor.input_storage [0]));
 sg13g2_dfrbp_1 \median_processor.input_storage[10]$_SDFFE_PN0P_  (.CLK(clknet_leaf_179_clk_p2c),
    .RESET_B(net497),
    .D(_00001_),
    .Q_N(_06800_),
    .Q(\median_processor.input_storage [10]));
 sg13g2_dfrbp_1 \median_processor.input_storage[11]$_SDFFE_PN0P_  (.CLK(clknet_leaf_180_clk_p2c),
    .RESET_B(net498),
    .D(_00002_),
    .Q_N(_06799_),
    .Q(\median_processor.input_storage [11]));
 sg13g2_dfrbp_1 \median_processor.input_storage[12]$_SDFFE_PN0P_  (.CLK(clknet_leaf_177_clk_p2c),
    .RESET_B(net499),
    .D(_00003_),
    .Q_N(_06798_),
    .Q(\median_processor.input_storage [12]));
 sg13g2_dfrbp_1 \median_processor.input_storage[13]$_SDFFE_PN0P_  (.CLK(clknet_leaf_176_clk_p2c),
    .RESET_B(net500),
    .D(_00004_),
    .Q_N(_06797_),
    .Q(\median_processor.input_storage [13]));
 sg13g2_dfrbp_1 \median_processor.input_storage[14]$_SDFFE_PN0P_  (.CLK(clknet_leaf_174_clk_p2c),
    .RESET_B(net501),
    .D(_00005_),
    .Q_N(_06796_),
    .Q(\median_processor.input_storage [14]));
 sg13g2_dfrbp_1 \median_processor.input_storage[15]$_SDFFE_PN0P_  (.CLK(clknet_leaf_174_clk_p2c),
    .RESET_B(net502),
    .D(_00006_),
    .Q_N(_06795_),
    .Q(\median_processor.input_storage [15]));
 sg13g2_dfrbp_1 \median_processor.input_storage[16]$_SDFFE_PN0P_  (.CLK(clknet_leaf_160_clk_p2c),
    .RESET_B(net503),
    .D(_00007_),
    .Q_N(_06794_),
    .Q(\median_processor.input_storage [16]));
 sg13g2_dfrbp_1 \median_processor.input_storage[17]$_SDFFE_PN0P_  (.CLK(clknet_leaf_160_clk_p2c),
    .RESET_B(net504),
    .D(_00008_),
    .Q_N(_06793_),
    .Q(\median_processor.input_storage [17]));
 sg13g2_dfrbp_1 \median_processor.input_storage[18]$_SDFFE_PN0P_  (.CLK(clknet_leaf_160_clk_p2c),
    .RESET_B(net505),
    .D(_00009_),
    .Q_N(_06792_),
    .Q(\median_processor.input_storage [18]));
 sg13g2_dfrbp_1 \median_processor.input_storage[19]$_SDFFE_PN0P_  (.CLK(clknet_leaf_182_clk_p2c),
    .RESET_B(net506),
    .D(_00010_),
    .Q_N(_06791_),
    .Q(\median_processor.input_storage [19]));
 sg13g2_dfrbp_1 \median_processor.input_storage[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_182_clk_p2c),
    .RESET_B(net507),
    .D(_00011_),
    .Q_N(_06790_),
    .Q(\median_processor.input_storage [1]));
 sg13g2_dfrbp_1 \median_processor.input_storage[20]$_SDFFE_PN0P_  (.CLK(clknet_leaf_171_clk_p2c),
    .RESET_B(net508),
    .D(_00012_),
    .Q_N(_06789_),
    .Q(\median_processor.input_storage [20]));
 sg13g2_dfrbp_1 \median_processor.input_storage[21]$_SDFFE_PN0P_  (.CLK(clknet_leaf_168_clk_p2c),
    .RESET_B(net509),
    .D(_00013_),
    .Q_N(_06788_),
    .Q(\median_processor.input_storage [21]));
 sg13g2_dfrbp_1 \median_processor.input_storage[22]$_SDFFE_PN0P_  (.CLK(clknet_leaf_168_clk_p2c),
    .RESET_B(net510),
    .D(_00014_),
    .Q_N(_06787_),
    .Q(\median_processor.input_storage [22]));
 sg13g2_dfrbp_1 \median_processor.input_storage[23]$_SDFFE_PN0P_  (.CLK(clknet_leaf_168_clk_p2c),
    .RESET_B(net511),
    .D(_00015_),
    .Q_N(_06786_),
    .Q(\median_processor.input_storage [23]));
 sg13g2_dfrbp_1 \median_processor.input_storage[24]$_SDFFE_PN0P_  (.CLK(clknet_leaf_160_clk_p2c),
    .RESET_B(net512),
    .D(_00016_),
    .Q_N(_06785_),
    .Q(\median_processor.input_storage [24]));
 sg13g2_dfrbp_1 \median_processor.input_storage[25]$_SDFFE_PN0P_  (.CLK(clknet_leaf_160_clk_p2c),
    .RESET_B(net513),
    .D(_00017_),
    .Q_N(_06784_),
    .Q(\median_processor.input_storage [25]));
 sg13g2_dfrbp_1 \median_processor.input_storage[26]$_SDFFE_PN0P_  (.CLK(clknet_leaf_161_clk_p2c),
    .RESET_B(net514),
    .D(_00018_),
    .Q_N(_06783_),
    .Q(\median_processor.input_storage [26]));
 sg13g2_dfrbp_1 \median_processor.input_storage[27]$_SDFFE_PN0P_  (.CLK(clknet_leaf_162_clk_p2c),
    .RESET_B(net515),
    .D(_00019_),
    .Q_N(_06782_),
    .Q(\median_processor.input_storage [27]));
 sg13g2_dfrbp_1 \median_processor.input_storage[28]$_SDFFE_PN0P_  (.CLK(clknet_leaf_172_clk_p2c),
    .RESET_B(net516),
    .D(_00020_),
    .Q_N(_06781_),
    .Q(\median_processor.input_storage [28]));
 sg13g2_dfrbp_1 \median_processor.input_storage[29]$_SDFFE_PN0P_  (.CLK(clknet_leaf_169_clk_p2c),
    .RESET_B(net517),
    .D(_00021_),
    .Q_N(_06780_),
    .Q(\median_processor.input_storage [29]));
 sg13g2_dfrbp_1 \median_processor.input_storage[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_181_clk_p2c),
    .RESET_B(net518),
    .D(_00022_),
    .Q_N(_06779_),
    .Q(\median_processor.input_storage [2]));
 sg13g2_dfrbp_1 \median_processor.input_storage[30]$_SDFFE_PN0P_  (.CLK(clknet_leaf_169_clk_p2c),
    .RESET_B(net519),
    .D(_00023_),
    .Q_N(_06778_),
    .Q(\median_processor.input_storage [30]));
 sg13g2_dfrbp_1 \median_processor.input_storage[31]$_SDFFE_PN0P_  (.CLK(clknet_leaf_168_clk_p2c),
    .RESET_B(net520),
    .D(_00024_),
    .Q_N(_06777_),
    .Q(\median_processor.input_storage [31]));
 sg13g2_dfrbp_1 \median_processor.input_storage[32]$_SDFFE_PN0P_  (.CLK(clknet_leaf_162_clk_p2c),
    .RESET_B(net521),
    .D(_00025_),
    .Q_N(_06776_),
    .Q(\median_processor.input_storage [32]));
 sg13g2_dfrbp_1 \median_processor.input_storage[33]$_SDFFE_PN0P_  (.CLK(clknet_leaf_162_clk_p2c),
    .RESET_B(net522),
    .D(_00026_),
    .Q_N(_06775_),
    .Q(\median_processor.input_storage [33]));
 sg13g2_dfrbp_1 \median_processor.input_storage[34]$_SDFFE_PN0P_  (.CLK(clknet_leaf_172_clk_p2c),
    .RESET_B(net523),
    .D(_00027_),
    .Q_N(_06774_),
    .Q(\median_processor.input_storage [34]));
 sg13g2_dfrbp_1 \median_processor.input_storage[35]$_SDFFE_PN0P_  (.CLK(clknet_leaf_172_clk_p2c),
    .RESET_B(net524),
    .D(_00028_),
    .Q_N(_06773_),
    .Q(\median_processor.input_storage [35]));
 sg13g2_dfrbp_1 \median_processor.input_storage[36]$_SDFFE_PN0P_  (.CLK(clknet_leaf_171_clk_p2c),
    .RESET_B(net525),
    .D(_00029_),
    .Q_N(_06772_),
    .Q(\median_processor.input_storage [36]));
 sg13g2_dfrbp_1 \median_processor.input_storage[37]$_SDFFE_PN0P_  (.CLK(clknet_leaf_169_clk_p2c),
    .RESET_B(net526),
    .D(_00030_),
    .Q_N(_06771_),
    .Q(\median_processor.input_storage [37]));
 sg13g2_dfrbp_1 \median_processor.input_storage[38]$_SDFFE_PN0P_  (.CLK(clknet_leaf_169_clk_p2c),
    .RESET_B(net527),
    .D(_00031_),
    .Q_N(_06770_),
    .Q(\median_processor.input_storage [38]));
 sg13g2_dfrbp_1 \median_processor.input_storage[39]$_SDFFE_PN0P_  (.CLK(clknet_leaf_169_clk_p2c),
    .RESET_B(net528),
    .D(_00032_),
    .Q_N(_06769_),
    .Q(\median_processor.input_storage [39]));
 sg13g2_dfrbp_1 \median_processor.input_storage[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_181_clk_p2c),
    .RESET_B(net529),
    .D(_00033_),
    .Q_N(_06768_),
    .Q(\median_processor.input_storage [3]));
 sg13g2_dfrbp_1 \median_processor.input_storage[40]$_SDFFE_PN0P_  (.CLK(clknet_leaf_173_clk_p2c),
    .RESET_B(net530),
    .D(_00034_),
    .Q_N(_06767_),
    .Q(\median_processor.input_storage [40]));
 sg13g2_dfrbp_1 \median_processor.input_storage[41]$_SDFFE_PN0P_  (.CLK(clknet_leaf_182_clk_p2c),
    .RESET_B(net531),
    .D(_00035_),
    .Q_N(_06766_),
    .Q(\median_processor.input_storage [41]));
 sg13g2_dfrbp_1 \median_processor.input_storage[42]$_SDFFE_PN0P_  (.CLK(clknet_leaf_173_clk_p2c),
    .RESET_B(net532),
    .D(_00036_),
    .Q_N(_06765_),
    .Q(\median_processor.input_storage [42]));
 sg13g2_dfrbp_1 \median_processor.input_storage[43]$_SDFFE_PN0P_  (.CLK(clknet_leaf_182_clk_p2c),
    .RESET_B(net533),
    .D(_00037_),
    .Q_N(_06764_),
    .Q(\median_processor.input_storage [43]));
 sg13g2_dfrbp_1 \median_processor.input_storage[44]$_SDFFE_PN0P_  (.CLK(clknet_leaf_173_clk_p2c),
    .RESET_B(net534),
    .D(_00038_),
    .Q_N(_06763_),
    .Q(\median_processor.input_storage [44]));
 sg13g2_dfrbp_1 \median_processor.input_storage[45]$_SDFFE_PN0P_  (.CLK(clknet_leaf_171_clk_p2c),
    .RESET_B(net535),
    .D(_00039_),
    .Q_N(_06762_),
    .Q(\median_processor.input_storage [45]));
 sg13g2_dfrbp_1 \median_processor.input_storage[46]$_SDFFE_PN0P_  (.CLK(clknet_leaf_170_clk_p2c),
    .RESET_B(net536),
    .D(_00040_),
    .Q_N(_06761_),
    .Q(\median_processor.input_storage [46]));
 sg13g2_dfrbp_1 \median_processor.input_storage[47]$_SDFFE_PN0P_  (.CLK(clknet_leaf_170_clk_p2c),
    .RESET_B(net537),
    .D(_00041_),
    .Q_N(_06760_),
    .Q(\median_processor.input_storage [47]));
 sg13g2_dfrbp_1 \median_processor.input_storage[48]$_SDFFE_PN0P_  (.CLK(clknet_leaf_173_clk_p2c),
    .RESET_B(net538),
    .D(_00042_),
    .Q_N(_06759_),
    .Q(\median_processor.input_storage [48]));
 sg13g2_dfrbp_1 \median_processor.input_storage[49]$_SDFFE_PN0P_  (.CLK(clknet_leaf_161_clk_p2c),
    .RESET_B(net539),
    .D(_00043_),
    .Q_N(_06758_),
    .Q(\median_processor.input_storage [49]));
 sg13g2_dfrbp_1 \median_processor.input_storage[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_174_clk_p2c),
    .RESET_B(net540),
    .D(_00044_),
    .Q_N(_06757_),
    .Q(\median_processor.input_storage [4]));
 sg13g2_dfrbp_1 \median_processor.input_storage[50]$_SDFFE_PN0P_  (.CLK(clknet_leaf_173_clk_p2c),
    .RESET_B(net541),
    .D(_00045_),
    .Q_N(_06756_),
    .Q(\median_processor.input_storage [50]));
 sg13g2_dfrbp_1 \median_processor.input_storage[51]$_SDFFE_PN0P_  (.CLK(clknet_leaf_172_clk_p2c),
    .RESET_B(net542),
    .D(_00046_),
    .Q_N(_06755_),
    .Q(\median_processor.input_storage [51]));
 sg13g2_dfrbp_1 \median_processor.input_storage[52]$_SDFFE_PN0P_  (.CLK(clknet_leaf_171_clk_p2c),
    .RESET_B(net543),
    .D(_00047_),
    .Q_N(_06754_),
    .Q(\median_processor.input_storage [52]));
 sg13g2_dfrbp_1 \median_processor.input_storage[53]$_SDFFE_PN0P_  (.CLK(clknet_leaf_170_clk_p2c),
    .RESET_B(net544),
    .D(_00048_),
    .Q_N(_06753_),
    .Q(\median_processor.input_storage [53]));
 sg13g2_dfrbp_1 \median_processor.input_storage[54]$_SDFFE_PN0P_  (.CLK(clknet_leaf_170_clk_p2c),
    .RESET_B(net545),
    .D(_00049_),
    .Q_N(_06752_),
    .Q(\median_processor.input_storage [54]));
 sg13g2_dfrbp_1 \median_processor.input_storage[55]$_SDFFE_PN0P_  (.CLK(clknet_leaf_171_clk_p2c),
    .RESET_B(net546),
    .D(_00050_),
    .Q_N(_06751_),
    .Q(\median_processor.input_storage [55]));
 sg13g2_dfrbp_1 \median_processor.input_storage[56]$_SDFFE_PN0P_  (.CLK(clknet_leaf_181_clk_p2c),
    .RESET_B(net547),
    .D(_00051_),
    .Q_N(_06750_),
    .Q(\median_processor.input_storage [56]));
 sg13g2_dfrbp_1 \median_processor.input_storage[57]$_SDFFE_PN0P_  (.CLK(clknet_leaf_180_clk_p2c),
    .RESET_B(net548),
    .D(_00052_),
    .Q_N(_06749_),
    .Q(\median_processor.input_storage [57]));
 sg13g2_dfrbp_1 \median_processor.input_storage[58]$_SDFFE_PN0P_  (.CLK(clknet_leaf_180_clk_p2c),
    .RESET_B(net549),
    .D(_00053_),
    .Q_N(_06748_),
    .Q(\median_processor.input_storage [58]));
 sg13g2_dfrbp_1 \median_processor.input_storage[59]$_SDFFE_PN0P_  (.CLK(clknet_leaf_177_clk_p2c),
    .RESET_B(net550),
    .D(_00054_),
    .Q_N(_06747_),
    .Q(\median_processor.input_storage [59]));
 sg13g2_dfrbp_1 \median_processor.input_storage[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_176_clk_p2c),
    .RESET_B(net551),
    .D(_00055_),
    .Q_N(_06746_),
    .Q(\median_processor.input_storage [5]));
 sg13g2_dfrbp_1 \median_processor.input_storage[60]$_SDFFE_PN0P_  (.CLK(clknet_leaf_176_clk_p2c),
    .RESET_B(net552),
    .D(_00056_),
    .Q_N(_06745_),
    .Q(\median_processor.input_storage [60]));
 sg13g2_dfrbp_1 \median_processor.input_storage[61]$_SDFFE_PN0P_  (.CLK(clknet_leaf_176_clk_p2c),
    .RESET_B(net553),
    .D(_00057_),
    .Q_N(_06744_),
    .Q(\median_processor.input_storage [61]));
 sg13g2_dfrbp_1 \median_processor.input_storage[62]$_SDFFE_PN0P_  (.CLK(clknet_leaf_176_clk_p2c),
    .RESET_B(net554),
    .D(_00058_),
    .Q_N(_06743_),
    .Q(\median_processor.input_storage [62]));
 sg13g2_dfrbp_1 \median_processor.input_storage[63]$_SDFFE_PN0P_  (.CLK(clknet_leaf_176_clk_p2c),
    .RESET_B(net555),
    .D(_00059_),
    .Q_N(_06742_),
    .Q(\median_processor.input_storage [63]));
 sg13g2_dfrbp_1 \median_processor.input_storage[6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_175_clk_p2c),
    .RESET_B(net556),
    .D(_00060_),
    .Q_N(_06741_),
    .Q(\median_processor.input_storage [6]));
 sg13g2_dfrbp_1 \median_processor.input_storage[7]$_SDFFE_PN0P_  (.CLK(clknet_leaf_174_clk_p2c),
    .RESET_B(net557),
    .D(_00061_),
    .Q_N(_06740_),
    .Q(\median_processor.input_storage [7]));
 sg13g2_dfrbp_1 \median_processor.input_storage[8]$_SDFFE_PN0P_  (.CLK(clknet_leaf_181_clk_p2c),
    .RESET_B(net558),
    .D(_00062_),
    .Q_N(_06739_),
    .Q(\median_processor.input_storage [8]));
 sg13g2_dfrbp_1 \median_processor.input_storage[9]$_SDFFE_PN0P_  (.CLK(clknet_leaf_181_clk_p2c),
    .RESET_B(net559),
    .D(_00063_),
    .Q_N(_06738_),
    .Q(\median_processor.input_storage [9]));
 sg13g2_dfrbp_1 \median_processor.median_processor.median_out[0]$_DFFE_PP_  (.CLK(clknet_leaf_179_clk_p2c),
    .RESET_B(net560),
    .D(_00064_),
    .Q_N(_06737_),
    .Q(\median_processor.median_processor.median_out [0]));
 sg13g2_dfrbp_1 \median_processor.median_processor.median_out[1]$_DFFE_PP_  (.CLK(clknet_leaf_180_clk_p2c),
    .RESET_B(net561),
    .D(_00065_),
    .Q_N(_06736_),
    .Q(\median_processor.median_processor.median_out [1]));
 sg13g2_dfrbp_1 \median_processor.median_processor.median_out[2]$_DFFE_PP_  (.CLK(clknet_leaf_180_clk_p2c),
    .RESET_B(net562),
    .D(_00066_),
    .Q_N(_06735_),
    .Q(\median_processor.median_processor.median_out [2]));
 sg13g2_dfrbp_1 \median_processor.median_processor.median_out[3]$_DFFE_PP_  (.CLK(clknet_leaf_177_clk_p2c),
    .RESET_B(net563),
    .D(_00067_),
    .Q_N(_06734_),
    .Q(\median_processor.median_processor.median_out [3]));
 sg13g2_dfrbp_1 \median_processor.median_processor.median_out[4]$_DFFE_PP_  (.CLK(clknet_leaf_177_clk_p2c),
    .RESET_B(net564),
    .D(_00068_),
    .Q_N(_06733_),
    .Q(\median_processor.median_processor.median_out [4]));
 sg13g2_dfrbp_1 \median_processor.median_processor.median_out[5]$_DFFE_PP_  (.CLK(clknet_leaf_175_clk_p2c),
    .RESET_B(net565),
    .D(_00069_),
    .Q_N(_06732_),
    .Q(\median_processor.median_processor.median_out [5]));
 sg13g2_dfrbp_1 \median_processor.median_processor.median_out[6]$_DFFE_PP_  (.CLK(clknet_leaf_175_clk_p2c),
    .RESET_B(net566),
    .D(_00070_),
    .Q_N(_06731_),
    .Q(\median_processor.median_processor.median_out [6]));
 sg13g2_dfrbp_1 \median_processor.median_processor.median_out[7]$_DFFE_PP_  (.CLK(clknet_leaf_175_clk_p2c),
    .RESET_B(net567),
    .D(_00071_),
    .Q_N(_06730_),
    .Q(\median_processor.median_processor.median_out [7]));
 sg13g2_IOPadIn port_aux_enable_cell (.p2c(aux_enable_p2c),
    .pad(aux_enable_pad));
 sg13g2_IOPadIn port_clk_cell (.p2c(clk_p2c),
    .pad(clk_pad));
 sg13g2_IOPadIn port_data_in1_cell (.p2c(data_in_p2c_1),
    .pad(data_in_pad[0]));
 sg13g2_IOPadIn port_data_in2_cell (.p2c(data_in_p2c_2),
    .pad(data_in_pad[1]));
 sg13g2_IOPadIn port_data_in3_cell (.p2c(data_in_p2c_3),
    .pad(data_in_pad[2]));
 sg13g2_IOPadIn port_data_in4_cell (.p2c(data_in_p2c_4),
    .pad(data_in_pad[3]));
 sg13g2_IOPadIn port_data_in5_cell (.p2c(data_in_p2c_5),
    .pad(data_in_pad[4]));
 sg13g2_IOPadIn port_data_in6_cell (.p2c(data_in_p2c_6),
    .pad(data_in_pad[5]));
 sg13g2_IOPadIn port_data_in7_cell (.p2c(data_in_p2c_7),
    .pad(data_in_pad[6]));
 sg13g2_IOPadIn port_data_in8_cell (.p2c(data_in_p2c_8),
    .pad(data_in_pad[7]));
 sg13g2_IOPadOut16mA port_data_out1_cell (.c2p(data_out_c2p[0]),
    .pad(data_out_pad[0]));
 sg13g2_IOPadOut16mA port_data_out2_cell (.c2p(data_out_c2p[1]),
    .pad(data_out_pad[1]));
 sg13g2_IOPadOut16mA port_data_out3_cell (.c2p(data_out_c2p[2]),
    .pad(data_out_pad[2]));
 sg13g2_IOPadOut16mA port_data_out4_cell (.c2p(data_out_c2p[3]),
    .pad(data_out_pad[3]));
 sg13g2_IOPadOut16mA port_data_out5_cell (.c2p(data_out_c2p[4]),
    .pad(data_out_pad[4]));
 sg13g2_IOPadOut16mA port_data_out6_cell (.c2p(data_out_c2p[5]),
    .pad(data_out_pad[5]));
 sg13g2_IOPadOut16mA port_data_out7_cell (.c2p(data_out_c2p[6]),
    .pad(data_out_pad[6]));
 sg13g2_IOPadOut16mA port_data_out8_cell (.c2p(data_out_c2p[7]),
    .pad(data_out_pad[7]));
 sg13g2_IOPadOut16mA port_lfsr_out_cell (.c2p(lfsr_out_c2p),
    .pad(lfsr_out_pad));
 sg13g2_IOPadIn port_out_select1_cell (.p2c(out_select_p2c_1),
    .pad(out_select_pad[0]));
 sg13g2_IOPadIn port_out_select2_cell (.p2c(out_select_p2c_2),
    .pad(out_select_pad[1]));
 sg13g2_IOPadIn port_reg_addr1_cell (.p2c(reg_addr_p2c_1),
    .pad(reg_addr_pad[0]));
 sg13g2_IOPadIn port_reg_addr2_cell (.p2c(reg_addr_p2c_2),
    .pad(reg_addr_pad[1]));
 sg13g2_IOPadIn port_reg_addr3_cell (.p2c(reg_addr_p2c_3),
    .pad(reg_addr_pad[2]));
 sg13g2_IOPadIn port_rst_cell (.p2c(\median_processor.rst ),
    .pad(rst_pad));
 sg13g2_IOPadIn port_shreg_in_cell (.p2c(\shift_storage.shreg_in ),
    .pad(shreg_in_pad));
 sg13g2_IOPadOut16mA port_shreg_out_cell (.c2p(\shift_storage.shreg_out ),
    .pad(shreg_out_pad));
 sg13g2_IOPadIn port_wr_enable_cell (.p2c(\median_processor.wr_enable ),
    .pad(wr_enable_pad));
 sg13g2_dfrbp_1 \rando_generator.lfsr_reg[0]$_SDFF_PN0_  (.CLK(clknet_leaf_86_clk_p2c),
    .RESET_B(net568),
    .D(_00072_),
    .Q_N(_06729_),
    .Q(lfsr_out_c2p));
 sg13g2_dfrbp_1 \rando_generator.lfsr_reg[10]$_SDFF_PN0_  (.CLK(clknet_leaf_83_clk_p2c),
    .RESET_B(net569),
    .D(_00073_),
    .Q_N(_06728_),
    .Q(\rando_generator.lfsr_reg [10]));
 sg13g2_dfrbp_1 \rando_generator.lfsr_reg[11]$_SDFF_PN0_  (.CLK(clknet_leaf_83_clk_p2c),
    .RESET_B(net570),
    .D(_00074_),
    .Q_N(_06727_),
    .Q(\rando_generator.lfsr_reg [11]));
 sg13g2_dfrbp_1 \rando_generator.lfsr_reg[12]$_SDFF_PN0_  (.CLK(clknet_leaf_83_clk_p2c),
    .RESET_B(net571),
    .D(_00075_),
    .Q_N(_06726_),
    .Q(\rando_generator.lfsr_reg [12]));
 sg13g2_dfrbp_1 \rando_generator.lfsr_reg[13]$_SDFF_PN0_  (.CLK(clknet_leaf_89_clk_p2c),
    .RESET_B(net572),
    .D(_00076_),
    .Q_N(_06725_),
    .Q(\rando_generator.lfsr_reg [13]));
 sg13g2_dfrbp_1 \rando_generator.lfsr_reg[14]$_SDFF_PN0_  (.CLK(clknet_leaf_89_clk_p2c),
    .RESET_B(net573),
    .D(_00077_),
    .Q_N(_06724_),
    .Q(\rando_generator.lfsr_reg [14]));
 sg13g2_dfrbp_1 \rando_generator.lfsr_reg[15]$_SDFF_PN0_  (.CLK(clknet_leaf_89_clk_p2c),
    .RESET_B(net574),
    .D(_00078_),
    .Q_N(_06723_),
    .Q(\rando_generator.lfsr_reg [15]));
 sg13g2_dfrbp_1 \rando_generator.lfsr_reg[16]$_SDFF_PN0_  (.CLK(clknet_leaf_87_clk_p2c),
    .RESET_B(net575),
    .D(_00079_),
    .Q_N(_06722_),
    .Q(\rando_generator.lfsr_reg [16]));
 sg13g2_dfrbp_1 \rando_generator.lfsr_reg[17]$_SDFF_PN0_  (.CLK(clknet_leaf_87_clk_p2c),
    .RESET_B(net576),
    .D(_00080_),
    .Q_N(_06721_),
    .Q(\rando_generator.lfsr_reg [17]));
 sg13g2_dfrbp_1 \rando_generator.lfsr_reg[18]$_SDFF_PN0_  (.CLK(clknet_leaf_87_clk_p2c),
    .RESET_B(net577),
    .D(_00081_),
    .Q_N(_06720_),
    .Q(\rando_generator.lfsr_reg [18]));
 sg13g2_dfrbp_1 \rando_generator.lfsr_reg[19]$_SDFF_PN0_  (.CLK(clknet_leaf_86_clk_p2c),
    .RESET_B(net578),
    .D(_00082_),
    .Q_N(_06719_),
    .Q(\rando_generator.lfsr_reg [19]));
 sg13g2_dfrbp_1 \rando_generator.lfsr_reg[1]$_SDFF_PN0_  (.CLK(clknet_leaf_84_clk_p2c),
    .RESET_B(net579),
    .D(_00083_),
    .Q_N(_06718_),
    .Q(\rando_generator.lfsr_reg [1]));
 sg13g2_dfrbp_1 \rando_generator.lfsr_reg[20]$_SDFF_PN0_  (.CLK(clknet_leaf_86_clk_p2c),
    .RESET_B(net580),
    .D(_00084_),
    .Q_N(_06717_),
    .Q(\rando_generator.lfsr_reg [20]));
 sg13g2_dfrbp_1 \rando_generator.lfsr_reg[21]$_SDFF_PN0_  (.CLK(clknet_leaf_87_clk_p2c),
    .RESET_B(net581),
    .D(_00085_),
    .Q_N(_06716_),
    .Q(\rando_generator.lfsr_reg [21]));
 sg13g2_dfrbp_1 \rando_generator.lfsr_reg[22]$_SDFF_PN0_  (.CLK(clknet_leaf_86_clk_p2c),
    .RESET_B(net582),
    .D(_00086_),
    .Q_N(_06715_),
    .Q(\rando_generator.lfsr_reg [22]));
 sg13g2_dfrbp_1 \rando_generator.lfsr_reg[23]$_SDFF_PN0_  (.CLK(clknet_leaf_86_clk_p2c),
    .RESET_B(net583),
    .D(_00087_),
    .Q_N(_06714_),
    .Q(\rando_generator.lfsr_reg [23]));
 sg13g2_dfrbp_1 \rando_generator.lfsr_reg[24]$_SDFF_PN0_  (.CLK(clknet_leaf_86_clk_p2c),
    .RESET_B(net584),
    .D(_00088_),
    .Q_N(_06713_),
    .Q(\rando_generator.lfsr_reg [24]));
 sg13g2_dfrbp_1 \rando_generator.lfsr_reg[25]$_SDFF_PN0_  (.CLK(clknet_leaf_86_clk_p2c),
    .RESET_B(net585),
    .D(_00089_),
    .Q_N(_06712_),
    .Q(\rando_generator.lfsr_reg [25]));
 sg13g2_dfrbp_1 \rando_generator.lfsr_reg[26]$_SDFF_PN0_  (.CLK(clknet_leaf_85_clk_p2c),
    .RESET_B(net586),
    .D(_00090_),
    .Q_N(_06711_),
    .Q(\rando_generator.lfsr_reg [26]));
 sg13g2_dfrbp_1 \rando_generator.lfsr_reg[27]$_SDFF_PN0_  (.CLK(clknet_leaf_85_clk_p2c),
    .RESET_B(net587),
    .D(_00091_),
    .Q_N(_06710_),
    .Q(\rando_generator.lfsr_reg [27]));
 sg13g2_dfrbp_1 \rando_generator.lfsr_reg[28]$_SDFF_PN0_  (.CLK(clknet_leaf_85_clk_p2c),
    .RESET_B(net588),
    .D(_00092_),
    .Q_N(_06709_),
    .Q(\rando_generator.lfsr_reg [28]));
 sg13g2_dfrbp_1 \rando_generator.lfsr_reg[29]$_SDFF_PN0_  (.CLK(clknet_leaf_85_clk_p2c),
    .RESET_B(net589),
    .D(_00093_),
    .Q_N(_06708_),
    .Q(\rando_generator.lfsr_reg [29]));
 sg13g2_dfrbp_1 \rando_generator.lfsr_reg[2]$_SDFF_PN0_  (.CLK(clknet_leaf_84_clk_p2c),
    .RESET_B(net590),
    .D(_00094_),
    .Q_N(_06707_),
    .Q(\rando_generator.lfsr_reg [2]));
 sg13g2_dfrbp_1 \rando_generator.lfsr_reg[30]$_SDFF_PN0_  (.CLK(clknet_leaf_85_clk_p2c),
    .RESET_B(net591),
    .D(_00095_),
    .Q_N(_06706_),
    .Q(\rando_generator.lfsr_reg [30]));
 sg13g2_dfrbp_1 \rando_generator.lfsr_reg[3]$_SDFF_PN0_  (.CLK(clknet_leaf_85_clk_p2c),
    .RESET_B(net592),
    .D(_00096_),
    .Q_N(_06705_),
    .Q(\rando_generator.lfsr_reg [3]));
 sg13g2_dfrbp_1 \rando_generator.lfsr_reg[4]$_SDFF_PN0_  (.CLK(clknet_leaf_84_clk_p2c),
    .RESET_B(net593),
    .D(_00097_),
    .Q_N(_06704_),
    .Q(\rando_generator.lfsr_reg [4]));
 sg13g2_dfrbp_1 \rando_generator.lfsr_reg[5]$_SDFF_PN0_  (.CLK(clknet_leaf_84_clk_p2c),
    .RESET_B(net594),
    .D(_00098_),
    .Q_N(_06703_),
    .Q(\rando_generator.lfsr_reg [5]));
 sg13g2_dfrbp_1 \rando_generator.lfsr_reg[6]$_SDFF_PN0_  (.CLK(clknet_leaf_84_clk_p2c),
    .RESET_B(net595),
    .D(_00099_),
    .Q_N(_06702_),
    .Q(\rando_generator.lfsr_reg [6]));
 sg13g2_dfrbp_1 \rando_generator.lfsr_reg[7]$_SDFF_PN0_  (.CLK(clknet_leaf_83_clk_p2c),
    .RESET_B(net596),
    .D(_00100_),
    .Q_N(_06701_),
    .Q(\rando_generator.lfsr_reg [7]));
 sg13g2_dfrbp_1 \rando_generator.lfsr_reg[8]$_SDFF_PN0_  (.CLK(clknet_leaf_83_clk_p2c),
    .RESET_B(net597),
    .D(_00101_),
    .Q_N(_06700_),
    .Q(\rando_generator.lfsr_reg [8]));
 sg13g2_dfrbp_1 \rando_generator.lfsr_reg[9]$_SDFF_PN0_  (.CLK(clknet_leaf_83_clk_p2c),
    .RESET_B(net598),
    .D(_00102_),
    .Q_N(_06699_),
    .Q(\rando_generator.lfsr_reg [9]));
 sg13g2_dfrbp_1 \shift_storage.storage[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_122_clk_p2c),
    .RESET_B(net599),
    .D(_00103_),
    .Q_N(_06698_),
    .Q(\shift_storage.storage [0]));
 sg13g2_dfrbp_1 \shift_storage.storage[1000]$_SDFFE_PN0P_  (.CLK(clknet_leaf_48_clk_p2c),
    .RESET_B(net600),
    .D(_00104_),
    .Q_N(_06697_),
    .Q(\shift_storage.storage [1000]));
 sg13g2_dfrbp_1 \shift_storage.storage[1001]$_SDFFE_PN0P_  (.CLK(clknet_leaf_48_clk_p2c),
    .RESET_B(net601),
    .D(_00105_),
    .Q_N(_06696_),
    .Q(\shift_storage.storage [1001]));
 sg13g2_dfrbp_1 \shift_storage.storage[1002]$_SDFFE_PN0P_  (.CLK(clknet_leaf_48_clk_p2c),
    .RESET_B(net602),
    .D(_00106_),
    .Q_N(_06695_),
    .Q(\shift_storage.storage [1002]));
 sg13g2_dfrbp_1 \shift_storage.storage[1003]$_SDFFE_PN0P_  (.CLK(clknet_leaf_122_clk_p2c),
    .RESET_B(net603),
    .D(_00107_),
    .Q_N(_06694_),
    .Q(\shift_storage.storage [1003]));
 sg13g2_dfrbp_1 \shift_storage.storage[1004]$_SDFFE_PN0P_  (.CLK(clknet_leaf_122_clk_p2c),
    .RESET_B(net604),
    .D(_00108_),
    .Q_N(_06693_),
    .Q(\shift_storage.storage [1004]));
 sg13g2_dfrbp_1 \shift_storage.storage[1005]$_SDFFE_PN0P_  (.CLK(clknet_leaf_50_clk_p2c),
    .RESET_B(net605),
    .D(_00109_),
    .Q_N(_06692_),
    .Q(\shift_storage.storage [1005]));
 sg13g2_dfrbp_1 \shift_storage.storage[1006]$_SDFFE_PN0P_  (.CLK(clknet_leaf_50_clk_p2c),
    .RESET_B(net606),
    .D(_00110_),
    .Q_N(_06691_),
    .Q(\shift_storage.storage [1006]));
 sg13g2_dfrbp_1 \shift_storage.storage[1007]$_SDFFE_PN0P_  (.CLK(clknet_leaf_49_clk_p2c),
    .RESET_B(net607),
    .D(_00111_),
    .Q_N(_06690_),
    .Q(\shift_storage.storage [1007]));
 sg13g2_dfrbp_1 \shift_storage.storage[1008]$_SDFFE_PN0P_  (.CLK(clknet_leaf_49_clk_p2c),
    .RESET_B(net608),
    .D(_00112_),
    .Q_N(_06689_),
    .Q(\shift_storage.storage [1008]));
 sg13g2_dfrbp_1 \shift_storage.storage[1009]$_SDFFE_PN0P_  (.CLK(clknet_leaf_49_clk_p2c),
    .RESET_B(net609),
    .D(_00113_),
    .Q_N(_06688_),
    .Q(\shift_storage.storage [1009]));
 sg13g2_dfrbp_1 \shift_storage.storage[100]$_SDFFE_PN0P_  (.CLK(clknet_leaf_49_clk_p2c),
    .RESET_B(net610),
    .D(_00114_),
    .Q_N(_06687_),
    .Q(\shift_storage.storage [100]));
 sg13g2_dfrbp_1 \shift_storage.storage[1010]$_SDFFE_PN0P_  (.CLK(clknet_leaf_48_clk_p2c),
    .RESET_B(net611),
    .D(_00115_),
    .Q_N(_06686_),
    .Q(\shift_storage.storage [1010]));
 sg13g2_dfrbp_1 \shift_storage.storage[1011]$_SDFFE_PN0P_  (.CLK(clknet_leaf_49_clk_p2c),
    .RESET_B(net612),
    .D(_00116_),
    .Q_N(_06685_),
    .Q(\shift_storage.storage [1011]));
 sg13g2_dfrbp_1 \shift_storage.storage[1012]$_SDFFE_PN0P_  (.CLK(clknet_leaf_49_clk_p2c),
    .RESET_B(net613),
    .D(_00117_),
    .Q_N(_06684_),
    .Q(\shift_storage.storage [1012]));
 sg13g2_dfrbp_1 \shift_storage.storage[1013]$_SDFFE_PN0P_  (.CLK(clknet_leaf_46_clk_p2c),
    .RESET_B(net614),
    .D(_00118_),
    .Q_N(_06683_),
    .Q(\shift_storage.storage [1013]));
 sg13g2_dfrbp_1 \shift_storage.storage[1014]$_SDFFE_PN0P_  (.CLK(clknet_leaf_46_clk_p2c),
    .RESET_B(net615),
    .D(_00119_),
    .Q_N(_06682_),
    .Q(\shift_storage.storage [1014]));
 sg13g2_dfrbp_1 \shift_storage.storage[1015]$_SDFFE_PN0P_  (.CLK(clknet_leaf_43_clk_p2c),
    .RESET_B(net616),
    .D(_00120_),
    .Q_N(_06681_),
    .Q(\shift_storage.storage [1015]));
 sg13g2_dfrbp_1 \shift_storage.storage[1016]$_SDFFE_PN0P_  (.CLK(clknet_leaf_51_clk_p2c),
    .RESET_B(net617),
    .D(_00121_),
    .Q_N(_06680_),
    .Q(\shift_storage.storage [1016]));
 sg13g2_dfrbp_1 \shift_storage.storage[1017]$_SDFFE_PN0P_  (.CLK(clknet_leaf_51_clk_p2c),
    .RESET_B(net618),
    .D(_00122_),
    .Q_N(_06679_),
    .Q(\shift_storage.storage [1017]));
 sg13g2_dfrbp_1 \shift_storage.storage[1018]$_SDFFE_PN0P_  (.CLK(clknet_leaf_42_clk_p2c),
    .RESET_B(net619),
    .D(_00123_),
    .Q_N(_06678_),
    .Q(\shift_storage.storage [1018]));
 sg13g2_dfrbp_1 \shift_storage.storage[1019]$_SDFFE_PN0P_  (.CLK(clknet_leaf_42_clk_p2c),
    .RESET_B(net620),
    .D(_00124_),
    .Q_N(_06677_),
    .Q(\shift_storage.storage [1019]));
 sg13g2_dfrbp_1 \shift_storage.storage[101]$_SDFFE_PN0P_  (.CLK(clknet_leaf_51_clk_p2c),
    .RESET_B(net621),
    .D(_00125_),
    .Q_N(_06676_),
    .Q(\shift_storage.storage [101]));
 sg13g2_dfrbp_1 \shift_storage.storage[1020]$_SDFFE_PN0P_  (.CLK(clknet_leaf_41_clk_p2c),
    .RESET_B(net622),
    .D(_00126_),
    .Q_N(_06675_),
    .Q(\shift_storage.storage [1020]));
 sg13g2_dfrbp_1 \shift_storage.storage[1021]$_SDFFE_PN0P_  (.CLK(clknet_leaf_52_clk_p2c),
    .RESET_B(net623),
    .D(_00127_),
    .Q_N(_06674_),
    .Q(\shift_storage.storage [1021]));
 sg13g2_dfrbp_1 \shift_storage.storage[1022]$_SDFFE_PN0P_  (.CLK(clknet_leaf_52_clk_p2c),
    .RESET_B(net624),
    .D(_00128_),
    .Q_N(_06673_),
    .Q(\shift_storage.storage [1022]));
 sg13g2_dfrbp_1 \shift_storage.storage[1023]$_SDFFE_PN0P_  (.CLK(clknet_leaf_52_clk_p2c),
    .RESET_B(net625),
    .D(_00129_),
    .Q_N(_06672_),
    .Q(\shift_storage.storage [1023]));
 sg13g2_dfrbp_1 \shift_storage.storage[1024]$_SDFFE_PN0P_  (.CLK(clknet_leaf_52_clk_p2c),
    .RESET_B(net626),
    .D(_00130_),
    .Q_N(_06671_),
    .Q(\shift_storage.storage [1024]));
 sg13g2_dfrbp_1 \shift_storage.storage[1025]$_SDFFE_PN0P_  (.CLK(clknet_leaf_51_clk_p2c),
    .RESET_B(net627),
    .D(_00131_),
    .Q_N(_06670_),
    .Q(\shift_storage.storage [1025]));
 sg13g2_dfrbp_1 \shift_storage.storage[1026]$_SDFFE_PN0P_  (.CLK(clknet_leaf_51_clk_p2c),
    .RESET_B(net628),
    .D(_00132_),
    .Q_N(_06669_),
    .Q(\shift_storage.storage [1026]));
 sg13g2_dfrbp_1 \shift_storage.storage[1027]$_SDFFE_PN0P_  (.CLK(clknet_leaf_51_clk_p2c),
    .RESET_B(net629),
    .D(_00133_),
    .Q_N(_06668_),
    .Q(\shift_storage.storage [1027]));
 sg13g2_dfrbp_1 \shift_storage.storage[1028]$_SDFFE_PN0P_  (.CLK(clknet_leaf_53_clk_p2c),
    .RESET_B(net630),
    .D(_00134_),
    .Q_N(_06667_),
    .Q(\shift_storage.storage [1028]));
 sg13g2_dfrbp_1 \shift_storage.storage[1029]$_SDFFE_PN0P_  (.CLK(clknet_leaf_53_clk_p2c),
    .RESET_B(net631),
    .D(_00135_),
    .Q_N(_06666_),
    .Q(\shift_storage.storage [1029]));
 sg13g2_dfrbp_1 \shift_storage.storage[102]$_SDFFE_PN0P_  (.CLK(clknet_leaf_50_clk_p2c),
    .RESET_B(net632),
    .D(_00136_),
    .Q_N(_06665_),
    .Q(\shift_storage.storage [102]));
 sg13g2_dfrbp_1 \shift_storage.storage[1030]$_SDFFE_PN0P_  (.CLK(clknet_leaf_55_clk_p2c),
    .RESET_B(net633),
    .D(_00137_),
    .Q_N(_06664_),
    .Q(\shift_storage.storage [1030]));
 sg13g2_dfrbp_1 \shift_storage.storage[1031]$_SDFFE_PN0P_  (.CLK(clknet_leaf_51_clk_p2c),
    .RESET_B(net634),
    .D(_00138_),
    .Q_N(_06663_),
    .Q(\shift_storage.storage [1031]));
 sg13g2_dfrbp_1 \shift_storage.storage[1032]$_SDFFE_PN0P_  (.CLK(clknet_leaf_55_clk_p2c),
    .RESET_B(net635),
    .D(_00139_),
    .Q_N(_06662_),
    .Q(\shift_storage.storage [1032]));
 sg13g2_dfrbp_1 \shift_storage.storage[1033]$_SDFFE_PN0P_  (.CLK(clknet_leaf_55_clk_p2c),
    .RESET_B(net636),
    .D(_00140_),
    .Q_N(_06661_),
    .Q(\shift_storage.storage [1033]));
 sg13g2_dfrbp_1 \shift_storage.storage[1034]$_SDFFE_PN0P_  (.CLK(clknet_leaf_50_clk_p2c),
    .RESET_B(net637),
    .D(_00141_),
    .Q_N(_06660_),
    .Q(\shift_storage.storage [1034]));
 sg13g2_dfrbp_1 \shift_storage.storage[1035]$_SDFFE_PN0P_  (.CLK(clknet_leaf_50_clk_p2c),
    .RESET_B(net638),
    .D(_00142_),
    .Q_N(_06659_),
    .Q(\shift_storage.storage [1035]));
 sg13g2_dfrbp_1 \shift_storage.storage[1036]$_SDFFE_PN0P_  (.CLK(clknet_leaf_50_clk_p2c),
    .RESET_B(net639),
    .D(_00143_),
    .Q_N(_06658_),
    .Q(\shift_storage.storage [1036]));
 sg13g2_dfrbp_1 \shift_storage.storage[1037]$_SDFFE_PN0P_  (.CLK(clknet_leaf_55_clk_p2c),
    .RESET_B(net640),
    .D(_00144_),
    .Q_N(_06657_),
    .Q(\shift_storage.storage [1037]));
 sg13g2_dfrbp_1 \shift_storage.storage[1038]$_SDFFE_PN0P_  (.CLK(clknet_leaf_56_clk_p2c),
    .RESET_B(net641),
    .D(_00145_),
    .Q_N(_06656_),
    .Q(\shift_storage.storage [1038]));
 sg13g2_dfrbp_1 \shift_storage.storage[1039]$_SDFFE_PN0P_  (.CLK(clknet_leaf_56_clk_p2c),
    .RESET_B(net642),
    .D(_00146_),
    .Q_N(_06655_),
    .Q(\shift_storage.storage [1039]));
 sg13g2_dfrbp_1 \shift_storage.storage[103]$_SDFFE_PN0P_  (.CLK(clknet_leaf_50_clk_p2c),
    .RESET_B(net643),
    .D(_00147_),
    .Q_N(_06654_),
    .Q(\shift_storage.storage [103]));
 sg13g2_dfrbp_1 \shift_storage.storage[1040]$_SDFFE_PN0P_  (.CLK(clknet_leaf_116_clk_p2c),
    .RESET_B(net644),
    .D(_00148_),
    .Q_N(_06653_),
    .Q(\shift_storage.storage [1040]));
 sg13g2_dfrbp_1 \shift_storage.storage[1041]$_SDFFE_PN0P_  (.CLK(clknet_leaf_116_clk_p2c),
    .RESET_B(net645),
    .D(_00149_),
    .Q_N(_06652_),
    .Q(\shift_storage.storage [1041]));
 sg13g2_dfrbp_1 \shift_storage.storage[1042]$_SDFFE_PN0P_  (.CLK(clknet_leaf_122_clk_p2c),
    .RESET_B(net646),
    .D(_00150_),
    .Q_N(_06651_),
    .Q(\shift_storage.storage [1042]));
 sg13g2_dfrbp_1 \shift_storage.storage[1043]$_SDFFE_PN0P_  (.CLK(clknet_leaf_122_clk_p2c),
    .RESET_B(net647),
    .D(_00151_),
    .Q_N(_06650_),
    .Q(\shift_storage.storage [1043]));
 sg13g2_dfrbp_1 \shift_storage.storage[1044]$_SDFFE_PN0P_  (.CLK(clknet_leaf_121_clk_p2c),
    .RESET_B(net648),
    .D(_00152_),
    .Q_N(_06649_),
    .Q(\shift_storage.storage [1044]));
 sg13g2_dfrbp_1 \shift_storage.storage[1045]$_SDFFE_PN0P_  (.CLK(clknet_leaf_121_clk_p2c),
    .RESET_B(net649),
    .D(_00153_),
    .Q_N(_06648_),
    .Q(\shift_storage.storage [1045]));
 sg13g2_dfrbp_1 \shift_storage.storage[1046]$_SDFFE_PN0P_  (.CLK(clknet_leaf_116_clk_p2c),
    .RESET_B(net650),
    .D(_00154_),
    .Q_N(_06647_),
    .Q(\shift_storage.storage [1046]));
 sg13g2_dfrbp_1 \shift_storage.storage[1047]$_SDFFE_PN0P_  (.CLK(clknet_leaf_116_clk_p2c),
    .RESET_B(net651),
    .D(_00155_),
    .Q_N(_06646_),
    .Q(\shift_storage.storage [1047]));
 sg13g2_dfrbp_1 \shift_storage.storage[1048]$_SDFFE_PN0P_  (.CLK(clknet_leaf_116_clk_p2c),
    .RESET_B(net652),
    .D(_00156_),
    .Q_N(_06645_),
    .Q(\shift_storage.storage [1048]));
 sg13g2_dfrbp_1 \shift_storage.storage[1049]$_SDFFE_PN0P_  (.CLK(clknet_leaf_117_clk_p2c),
    .RESET_B(net653),
    .D(_00157_),
    .Q_N(_06644_),
    .Q(\shift_storage.storage [1049]));
 sg13g2_dfrbp_1 \shift_storage.storage[104]$_SDFFE_PN0P_  (.CLK(clknet_leaf_122_clk_p2c),
    .RESET_B(net654),
    .D(_00158_),
    .Q_N(_06643_),
    .Q(\shift_storage.storage [104]));
 sg13g2_dfrbp_1 \shift_storage.storage[1050]$_SDFFE_PN0P_  (.CLK(clknet_leaf_121_clk_p2c),
    .RESET_B(net655),
    .D(_00159_),
    .Q_N(_06642_),
    .Q(\shift_storage.storage [1050]));
 sg13g2_dfrbp_1 \shift_storage.storage[1051]$_SDFFE_PN0P_  (.CLK(clknet_leaf_121_clk_p2c),
    .RESET_B(net656),
    .D(_00160_),
    .Q_N(_06641_),
    .Q(\shift_storage.storage [1051]));
 sg13g2_dfrbp_1 \shift_storage.storage[1052]$_SDFFE_PN0P_  (.CLK(clknet_leaf_120_clk_p2c),
    .RESET_B(net657),
    .D(_00161_),
    .Q_N(_06640_),
    .Q(\shift_storage.storage [1052]));
 sg13g2_dfrbp_1 \shift_storage.storage[1053]$_SDFFE_PN0P_  (.CLK(clknet_leaf_119_clk_p2c),
    .RESET_B(net658),
    .D(_00162_),
    .Q_N(_06639_),
    .Q(\shift_storage.storage [1053]));
 sg13g2_dfrbp_1 \shift_storage.storage[1054]$_SDFFE_PN0P_  (.CLK(clknet_leaf_119_clk_p2c),
    .RESET_B(net659),
    .D(_00163_),
    .Q_N(_06638_),
    .Q(\shift_storage.storage [1054]));
 sg13g2_dfrbp_1 \shift_storage.storage[1055]$_SDFFE_PN0P_  (.CLK(clknet_leaf_120_clk_p2c),
    .RESET_B(net660),
    .D(_00164_),
    .Q_N(_06637_),
    .Q(\shift_storage.storage [1055]));
 sg13g2_dfrbp_1 \shift_storage.storage[1056]$_SDFFE_PN0P_  (.CLK(clknet_leaf_120_clk_p2c),
    .RESET_B(net661),
    .D(_00165_),
    .Q_N(_06636_),
    .Q(\shift_storage.storage [1056]));
 sg13g2_dfrbp_1 \shift_storage.storage[1057]$_SDFFE_PN0P_  (.CLK(clknet_leaf_120_clk_p2c),
    .RESET_B(net662),
    .D(_00166_),
    .Q_N(_06635_),
    .Q(\shift_storage.storage [1057]));
 sg13g2_dfrbp_1 \shift_storage.storage[1058]$_SDFFE_PN0P_  (.CLK(clknet_leaf_120_clk_p2c),
    .RESET_B(net663),
    .D(_00167_),
    .Q_N(_06634_),
    .Q(\shift_storage.storage [1058]));
 sg13g2_dfrbp_1 \shift_storage.storage[1059]$_SDFFE_PN0P_  (.CLK(clknet_leaf_120_clk_p2c),
    .RESET_B(net664),
    .D(_00168_),
    .Q_N(_06633_),
    .Q(\shift_storage.storage [1059]));
 sg13g2_dfrbp_1 \shift_storage.storage[105]$_SDFFE_PN0P_  (.CLK(clknet_leaf_123_clk_p2c),
    .RESET_B(net665),
    .D(_00169_),
    .Q_N(_06632_),
    .Q(\shift_storage.storage [105]));
 sg13g2_dfrbp_1 \shift_storage.storage[1060]$_SDFFE_PN0P_  (.CLK(clknet_leaf_123_clk_p2c),
    .RESET_B(net666),
    .D(_00170_),
    .Q_N(_06631_),
    .Q(\shift_storage.storage [1060]));
 sg13g2_dfrbp_1 \shift_storage.storage[1061]$_SDFFE_PN0P_  (.CLK(clknet_leaf_123_clk_p2c),
    .RESET_B(net667),
    .D(_00171_),
    .Q_N(_06630_),
    .Q(\shift_storage.storage [1061]));
 sg13g2_dfrbp_1 \shift_storage.storage[1062]$_SDFFE_PN0P_  (.CLK(clknet_leaf_123_clk_p2c),
    .RESET_B(net668),
    .D(_00172_),
    .Q_N(_06629_),
    .Q(\shift_storage.storage [1062]));
 sg13g2_dfrbp_1 \shift_storage.storage[1063]$_SDFFE_PN0P_  (.CLK(clknet_leaf_123_clk_p2c),
    .RESET_B(net669),
    .D(_00173_),
    .Q_N(_06628_),
    .Q(\shift_storage.storage [1063]));
 sg13g2_dfrbp_1 \shift_storage.storage[1064]$_SDFFE_PN0P_  (.CLK(clknet_leaf_123_clk_p2c),
    .RESET_B(net670),
    .D(_00174_),
    .Q_N(_06627_),
    .Q(\shift_storage.storage [1064]));
 sg13g2_dfrbp_1 \shift_storage.storage[1065]$_SDFFE_PN0P_  (.CLK(clknet_leaf_126_clk_p2c),
    .RESET_B(net671),
    .D(_00175_),
    .Q_N(_06626_),
    .Q(\shift_storage.storage [1065]));
 sg13g2_dfrbp_1 \shift_storage.storage[1066]$_SDFFE_PN0P_  (.CLK(clknet_leaf_126_clk_p2c),
    .RESET_B(net672),
    .D(_00176_),
    .Q_N(_06625_),
    .Q(\shift_storage.storage [1066]));
 sg13g2_dfrbp_1 \shift_storage.storage[1067]$_SDFFE_PN0P_  (.CLK(clknet_leaf_125_clk_p2c),
    .RESET_B(net673),
    .D(_00177_),
    .Q_N(_06624_),
    .Q(\shift_storage.storage [1067]));
 sg13g2_dfrbp_1 \shift_storage.storage[1068]$_SDFFE_PN0P_  (.CLK(clknet_leaf_125_clk_p2c),
    .RESET_B(net674),
    .D(_00178_),
    .Q_N(_06623_),
    .Q(\shift_storage.storage [1068]));
 sg13g2_dfrbp_1 \shift_storage.storage[1069]$_SDFFE_PN0P_  (.CLK(clknet_leaf_124_clk_p2c),
    .RESET_B(net675),
    .D(_00179_),
    .Q_N(_06622_),
    .Q(\shift_storage.storage [1069]));
 sg13g2_dfrbp_1 \shift_storage.storage[106]$_SDFFE_PN0P_  (.CLK(clknet_leaf_124_clk_p2c),
    .RESET_B(net676),
    .D(_00180_),
    .Q_N(_06621_),
    .Q(\shift_storage.storage [106]));
 sg13g2_dfrbp_1 \shift_storage.storage[1070]$_SDFFE_PN0P_  (.CLK(clknet_leaf_124_clk_p2c),
    .RESET_B(net677),
    .D(_00181_),
    .Q_N(_06620_),
    .Q(\shift_storage.storage [1070]));
 sg13g2_dfrbp_1 \shift_storage.storage[1071]$_SDFFE_PN0P_  (.CLK(clknet_leaf_124_clk_p2c),
    .RESET_B(net678),
    .D(_00182_),
    .Q_N(_06619_),
    .Q(\shift_storage.storage [1071]));
 sg13g2_dfrbp_1 \shift_storage.storage[1072]$_SDFFE_PN0P_  (.CLK(clknet_leaf_124_clk_p2c),
    .RESET_B(net679),
    .D(_00183_),
    .Q_N(_06618_),
    .Q(\shift_storage.storage [1072]));
 sg13g2_dfrbp_1 \shift_storage.storage[1073]$_SDFFE_PN0P_  (.CLK(clknet_leaf_193_clk_p2c),
    .RESET_B(net680),
    .D(_00184_),
    .Q_N(_06617_),
    .Q(\shift_storage.storage [1073]));
 sg13g2_dfrbp_1 \shift_storage.storage[1074]$_SDFFE_PN0P_  (.CLK(clknet_leaf_193_clk_p2c),
    .RESET_B(net681),
    .D(_00185_),
    .Q_N(_06616_),
    .Q(\shift_storage.storage [1074]));
 sg13g2_dfrbp_1 \shift_storage.storage[1075]$_SDFFE_PN0P_  (.CLK(clknet_leaf_124_clk_p2c),
    .RESET_B(net682),
    .D(_00186_),
    .Q_N(_06615_),
    .Q(\shift_storage.storage [1075]));
 sg13g2_dfrbp_1 \shift_storage.storage[1076]$_SDFFE_PN0P_  (.CLK(clknet_leaf_124_clk_p2c),
    .RESET_B(net683),
    .D(_00187_),
    .Q_N(_06614_),
    .Q(\shift_storage.storage [1076]));
 sg13g2_dfrbp_1 \shift_storage.storage[1077]$_SDFFE_PN0P_  (.CLK(clknet_leaf_47_clk_p2c),
    .RESET_B(net684),
    .D(_00188_),
    .Q_N(_06613_),
    .Q(\shift_storage.storage [1077]));
 sg13g2_dfrbp_1 \shift_storage.storage[1078]$_SDFFE_PN0P_  (.CLK(clknet_leaf_47_clk_p2c),
    .RESET_B(net685),
    .D(_00189_),
    .Q_N(_06612_),
    .Q(\shift_storage.storage [1078]));
 sg13g2_dfrbp_1 \shift_storage.storage[1079]$_SDFFE_PN0P_  (.CLK(clknet_leaf_47_clk_p2c),
    .RESET_B(net686),
    .D(_00190_),
    .Q_N(_06611_),
    .Q(\shift_storage.storage [1079]));
 sg13g2_dfrbp_1 \shift_storage.storage[107]$_SDFFE_PN0P_  (.CLK(clknet_leaf_48_clk_p2c),
    .RESET_B(net687),
    .D(_00191_),
    .Q_N(_06610_),
    .Q(\shift_storage.storage [107]));
 sg13g2_dfrbp_1 \shift_storage.storage[1080]$_SDFFE_PN0P_  (.CLK(clknet_leaf_245_clk_p2c),
    .RESET_B(net688),
    .D(_00192_),
    .Q_N(_06609_),
    .Q(\shift_storage.storage [1080]));
 sg13g2_dfrbp_1 \shift_storage.storage[1081]$_SDFFE_PN0P_  (.CLK(clknet_leaf_47_clk_p2c),
    .RESET_B(net689),
    .D(_00193_),
    .Q_N(_06608_),
    .Q(\shift_storage.storage [1081]));
 sg13g2_dfrbp_1 \shift_storage.storage[1082]$_SDFFE_PN0P_  (.CLK(clknet_leaf_47_clk_p2c),
    .RESET_B(net690),
    .D(_00194_),
    .Q_N(_06607_),
    .Q(\shift_storage.storage [1082]));
 sg13g2_dfrbp_1 \shift_storage.storage[1083]$_SDFFE_PN0P_  (.CLK(clknet_leaf_48_clk_p2c),
    .RESET_B(net691),
    .D(_00195_),
    .Q_N(_06606_),
    .Q(\shift_storage.storage [1083]));
 sg13g2_dfrbp_1 \shift_storage.storage[1084]$_SDFFE_PN0P_  (.CLK(clknet_leaf_48_clk_p2c),
    .RESET_B(net692),
    .D(_00196_),
    .Q_N(_06605_),
    .Q(\shift_storage.storage [1084]));
 sg13g2_dfrbp_1 \shift_storage.storage[1085]$_SDFFE_PN0P_  (.CLK(clknet_leaf_46_clk_p2c),
    .RESET_B(net693),
    .D(_00197_),
    .Q_N(_06604_),
    .Q(\shift_storage.storage [1085]));
 sg13g2_dfrbp_1 \shift_storage.storage[1086]$_SDFFE_PN0P_  (.CLK(clknet_leaf_46_clk_p2c),
    .RESET_B(net694),
    .D(_00198_),
    .Q_N(_06603_),
    .Q(\shift_storage.storage [1086]));
 sg13g2_dfrbp_1 \shift_storage.storage[1087]$_SDFFE_PN0P_  (.CLK(clknet_leaf_46_clk_p2c),
    .RESET_B(net695),
    .D(_00199_),
    .Q_N(_06602_),
    .Q(\shift_storage.storage [1087]));
 sg13g2_dfrbp_1 \shift_storage.storage[1088]$_SDFFE_PN0P_  (.CLK(clknet_leaf_47_clk_p2c),
    .RESET_B(net696),
    .D(_00200_),
    .Q_N(_06601_),
    .Q(\shift_storage.storage [1088]));
 sg13g2_dfrbp_1 \shift_storage.storage[1089]$_SDFFE_PN0P_  (.CLK(clknet_leaf_246_clk_p2c),
    .RESET_B(net697),
    .D(_00201_),
    .Q_N(_06600_),
    .Q(\shift_storage.storage [1089]));
 sg13g2_dfrbp_1 \shift_storage.storage[108]$_SDFFE_PN0P_  (.CLK(clknet_leaf_246_clk_p2c),
    .RESET_B(net698),
    .D(_00202_),
    .Q_N(_06599_),
    .Q(\shift_storage.storage [108]));
 sg13g2_dfrbp_1 \shift_storage.storage[1090]$_SDFFE_PN0P_  (.CLK(clknet_leaf_246_clk_p2c),
    .RESET_B(net699),
    .D(_00203_),
    .Q_N(_06598_),
    .Q(\shift_storage.storage [1090]));
 sg13g2_dfrbp_1 \shift_storage.storage[1091]$_SDFFE_PN0P_  (.CLK(clknet_leaf_247_clk_p2c),
    .RESET_B(net700),
    .D(_00204_),
    .Q_N(_06597_),
    .Q(\shift_storage.storage [1091]));
 sg13g2_dfrbp_1 \shift_storage.storage[1092]$_SDFFE_PN0P_  (.CLK(clknet_leaf_248_clk_p2c),
    .RESET_B(net701),
    .D(_00205_),
    .Q_N(_06596_),
    .Q(\shift_storage.storage [1092]));
 sg13g2_dfrbp_1 \shift_storage.storage[1093]$_SDFFE_PN0P_  (.CLK(clknet_leaf_247_clk_p2c),
    .RESET_B(net702),
    .D(_00206_),
    .Q_N(_06595_),
    .Q(\shift_storage.storage [1093]));
 sg13g2_dfrbp_1 \shift_storage.storage[1094]$_SDFFE_PN0P_  (.CLK(clknet_leaf_247_clk_p2c),
    .RESET_B(net703),
    .D(_00207_),
    .Q_N(_06594_),
    .Q(\shift_storage.storage [1094]));
 sg13g2_dfrbp_1 \shift_storage.storage[1095]$_SDFFE_PN0P_  (.CLK(clknet_leaf_246_clk_p2c),
    .RESET_B(net704),
    .D(_00208_),
    .Q_N(_06593_),
    .Q(\shift_storage.storage [1095]));
 sg13g2_dfrbp_1 \shift_storage.storage[1096]$_SDFFE_PN0P_  (.CLK(clknet_leaf_244_clk_p2c),
    .RESET_B(net705),
    .D(_00209_),
    .Q_N(_06592_),
    .Q(\shift_storage.storage [1096]));
 sg13g2_dfrbp_1 \shift_storage.storage[1097]$_SDFFE_PN0P_  (.CLK(clknet_leaf_244_clk_p2c),
    .RESET_B(net706),
    .D(_00210_),
    .Q_N(_06591_),
    .Q(\shift_storage.storage [1097]));
 sg13g2_dfrbp_1 \shift_storage.storage[1098]$_SDFFE_PN0P_  (.CLK(clknet_leaf_244_clk_p2c),
    .RESET_B(net707),
    .D(_00211_),
    .Q_N(_06590_),
    .Q(\shift_storage.storage [1098]));
 sg13g2_dfrbp_1 \shift_storage.storage[1099]$_SDFFE_PN0P_  (.CLK(clknet_leaf_246_clk_p2c),
    .RESET_B(net708),
    .D(_00212_),
    .Q_N(_06589_),
    .Q(\shift_storage.storage [1099]));
 sg13g2_dfrbp_1 \shift_storage.storage[109]$_SDFFE_PN0P_  (.CLK(clknet_leaf_245_clk_p2c),
    .RESET_B(net709),
    .D(_00213_),
    .Q_N(_06588_),
    .Q(\shift_storage.storage [109]));
 sg13g2_dfrbp_1 \shift_storage.storage[10]$_SDFFE_PN0P_  (.CLK(clknet_leaf_244_clk_p2c),
    .RESET_B(net710),
    .D(_00214_),
    .Q_N(_06587_),
    .Q(\shift_storage.storage [10]));
 sg13g2_dfrbp_1 \shift_storage.storage[1100]$_SDFFE_PN0P_  (.CLK(clknet_leaf_246_clk_p2c),
    .RESET_B(net711),
    .D(_00215_),
    .Q_N(_06586_),
    .Q(\shift_storage.storage [1100]));
 sg13g2_dfrbp_1 \shift_storage.storage[1101]$_SDFFE_PN0P_  (.CLK(clknet_leaf_245_clk_p2c),
    .RESET_B(net712),
    .D(_00216_),
    .Q_N(_06585_),
    .Q(\shift_storage.storage [1101]));
 sg13g2_dfrbp_1 \shift_storage.storage[1102]$_SDFFE_PN0P_  (.CLK(clknet_leaf_245_clk_p2c),
    .RESET_B(net713),
    .D(_00217_),
    .Q_N(_06584_),
    .Q(\shift_storage.storage [1102]));
 sg13g2_dfrbp_1 \shift_storage.storage[1103]$_SDFFE_PN0P_  (.CLK(clknet_leaf_245_clk_p2c),
    .RESET_B(net714),
    .D(_00218_),
    .Q_N(_06583_),
    .Q(\shift_storage.storage [1103]));
 sg13g2_dfrbp_1 \shift_storage.storage[1104]$_SDFFE_PN0P_  (.CLK(clknet_leaf_245_clk_p2c),
    .RESET_B(net715),
    .D(_00219_),
    .Q_N(_06582_),
    .Q(\shift_storage.storage [1104]));
 sg13g2_dfrbp_1 \shift_storage.storage[1105]$_SDFFE_PN0P_  (.CLK(clknet_leaf_194_clk_p2c),
    .RESET_B(net716),
    .D(_00220_),
    .Q_N(_06581_),
    .Q(\shift_storage.storage [1105]));
 sg13g2_dfrbp_1 \shift_storage.storage[1106]$_SDFFE_PN0P_  (.CLK(clknet_leaf_194_clk_p2c),
    .RESET_B(net717),
    .D(_00221_),
    .Q_N(_06580_),
    .Q(\shift_storage.storage [1106]));
 sg13g2_dfrbp_1 \shift_storage.storage[1107]$_SDFFE_PN0P_  (.CLK(clknet_leaf_195_clk_p2c),
    .RESET_B(net718),
    .D(_00222_),
    .Q_N(_06579_),
    .Q(\shift_storage.storage [1107]));
 sg13g2_dfrbp_1 \shift_storage.storage[1108]$_SDFFE_PN0P_  (.CLK(clknet_leaf_195_clk_p2c),
    .RESET_B(net719),
    .D(_00223_),
    .Q_N(_06578_),
    .Q(\shift_storage.storage [1108]));
 sg13g2_dfrbp_1 \shift_storage.storage[1109]$_SDFFE_PN0P_  (.CLK(clknet_leaf_195_clk_p2c),
    .RESET_B(net720),
    .D(_00224_),
    .Q_N(_06577_),
    .Q(\shift_storage.storage [1109]));
 sg13g2_dfrbp_1 \shift_storage.storage[110]$_SDFFE_PN0P_  (.CLK(clknet_leaf_243_clk_p2c),
    .RESET_B(net721),
    .D(_00225_),
    .Q_N(_06576_),
    .Q(\shift_storage.storage [110]));
 sg13g2_dfrbp_1 \shift_storage.storage[1110]$_SDFFE_PN0P_  (.CLK(clknet_leaf_195_clk_p2c),
    .RESET_B(net722),
    .D(_00226_),
    .Q_N(_06575_),
    .Q(\shift_storage.storage [1110]));
 sg13g2_dfrbp_1 \shift_storage.storage[1111]$_SDFFE_PN0P_  (.CLK(clknet_leaf_243_clk_p2c),
    .RESET_B(net723),
    .D(_00227_),
    .Q_N(_06574_),
    .Q(\shift_storage.storage [1111]));
 sg13g2_dfrbp_1 \shift_storage.storage[1112]$_SDFFE_PN0P_  (.CLK(clknet_leaf_243_clk_p2c),
    .RESET_B(net724),
    .D(_00228_),
    .Q_N(_06573_),
    .Q(\shift_storage.storage [1112]));
 sg13g2_dfrbp_1 \shift_storage.storage[1113]$_SDFFE_PN0P_  (.CLK(clknet_leaf_243_clk_p2c),
    .RESET_B(net725),
    .D(_00229_),
    .Q_N(_06572_),
    .Q(\shift_storage.storage [1113]));
 sg13g2_dfrbp_1 \shift_storage.storage[1114]$_SDFFE_PN0P_  (.CLK(clknet_leaf_242_clk_p2c),
    .RESET_B(net726),
    .D(_00230_),
    .Q_N(_06571_),
    .Q(\shift_storage.storage [1114]));
 sg13g2_dfrbp_1 \shift_storage.storage[1115]$_SDFFE_PN0P_  (.CLK(clknet_leaf_243_clk_p2c),
    .RESET_B(net727),
    .D(_00231_),
    .Q_N(_06570_),
    .Q(\shift_storage.storage [1115]));
 sg13g2_dfrbp_1 \shift_storage.storage[1116]$_SDFFE_PN0P_  (.CLK(clknet_leaf_243_clk_p2c),
    .RESET_B(net728),
    .D(_00232_),
    .Q_N(_06569_),
    .Q(\shift_storage.storage [1116]));
 sg13g2_dfrbp_1 \shift_storage.storage[1117]$_SDFFE_PN0P_  (.CLK(clknet_leaf_241_clk_p2c),
    .RESET_B(net729),
    .D(_00233_),
    .Q_N(_06568_),
    .Q(\shift_storage.storage [1117]));
 sg13g2_dfrbp_1 \shift_storage.storage[1118]$_SDFFE_PN0P_  (.CLK(clknet_leaf_241_clk_p2c),
    .RESET_B(net730),
    .D(_00234_),
    .Q_N(_06567_),
    .Q(\shift_storage.storage [1118]));
 sg13g2_dfrbp_1 \shift_storage.storage[1119]$_SDFFE_PN0P_  (.CLK(clknet_leaf_242_clk_p2c),
    .RESET_B(net731),
    .D(_00235_),
    .Q_N(_06566_),
    .Q(\shift_storage.storage [1119]));
 sg13g2_dfrbp_1 \shift_storage.storage[111]$_SDFFE_PN0P_  (.CLK(clknet_leaf_244_clk_p2c),
    .RESET_B(net732),
    .D(_00236_),
    .Q_N(_06565_),
    .Q(\shift_storage.storage [111]));
 sg13g2_dfrbp_1 \shift_storage.storage[1120]$_SDFFE_PN0P_  (.CLK(clknet_leaf_242_clk_p2c),
    .RESET_B(net733),
    .D(_00237_),
    .Q_N(_06564_),
    .Q(\shift_storage.storage [1120]));
 sg13g2_dfrbp_1 \shift_storage.storage[1121]$_SDFFE_PN0P_  (.CLK(clknet_leaf_242_clk_p2c),
    .RESET_B(net734),
    .D(_00238_),
    .Q_N(_06563_),
    .Q(\shift_storage.storage [1121]));
 sg13g2_dfrbp_1 \shift_storage.storage[1122]$_SDFFE_PN0P_  (.CLK(clknet_leaf_241_clk_p2c),
    .RESET_B(net735),
    .D(_00239_),
    .Q_N(_06562_),
    .Q(\shift_storage.storage [1122]));
 sg13g2_dfrbp_1 \shift_storage.storage[1123]$_SDFFE_PN0P_  (.CLK(clknet_leaf_236_clk_p2c),
    .RESET_B(net736),
    .D(_00240_),
    .Q_N(_06561_),
    .Q(\shift_storage.storage [1123]));
 sg13g2_dfrbp_1 \shift_storage.storage[1124]$_SDFFE_PN0P_  (.CLK(clknet_leaf_240_clk_p2c),
    .RESET_B(net737),
    .D(_00241_),
    .Q_N(_06560_),
    .Q(\shift_storage.storage [1124]));
 sg13g2_dfrbp_1 \shift_storage.storage[1125]$_SDFFE_PN0P_  (.CLK(clknet_leaf_241_clk_p2c),
    .RESET_B(net738),
    .D(_00242_),
    .Q_N(_06559_),
    .Q(\shift_storage.storage [1125]));
 sg13g2_dfrbp_1 \shift_storage.storage[1126]$_SDFFE_PN0P_  (.CLK(clknet_leaf_241_clk_p2c),
    .RESET_B(net739),
    .D(_00243_),
    .Q_N(_06558_),
    .Q(\shift_storage.storage [1126]));
 sg13g2_dfrbp_1 \shift_storage.storage[1127]$_SDFFE_PN0P_  (.CLK(clknet_leaf_240_clk_p2c),
    .RESET_B(net740),
    .D(_00244_),
    .Q_N(_06557_),
    .Q(\shift_storage.storage [1127]));
 sg13g2_dfrbp_1 \shift_storage.storage[1128]$_SDFFE_PN0P_  (.CLK(clknet_leaf_240_clk_p2c),
    .RESET_B(net741),
    .D(_00245_),
    .Q_N(_06556_),
    .Q(\shift_storage.storage [1128]));
 sg13g2_dfrbp_1 \shift_storage.storage[1129]$_SDFFE_PN0P_  (.CLK(clknet_leaf_250_clk_p2c),
    .RESET_B(net742),
    .D(_00246_),
    .Q_N(_06555_),
    .Q(\shift_storage.storage [1129]));
 sg13g2_dfrbp_1 \shift_storage.storage[112]$_SDFFE_PN0P_  (.CLK(clknet_leaf_241_clk_p2c),
    .RESET_B(net743),
    .D(_00247_),
    .Q_N(_06554_),
    .Q(\shift_storage.storage [112]));
 sg13g2_dfrbp_1 \shift_storage.storage[1130]$_SDFFE_PN0P_  (.CLK(clknet_leaf_240_clk_p2c),
    .RESET_B(net744),
    .D(_00248_),
    .Q_N(_06553_),
    .Q(\shift_storage.storage [1130]));
 sg13g2_dfrbp_1 \shift_storage.storage[1131]$_SDFFE_PN0P_  (.CLK(clknet_leaf_240_clk_p2c),
    .RESET_B(net745),
    .D(_00249_),
    .Q_N(_06552_),
    .Q(\shift_storage.storage [1131]));
 sg13g2_dfrbp_1 \shift_storage.storage[1132]$_SDFFE_PN0P_  (.CLK(clknet_leaf_240_clk_p2c),
    .RESET_B(net746),
    .D(_00250_),
    .Q_N(_06551_),
    .Q(\shift_storage.storage [1132]));
 sg13g2_dfrbp_1 \shift_storage.storage[1133]$_SDFFE_PN0P_  (.CLK(clknet_leaf_244_clk_p2c),
    .RESET_B(net747),
    .D(_00251_),
    .Q_N(_06550_),
    .Q(\shift_storage.storage [1133]));
 sg13g2_dfrbp_1 \shift_storage.storage[1134]$_SDFFE_PN0P_  (.CLK(clknet_leaf_247_clk_p2c),
    .RESET_B(net748),
    .D(_00252_),
    .Q_N(_06549_),
    .Q(\shift_storage.storage [1134]));
 sg13g2_dfrbp_1 \shift_storage.storage[1135]$_SDFFE_PN0P_  (.CLK(clknet_leaf_247_clk_p2c),
    .RESET_B(net749),
    .D(_00253_),
    .Q_N(_06548_),
    .Q(\shift_storage.storage [1135]));
 sg13g2_dfrbp_1 \shift_storage.storage[1136]$_SDFFE_PN0P_  (.CLK(clknet_leaf_249_clk_p2c),
    .RESET_B(net750),
    .D(_00254_),
    .Q_N(_06547_),
    .Q(\shift_storage.storage [1136]));
 sg13g2_dfrbp_1 \shift_storage.storage[1137]$_SDFFE_PN0P_  (.CLK(clknet_leaf_249_clk_p2c),
    .RESET_B(net751),
    .D(_00255_),
    .Q_N(_06546_),
    .Q(\shift_storage.storage [1137]));
 sg13g2_dfrbp_1 \shift_storage.storage[1138]$_SDFFE_PN0P_  (.CLK(clknet_leaf_248_clk_p2c),
    .RESET_B(net752),
    .D(_00256_),
    .Q_N(_06545_),
    .Q(\shift_storage.storage [1138]));
 sg13g2_dfrbp_1 \shift_storage.storage[1139]$_SDFFE_PN0P_  (.CLK(clknet_leaf_247_clk_p2c),
    .RESET_B(net753),
    .D(_00257_),
    .Q_N(_06544_),
    .Q(\shift_storage.storage [1139]));
 sg13g2_dfrbp_1 \shift_storage.storage[113]$_SDFFE_PN0P_  (.CLK(clknet_leaf_249_clk_p2c),
    .RESET_B(net754),
    .D(_00258_),
    .Q_N(_06543_),
    .Q(\shift_storage.storage [113]));
 sg13g2_dfrbp_1 \shift_storage.storage[1140]$_SDFFE_PN0P_  (.CLK(clknet_leaf_248_clk_p2c),
    .RESET_B(net755),
    .D(_00259_),
    .Q_N(_06542_),
    .Q(\shift_storage.storage [1140]));
 sg13g2_dfrbp_1 \shift_storage.storage[1141]$_SDFFE_PN0P_  (.CLK(clknet_leaf_248_clk_p2c),
    .RESET_B(net756),
    .D(_00260_),
    .Q_N(_06541_),
    .Q(\shift_storage.storage [1141]));
 sg13g2_dfrbp_1 \shift_storage.storage[1142]$_SDFFE_PN0P_  (.CLK(clknet_leaf_248_clk_p2c),
    .RESET_B(net757),
    .D(_00261_),
    .Q_N(_06540_),
    .Q(\shift_storage.storage [1142]));
 sg13g2_dfrbp_1 \shift_storage.storage[1143]$_SDFFE_PN0P_  (.CLK(clknet_leaf_248_clk_p2c),
    .RESET_B(net758),
    .D(_00262_),
    .Q_N(_06539_),
    .Q(\shift_storage.storage [1143]));
 sg13g2_dfrbp_1 \shift_storage.storage[1144]$_SDFFE_PN0P_  (.CLK(clknet_leaf_253_clk_p2c),
    .RESET_B(net759),
    .D(_00263_),
    .Q_N(_06538_),
    .Q(\shift_storage.storage [1144]));
 sg13g2_dfrbp_1 \shift_storage.storage[1145]$_SDFFE_PN0P_  (.CLK(clknet_leaf_253_clk_p2c),
    .RESET_B(net760),
    .D(_00264_),
    .Q_N(_06537_),
    .Q(\shift_storage.storage [1145]));
 sg13g2_dfrbp_1 \shift_storage.storage[1146]$_SDFFE_PN0P_  (.CLK(clknet_leaf_249_clk_p2c),
    .RESET_B(net761),
    .D(_00265_),
    .Q_N(_06536_),
    .Q(\shift_storage.storage [1146]));
 sg13g2_dfrbp_1 \shift_storage.storage[1147]$_SDFFE_PN0P_  (.CLK(clknet_leaf_249_clk_p2c),
    .RESET_B(net762),
    .D(_00266_),
    .Q_N(_06535_),
    .Q(\shift_storage.storage [1147]));
 sg13g2_dfrbp_1 \shift_storage.storage[1148]$_SDFFE_PN0P_  (.CLK(clknet_leaf_249_clk_p2c),
    .RESET_B(net763),
    .D(_00267_),
    .Q_N(_06534_),
    .Q(\shift_storage.storage [1148]));
 sg13g2_dfrbp_1 \shift_storage.storage[1149]$_SDFFE_PN0P_  (.CLK(clknet_leaf_250_clk_p2c),
    .RESET_B(net764),
    .D(_00268_),
    .Q_N(_06533_),
    .Q(\shift_storage.storage [1149]));
 sg13g2_dfrbp_1 \shift_storage.storage[114]$_SDFFE_PN0P_  (.CLK(clknet_leaf_250_clk_p2c),
    .RESET_B(net765),
    .D(_00269_),
    .Q_N(_06532_),
    .Q(\shift_storage.storage [114]));
 sg13g2_dfrbp_1 \shift_storage.storage[1150]$_SDFFE_PN0P_  (.CLK(clknet_leaf_250_clk_p2c),
    .RESET_B(net766),
    .D(_00270_),
    .Q_N(_06531_),
    .Q(\shift_storage.storage [1150]));
 sg13g2_dfrbp_1 \shift_storage.storage[1151]$_SDFFE_PN0P_  (.CLK(clknet_leaf_250_clk_p2c),
    .RESET_B(net767),
    .D(_00271_),
    .Q_N(_06530_),
    .Q(\shift_storage.storage [1151]));
 sg13g2_dfrbp_1 \shift_storage.storage[1152]$_SDFFE_PN0P_  (.CLK(clknet_leaf_253_clk_p2c),
    .RESET_B(net768),
    .D(_00272_),
    .Q_N(_06529_),
    .Q(\shift_storage.storage [1152]));
 sg13g2_dfrbp_1 \shift_storage.storage[1153]$_SDFFE_PN0P_  (.CLK(clknet_leaf_253_clk_p2c),
    .RESET_B(net769),
    .D(_00273_),
    .Q_N(_06528_),
    .Q(\shift_storage.storage [1153]));
 sg13g2_dfrbp_1 \shift_storage.storage[1154]$_SDFFE_PN0P_  (.CLK(clknet_leaf_252_clk_p2c),
    .RESET_B(net770),
    .D(_00274_),
    .Q_N(_06527_),
    .Q(\shift_storage.storage [1154]));
 sg13g2_dfrbp_1 \shift_storage.storage[1155]$_SDFFE_PN0P_  (.CLK(clknet_leaf_252_clk_p2c),
    .RESET_B(net771),
    .D(_00275_),
    .Q_N(_06526_),
    .Q(\shift_storage.storage [1155]));
 sg13g2_dfrbp_1 \shift_storage.storage[1156]$_SDFFE_PN0P_  (.CLK(clknet_leaf_251_clk_p2c),
    .RESET_B(net772),
    .D(_00276_),
    .Q_N(_06525_),
    .Q(\shift_storage.storage [1156]));
 sg13g2_dfrbp_1 \shift_storage.storage[1157]$_SDFFE_PN0P_  (.CLK(clknet_leaf_251_clk_p2c),
    .RESET_B(net773),
    .D(_00277_),
    .Q_N(_06524_),
    .Q(\shift_storage.storage [1157]));
 sg13g2_dfrbp_1 \shift_storage.storage[1158]$_SDFFE_PN0P_  (.CLK(clknet_leaf_251_clk_p2c),
    .RESET_B(net774),
    .D(_00278_),
    .Q_N(_06523_),
    .Q(\shift_storage.storage [1158]));
 sg13g2_dfrbp_1 \shift_storage.storage[1159]$_SDFFE_PN0P_  (.CLK(clknet_leaf_251_clk_p2c),
    .RESET_B(net775),
    .D(_00279_),
    .Q_N(_06522_),
    .Q(\shift_storage.storage [1159]));
 sg13g2_dfrbp_1 \shift_storage.storage[115]$_SDFFE_PN0P_  (.CLK(clknet_leaf_239_clk_p2c),
    .RESET_B(net776),
    .D(_00280_),
    .Q_N(_06521_),
    .Q(\shift_storage.storage [115]));
 sg13g2_dfrbp_1 \shift_storage.storage[1160]$_SDFFE_PN0P_  (.CLK(clknet_leaf_251_clk_p2c),
    .RESET_B(net777),
    .D(_00281_),
    .Q_N(_06520_),
    .Q(\shift_storage.storage [1160]));
 sg13g2_dfrbp_1 \shift_storage.storage[1161]$_SDFFE_PN0P_  (.CLK(clknet_leaf_239_clk_p2c),
    .RESET_B(net778),
    .D(_00282_),
    .Q_N(_06519_),
    .Q(\shift_storage.storage [1161]));
 sg13g2_dfrbp_1 \shift_storage.storage[1162]$_SDFFE_PN0P_  (.CLK(clknet_leaf_239_clk_p2c),
    .RESET_B(net779),
    .D(_00283_),
    .Q_N(_06518_),
    .Q(\shift_storage.storage [1162]));
 sg13g2_dfrbp_1 \shift_storage.storage[1163]$_SDFFE_PN0P_  (.CLK(clknet_leaf_239_clk_p2c),
    .RESET_B(net780),
    .D(_00284_),
    .Q_N(_06517_),
    .Q(\shift_storage.storage [1163]));
 sg13g2_dfrbp_1 \shift_storage.storage[1164]$_SDFFE_PN0P_  (.CLK(clknet_leaf_239_clk_p2c),
    .RESET_B(net781),
    .D(_00285_),
    .Q_N(_06516_),
    .Q(\shift_storage.storage [1164]));
 sg13g2_dfrbp_1 \shift_storage.storage[1165]$_SDFFE_PN0P_  (.CLK(clknet_leaf_239_clk_p2c),
    .RESET_B(net782),
    .D(_00286_),
    .Q_N(_06515_),
    .Q(\shift_storage.storage [1165]));
 sg13g2_dfrbp_1 \shift_storage.storage[1166]$_SDFFE_PN0P_  (.CLK(clknet_leaf_228_clk_p2c),
    .RESET_B(net783),
    .D(_00287_),
    .Q_N(_06514_),
    .Q(\shift_storage.storage [1166]));
 sg13g2_dfrbp_1 \shift_storage.storage[1167]$_SDFFE_PN0P_  (.CLK(clknet_leaf_238_clk_p2c),
    .RESET_B(net784),
    .D(_00288_),
    .Q_N(_06513_),
    .Q(\shift_storage.storage [1167]));
 sg13g2_dfrbp_1 \shift_storage.storage[1168]$_SDFFE_PN0P_  (.CLK(clknet_leaf_238_clk_p2c),
    .RESET_B(net785),
    .D(_00289_),
    .Q_N(_06512_),
    .Q(\shift_storage.storage [1168]));
 sg13g2_dfrbp_1 \shift_storage.storage[1169]$_SDFFE_PN0P_  (.CLK(clknet_leaf_238_clk_p2c),
    .RESET_B(net786),
    .D(_00290_),
    .Q_N(_06511_),
    .Q(\shift_storage.storage [1169]));
 sg13g2_dfrbp_1 \shift_storage.storage[116]$_SDFFE_PN0P_  (.CLK(clknet_leaf_238_clk_p2c),
    .RESET_B(net787),
    .D(_00291_),
    .Q_N(_06510_),
    .Q(\shift_storage.storage [116]));
 sg13g2_dfrbp_1 \shift_storage.storage[1170]$_SDFFE_PN0P_  (.CLK(clknet_leaf_238_clk_p2c),
    .RESET_B(net788),
    .D(_00292_),
    .Q_N(_06509_),
    .Q(\shift_storage.storage [1170]));
 sg13g2_dfrbp_1 \shift_storage.storage[1171]$_SDFFE_PN0P_  (.CLK(clknet_leaf_238_clk_p2c),
    .RESET_B(net789),
    .D(_00293_),
    .Q_N(_06508_),
    .Q(\shift_storage.storage [1171]));
 sg13g2_dfrbp_1 \shift_storage.storage[1172]$_SDFFE_PN0P_  (.CLK(clknet_leaf_237_clk_p2c),
    .RESET_B(net790),
    .D(_00294_),
    .Q_N(_06507_),
    .Q(\shift_storage.storage [1172]));
 sg13g2_dfrbp_1 \shift_storage.storage[1173]$_SDFFE_PN0P_  (.CLK(clknet_leaf_237_clk_p2c),
    .RESET_B(net791),
    .D(_00295_),
    .Q_N(_06506_),
    .Q(\shift_storage.storage [1173]));
 sg13g2_dfrbp_1 \shift_storage.storage[1174]$_SDFFE_PN0P_  (.CLK(clknet_leaf_229_clk_p2c),
    .RESET_B(net792),
    .D(_00296_),
    .Q_N(_06505_),
    .Q(\shift_storage.storage [1174]));
 sg13g2_dfrbp_1 \shift_storage.storage[1175]$_SDFFE_PN0P_  (.CLK(clknet_leaf_228_clk_p2c),
    .RESET_B(net793),
    .D(_00297_),
    .Q_N(_06504_),
    .Q(\shift_storage.storage [1175]));
 sg13g2_dfrbp_1 \shift_storage.storage[1176]$_SDFFE_PN0P_  (.CLK(clknet_leaf_229_clk_p2c),
    .RESET_B(net794),
    .D(_00298_),
    .Q_N(_06503_),
    .Q(\shift_storage.storage [1176]));
 sg13g2_dfrbp_1 \shift_storage.storage[1177]$_SDFFE_PN0P_  (.CLK(clknet_leaf_229_clk_p2c),
    .RESET_B(net795),
    .D(_00299_),
    .Q_N(_06502_),
    .Q(\shift_storage.storage [1177]));
 sg13g2_dfrbp_1 \shift_storage.storage[1178]$_SDFFE_PN0P_  (.CLK(clknet_leaf_229_clk_p2c),
    .RESET_B(net796),
    .D(_00300_),
    .Q_N(_06501_),
    .Q(\shift_storage.storage [1178]));
 sg13g2_dfrbp_1 \shift_storage.storage[1179]$_SDFFE_PN0P_  (.CLK(clknet_leaf_229_clk_p2c),
    .RESET_B(net797),
    .D(_00301_),
    .Q_N(_06500_),
    .Q(\shift_storage.storage [1179]));
 sg13g2_dfrbp_1 \shift_storage.storage[117]$_SDFFE_PN0P_  (.CLK(clknet_leaf_236_clk_p2c),
    .RESET_B(net798),
    .D(_00302_),
    .Q_N(_06499_),
    .Q(\shift_storage.storage [117]));
 sg13g2_dfrbp_1 \shift_storage.storage[1180]$_SDFFE_PN0P_  (.CLK(clknet_leaf_231_clk_p2c),
    .RESET_B(net799),
    .D(_00303_),
    .Q_N(_06498_),
    .Q(\shift_storage.storage [1180]));
 sg13g2_dfrbp_1 \shift_storage.storage[1181]$_SDFFE_PN0P_  (.CLK(clknet_leaf_231_clk_p2c),
    .RESET_B(net800),
    .D(_00304_),
    .Q_N(_06497_),
    .Q(\shift_storage.storage [1181]));
 sg13g2_dfrbp_1 \shift_storage.storage[1182]$_SDFFE_PN0P_  (.CLK(clknet_leaf_234_clk_p2c),
    .RESET_B(net801),
    .D(_00305_),
    .Q_N(_06496_),
    .Q(\shift_storage.storage [1182]));
 sg13g2_dfrbp_1 \shift_storage.storage[1183]$_SDFFE_PN0P_  (.CLK(clknet_leaf_237_clk_p2c),
    .RESET_B(net802),
    .D(_00306_),
    .Q_N(_06495_),
    .Q(\shift_storage.storage [1183]));
 sg13g2_dfrbp_1 \shift_storage.storage[1184]$_SDFFE_PN0P_  (.CLK(clknet_leaf_237_clk_p2c),
    .RESET_B(net803),
    .D(_00307_),
    .Q_N(_06494_),
    .Q(\shift_storage.storage [1184]));
 sg13g2_dfrbp_1 \shift_storage.storage[1185]$_SDFFE_PN0P_  (.CLK(clknet_leaf_237_clk_p2c),
    .RESET_B(net804),
    .D(_00308_),
    .Q_N(_06493_),
    .Q(\shift_storage.storage [1185]));
 sg13g2_dfrbp_1 \shift_storage.storage[1186]$_SDFFE_PN0P_  (.CLK(clknet_leaf_237_clk_p2c),
    .RESET_B(net805),
    .D(_00309_),
    .Q_N(_06492_),
    .Q(\shift_storage.storage [1186]));
 sg13g2_dfrbp_1 \shift_storage.storage[1187]$_SDFFE_PN0P_  (.CLK(clknet_leaf_234_clk_p2c),
    .RESET_B(net806),
    .D(_00310_),
    .Q_N(_06491_),
    .Q(\shift_storage.storage [1187]));
 sg13g2_dfrbp_1 \shift_storage.storage[1188]$_SDFFE_PN0P_  (.CLK(clknet_leaf_234_clk_p2c),
    .RESET_B(net807),
    .D(_00311_),
    .Q_N(_06490_),
    .Q(\shift_storage.storage [1188]));
 sg13g2_dfrbp_1 \shift_storage.storage[1189]$_SDFFE_PN0P_  (.CLK(clknet_leaf_234_clk_p2c),
    .RESET_B(net808),
    .D(_00312_),
    .Q_N(_06489_),
    .Q(\shift_storage.storage [1189]));
 sg13g2_dfrbp_1 \shift_storage.storage[118]$_SDFFE_PN0P_  (.CLK(clknet_leaf_235_clk_p2c),
    .RESET_B(net809),
    .D(_00313_),
    .Q_N(_06488_),
    .Q(\shift_storage.storage [118]));
 sg13g2_dfrbp_1 \shift_storage.storage[1190]$_SDFFE_PN0P_  (.CLK(clknet_leaf_235_clk_p2c),
    .RESET_B(net810),
    .D(_00314_),
    .Q_N(_06487_),
    .Q(\shift_storage.storage [1190]));
 sg13g2_dfrbp_1 \shift_storage.storage[1191]$_SDFFE_PN0P_  (.CLK(clknet_leaf_234_clk_p2c),
    .RESET_B(net811),
    .D(_00315_),
    .Q_N(_06486_),
    .Q(\shift_storage.storage [1191]));
 sg13g2_dfrbp_1 \shift_storage.storage[1192]$_SDFFE_PN0P_  (.CLK(clknet_leaf_236_clk_p2c),
    .RESET_B(net812),
    .D(_00316_),
    .Q_N(_06485_),
    .Q(\shift_storage.storage [1192]));
 sg13g2_dfrbp_1 \shift_storage.storage[1193]$_SDFFE_PN0P_  (.CLK(clknet_leaf_236_clk_p2c),
    .RESET_B(net813),
    .D(_00317_),
    .Q_N(_06484_),
    .Q(\shift_storage.storage [1193]));
 sg13g2_dfrbp_1 \shift_storage.storage[1194]$_SDFFE_PN0P_  (.CLK(clknet_leaf_236_clk_p2c),
    .RESET_B(net814),
    .D(_00318_),
    .Q_N(_06483_),
    .Q(\shift_storage.storage [1194]));
 sg13g2_dfrbp_1 \shift_storage.storage[1195]$_SDFFE_PN0P_  (.CLK(clknet_leaf_242_clk_p2c),
    .RESET_B(net815),
    .D(_00319_),
    .Q_N(_06482_),
    .Q(\shift_storage.storage [1195]));
 sg13g2_dfrbp_1 \shift_storage.storage[1196]$_SDFFE_PN0P_  (.CLK(clknet_leaf_235_clk_p2c),
    .RESET_B(net816),
    .D(_00320_),
    .Q_N(_06481_),
    .Q(\shift_storage.storage [1196]));
 sg13g2_dfrbp_1 \shift_storage.storage[1197]$_SDFFE_PN0P_  (.CLK(clknet_leaf_201_clk_p2c),
    .RESET_B(net817),
    .D(_00321_),
    .Q_N(_06480_),
    .Q(\shift_storage.storage [1197]));
 sg13g2_dfrbp_1 \shift_storage.storage[1198]$_SDFFE_PN0P_  (.CLK(clknet_leaf_201_clk_p2c),
    .RESET_B(net818),
    .D(_00322_),
    .Q_N(_06479_),
    .Q(\shift_storage.storage [1198]));
 sg13g2_dfrbp_1 \shift_storage.storage[1199]$_SDFFE_PN0P_  (.CLK(clknet_leaf_242_clk_p2c),
    .RESET_B(net819),
    .D(_00323_),
    .Q_N(_06478_),
    .Q(\shift_storage.storage [1199]));
 sg13g2_dfrbp_1 \shift_storage.storage[119]$_SDFFE_PN0P_  (.CLK(clknet_leaf_235_clk_p2c),
    .RESET_B(net820),
    .D(_00324_),
    .Q_N(_06477_),
    .Q(\shift_storage.storage [119]));
 sg13g2_dfrbp_1 \shift_storage.storage[11]$_SDFFE_PN0P_  (.CLK(clknet_leaf_196_clk_p2c),
    .RESET_B(net821),
    .D(_00325_),
    .Q_N(_06476_),
    .Q(\shift_storage.storage [11]));
 sg13g2_dfrbp_1 \shift_storage.storage[1200]$_SDFFE_PN0P_  (.CLK(clknet_leaf_196_clk_p2c),
    .RESET_B(net822),
    .D(_00326_),
    .Q_N(_06475_),
    .Q(\shift_storage.storage [1200]));
 sg13g2_dfrbp_1 \shift_storage.storage[1201]$_SDFFE_PN0P_  (.CLK(clknet_leaf_195_clk_p2c),
    .RESET_B(net823),
    .D(_00327_),
    .Q_N(_06474_),
    .Q(\shift_storage.storage [1201]));
 sg13g2_dfrbp_1 \shift_storage.storage[1202]$_SDFFE_PN0P_  (.CLK(clknet_leaf_196_clk_p2c),
    .RESET_B(net824),
    .D(_00328_),
    .Q_N(_06473_),
    .Q(\shift_storage.storage [1202]));
 sg13g2_dfrbp_1 \shift_storage.storage[1203]$_SDFFE_PN0P_  (.CLK(clknet_leaf_200_clk_p2c),
    .RESET_B(net825),
    .D(_00329_),
    .Q_N(_06472_),
    .Q(\shift_storage.storage [1203]));
 sg13g2_dfrbp_1 \shift_storage.storage[1204]$_SDFFE_PN0P_  (.CLK(clknet_leaf_200_clk_p2c),
    .RESET_B(net826),
    .D(_00330_),
    .Q_N(_06471_),
    .Q(\shift_storage.storage [1204]));
 sg13g2_dfrbp_1 \shift_storage.storage[1205]$_SDFFE_PN0P_  (.CLK(clknet_leaf_201_clk_p2c),
    .RESET_B(net827),
    .D(_00331_),
    .Q_N(_06470_),
    .Q(\shift_storage.storage [1205]));
 sg13g2_dfrbp_1 \shift_storage.storage[1206]$_SDFFE_PN0P_  (.CLK(clknet_leaf_201_clk_p2c),
    .RESET_B(net828),
    .D(_00332_),
    .Q_N(_06469_),
    .Q(\shift_storage.storage [1206]));
 sg13g2_dfrbp_1 \shift_storage.storage[1207]$_SDFFE_PN0P_  (.CLK(clknet_leaf_201_clk_p2c),
    .RESET_B(net829),
    .D(_00333_),
    .Q_N(_06468_),
    .Q(\shift_storage.storage [1207]));
 sg13g2_dfrbp_1 \shift_storage.storage[1208]$_SDFFE_PN0P_  (.CLK(clknet_leaf_202_clk_p2c),
    .RESET_B(net830),
    .D(_00334_),
    .Q_N(_06467_),
    .Q(\shift_storage.storage [1208]));
 sg13g2_dfrbp_1 \shift_storage.storage[1209]$_SDFFE_PN0P_  (.CLK(clknet_leaf_202_clk_p2c),
    .RESET_B(net831),
    .D(_00335_),
    .Q_N(_06466_),
    .Q(\shift_storage.storage [1209]));
 sg13g2_dfrbp_1 \shift_storage.storage[120]$_SDFFE_PN0P_  (.CLK(clknet_leaf_235_clk_p2c),
    .RESET_B(net832),
    .D(_00336_),
    .Q_N(_06465_),
    .Q(\shift_storage.storage [120]));
 sg13g2_dfrbp_1 \shift_storage.storage[1210]$_SDFFE_PN0P_  (.CLK(clknet_leaf_202_clk_p2c),
    .RESET_B(net833),
    .D(_00337_),
    .Q_N(_06464_),
    .Q(\shift_storage.storage [1210]));
 sg13g2_dfrbp_1 \shift_storage.storage[1211]$_SDFFE_PN0P_  (.CLK(clknet_leaf_202_clk_p2c),
    .RESET_B(net834),
    .D(_00338_),
    .Q_N(_06463_),
    .Q(\shift_storage.storage [1211]));
 sg13g2_dfrbp_1 \shift_storage.storage[1212]$_SDFFE_PN0P_  (.CLK(clknet_leaf_235_clk_p2c),
    .RESET_B(net835),
    .D(_00339_),
    .Q_N(_06462_),
    .Q(\shift_storage.storage [1212]));
 sg13g2_dfrbp_1 \shift_storage.storage[1213]$_SDFFE_PN0P_  (.CLK(clknet_leaf_233_clk_p2c),
    .RESET_B(net836),
    .D(_00340_),
    .Q_N(_06461_),
    .Q(\shift_storage.storage [1213]));
 sg13g2_dfrbp_1 \shift_storage.storage[1214]$_SDFFE_PN0P_  (.CLK(clknet_leaf_204_clk_p2c),
    .RESET_B(net837),
    .D(_00341_),
    .Q_N(_06460_),
    .Q(\shift_storage.storage [1214]));
 sg13g2_dfrbp_1 \shift_storage.storage[1215]$_SDFFE_PN0P_  (.CLK(clknet_leaf_204_clk_p2c),
    .RESET_B(net838),
    .D(_00342_),
    .Q_N(_06459_),
    .Q(\shift_storage.storage [1215]));
 sg13g2_dfrbp_1 \shift_storage.storage[1216]$_SDFFE_PN0P_  (.CLK(clknet_leaf_204_clk_p2c),
    .RESET_B(net839),
    .D(_00343_),
    .Q_N(_06458_),
    .Q(\shift_storage.storage [1216]));
 sg13g2_dfrbp_1 \shift_storage.storage[1217]$_SDFFE_PN0P_  (.CLK(clknet_leaf_204_clk_p2c),
    .RESET_B(net840),
    .D(_00344_),
    .Q_N(_06457_),
    .Q(\shift_storage.storage [1217]));
 sg13g2_dfrbp_1 \shift_storage.storage[1218]$_SDFFE_PN0P_  (.CLK(clknet_leaf_233_clk_p2c),
    .RESET_B(net841),
    .D(_00345_),
    .Q_N(_06456_),
    .Q(\shift_storage.storage [1218]));
 sg13g2_dfrbp_1 \shift_storage.storage[1219]$_SDFFE_PN0P_  (.CLK(clknet_leaf_205_clk_p2c),
    .RESET_B(net842),
    .D(_00346_),
    .Q_N(_06455_),
    .Q(\shift_storage.storage [1219]));
 sg13g2_dfrbp_1 \shift_storage.storage[121]$_SDFFE_PN0P_  (.CLK(clknet_leaf_233_clk_p2c),
    .RESET_B(net843),
    .D(_00347_),
    .Q_N(_06454_),
    .Q(\shift_storage.storage [121]));
 sg13g2_dfrbp_1 \shift_storage.storage[1220]$_SDFFE_PN0P_  (.CLK(clknet_leaf_205_clk_p2c),
    .RESET_B(net844),
    .D(_00348_),
    .Q_N(_06453_),
    .Q(\shift_storage.storage [1220]));
 sg13g2_dfrbp_1 \shift_storage.storage[1221]$_SDFFE_PN0P_  (.CLK(clknet_leaf_232_clk_p2c),
    .RESET_B(net845),
    .D(_00349_),
    .Q_N(_06452_),
    .Q(\shift_storage.storage [1221]));
 sg13g2_dfrbp_1 \shift_storage.storage[1222]$_SDFFE_PN0P_  (.CLK(clknet_leaf_232_clk_p2c),
    .RESET_B(net846),
    .D(_00350_),
    .Q_N(_06451_),
    .Q(\shift_storage.storage [1222]));
 sg13g2_dfrbp_1 \shift_storage.storage[1223]$_SDFFE_PN0P_  (.CLK(clknet_leaf_233_clk_p2c),
    .RESET_B(net847),
    .D(_00351_),
    .Q_N(_06450_),
    .Q(\shift_storage.storage [1223]));
 sg13g2_dfrbp_1 \shift_storage.storage[1224]$_SDFFE_PN0P_  (.CLK(clknet_leaf_233_clk_p2c),
    .RESET_B(net848),
    .D(_00352_),
    .Q_N(_06449_),
    .Q(\shift_storage.storage [1224]));
 sg13g2_dfrbp_1 \shift_storage.storage[1225]$_SDFFE_PN0P_  (.CLK(clknet_leaf_233_clk_p2c),
    .RESET_B(net849),
    .D(_00353_),
    .Q_N(_06448_),
    .Q(\shift_storage.storage [1225]));
 sg13g2_dfrbp_1 \shift_storage.storage[1226]$_SDFFE_PN0P_  (.CLK(clknet_leaf_234_clk_p2c),
    .RESET_B(net850),
    .D(_00354_),
    .Q_N(_06447_),
    .Q(\shift_storage.storage [1226]));
 sg13g2_dfrbp_1 \shift_storage.storage[1227]$_SDFFE_PN0P_  (.CLK(clknet_leaf_231_clk_p2c),
    .RESET_B(net851),
    .D(_00355_),
    .Q_N(_06446_),
    .Q(\shift_storage.storage [1227]));
 sg13g2_dfrbp_1 \shift_storage.storage[1228]$_SDFFE_PN0P_  (.CLK(clknet_leaf_232_clk_p2c),
    .RESET_B(net852),
    .D(_00356_),
    .Q_N(_06445_),
    .Q(\shift_storage.storage [1228]));
 sg13g2_dfrbp_1 \shift_storage.storage[1229]$_SDFFE_PN0P_  (.CLK(clknet_leaf_232_clk_p2c),
    .RESET_B(net853),
    .D(_00357_),
    .Q_N(_06444_),
    .Q(\shift_storage.storage [1229]));
 sg13g2_dfrbp_1 \shift_storage.storage[122]$_SDFFE_PN0P_  (.CLK(clknet_leaf_232_clk_p2c),
    .RESET_B(net854),
    .D(_00358_),
    .Q_N(_06443_),
    .Q(\shift_storage.storage [122]));
 sg13g2_dfrbp_1 \shift_storage.storage[1230]$_SDFFE_PN0P_  (.CLK(clknet_leaf_231_clk_p2c),
    .RESET_B(net855),
    .D(_00359_),
    .Q_N(_06442_),
    .Q(\shift_storage.storage [1230]));
 sg13g2_dfrbp_1 \shift_storage.storage[1231]$_SDFFE_PN0P_  (.CLK(clknet_leaf_230_clk_p2c),
    .RESET_B(net856),
    .D(_00360_),
    .Q_N(_06441_),
    .Q(\shift_storage.storage [1231]));
 sg13g2_dfrbp_1 \shift_storage.storage[1232]$_SDFFE_PN0P_  (.CLK(clknet_leaf_231_clk_p2c),
    .RESET_B(net857),
    .D(_00361_),
    .Q_N(_06440_),
    .Q(\shift_storage.storage [1232]));
 sg13g2_dfrbp_1 \shift_storage.storage[1233]$_SDFFE_PN0P_  (.CLK(clknet_leaf_231_clk_p2c),
    .RESET_B(net858),
    .D(_00362_),
    .Q_N(_06439_),
    .Q(\shift_storage.storage [1233]));
 sg13g2_dfrbp_1 \shift_storage.storage[1234]$_SDFFE_PN0P_  (.CLK(clknet_leaf_230_clk_p2c),
    .RESET_B(net859),
    .D(_00363_),
    .Q_N(_06438_),
    .Q(\shift_storage.storage [1234]));
 sg13g2_dfrbp_1 \shift_storage.storage[1235]$_SDFFE_PN0P_  (.CLK(clknet_leaf_230_clk_p2c),
    .RESET_B(net860),
    .D(_00364_),
    .Q_N(_06437_),
    .Q(\shift_storage.storage [1235]));
 sg13g2_dfrbp_1 \shift_storage.storage[1236]$_SDFFE_PN0P_  (.CLK(clknet_leaf_230_clk_p2c),
    .RESET_B(net861),
    .D(_00365_),
    .Q_N(_06436_),
    .Q(\shift_storage.storage [1236]));
 sg13g2_dfrbp_1 \shift_storage.storage[1237]$_SDFFE_PN0P_  (.CLK(clknet_leaf_230_clk_p2c),
    .RESET_B(net862),
    .D(_00366_),
    .Q_N(_06435_),
    .Q(\shift_storage.storage [1237]));
 sg13g2_dfrbp_1 \shift_storage.storage[1238]$_SDFFE_PN0P_  (.CLK(clknet_leaf_224_clk_p2c),
    .RESET_B(net863),
    .D(_00367_),
    .Q_N(_06434_),
    .Q(\shift_storage.storage [1238]));
 sg13g2_dfrbp_1 \shift_storage.storage[1239]$_SDFFE_PN0P_  (.CLK(clknet_leaf_223_clk_p2c),
    .RESET_B(net864),
    .D(_00368_),
    .Q_N(_06433_),
    .Q(\shift_storage.storage [1239]));
 sg13g2_dfrbp_1 \shift_storage.storage[123]$_SDFFE_PN0P_  (.CLK(clknet_leaf_232_clk_p2c),
    .RESET_B(net865),
    .D(_00369_),
    .Q_N(_06432_),
    .Q(\shift_storage.storage [123]));
 sg13g2_dfrbp_1 \shift_storage.storage[1240]$_SDFFE_PN0P_  (.CLK(clknet_leaf_223_clk_p2c),
    .RESET_B(net866),
    .D(_00370_),
    .Q_N(_06431_),
    .Q(\shift_storage.storage [1240]));
 sg13g2_dfrbp_1 \shift_storage.storage[1241]$_SDFFE_PN0P_  (.CLK(clknet_leaf_223_clk_p2c),
    .RESET_B(net867),
    .D(_00371_),
    .Q_N(_06430_),
    .Q(\shift_storage.storage [1241]));
 sg13g2_dfrbp_1 \shift_storage.storage[1242]$_SDFFE_PN0P_  (.CLK(clknet_leaf_223_clk_p2c),
    .RESET_B(net868),
    .D(_00372_),
    .Q_N(_06429_),
    .Q(\shift_storage.storage [1242]));
 sg13g2_dfrbp_1 \shift_storage.storage[1243]$_SDFFE_PN0P_  (.CLK(clknet_leaf_222_clk_p2c),
    .RESET_B(net869),
    .D(_00373_),
    .Q_N(_06428_),
    .Q(\shift_storage.storage [1243]));
 sg13g2_dfrbp_1 \shift_storage.storage[1244]$_SDFFE_PN0P_  (.CLK(clknet_leaf_222_clk_p2c),
    .RESET_B(net870),
    .D(_00374_),
    .Q_N(_06427_),
    .Q(\shift_storage.storage [1244]));
 sg13g2_dfrbp_1 \shift_storage.storage[1245]$_SDFFE_PN0P_  (.CLK(clknet_leaf_223_clk_p2c),
    .RESET_B(net871),
    .D(_00375_),
    .Q_N(_06426_),
    .Q(\shift_storage.storage [1245]));
 sg13g2_dfrbp_1 \shift_storage.storage[1246]$_SDFFE_PN0P_  (.CLK(clknet_leaf_222_clk_p2c),
    .RESET_B(net872),
    .D(_00376_),
    .Q_N(_06425_),
    .Q(\shift_storage.storage [1246]));
 sg13g2_dfrbp_1 \shift_storage.storage[1247]$_SDFFE_PN0P_  (.CLK(clknet_leaf_223_clk_p2c),
    .RESET_B(net873),
    .D(_00377_),
    .Q_N(_06424_),
    .Q(\shift_storage.storage [1247]));
 sg13g2_dfrbp_1 \shift_storage.storage[1248]$_SDFFE_PN0P_  (.CLK(clknet_leaf_222_clk_p2c),
    .RESET_B(net874),
    .D(_00378_),
    .Q_N(_06423_),
    .Q(\shift_storage.storage [1248]));
 sg13g2_dfrbp_1 \shift_storage.storage[1249]$_SDFFE_PN0P_  (.CLK(clknet_leaf_222_clk_p2c),
    .RESET_B(net875),
    .D(_00379_),
    .Q_N(_06422_),
    .Q(\shift_storage.storage [1249]));
 sg13g2_dfrbp_1 \shift_storage.storage[124]$_SDFFE_PN0P_  (.CLK(clknet_leaf_221_clk_p2c),
    .RESET_B(net876),
    .D(_00380_),
    .Q_N(_06421_),
    .Q(\shift_storage.storage [124]));
 sg13g2_dfrbp_1 \shift_storage.storage[1250]$_SDFFE_PN0P_  (.CLK(clknet_leaf_222_clk_p2c),
    .RESET_B(net877),
    .D(_00381_),
    .Q_N(_06420_),
    .Q(\shift_storage.storage [1250]));
 sg13g2_dfrbp_1 \shift_storage.storage[1251]$_SDFFE_PN0P_  (.CLK(clknet_leaf_220_clk_p2c),
    .RESET_B(net878),
    .D(_00382_),
    .Q_N(_06419_),
    .Q(\shift_storage.storage [1251]));
 sg13g2_dfrbp_1 \shift_storage.storage[1252]$_SDFFE_PN0P_  (.CLK(clknet_leaf_220_clk_p2c),
    .RESET_B(net879),
    .D(_00383_),
    .Q_N(_06418_),
    .Q(\shift_storage.storage [1252]));
 sg13g2_dfrbp_1 \shift_storage.storage[1253]$_SDFFE_PN0P_  (.CLK(clknet_leaf_220_clk_p2c),
    .RESET_B(net880),
    .D(_00384_),
    .Q_N(_06417_),
    .Q(\shift_storage.storage [1253]));
 sg13g2_dfrbp_1 \shift_storage.storage[1254]$_SDFFE_PN0P_  (.CLK(clknet_leaf_220_clk_p2c),
    .RESET_B(net881),
    .D(_00385_),
    .Q_N(_06416_),
    .Q(\shift_storage.storage [1254]));
 sg13g2_dfrbp_1 \shift_storage.storage[1255]$_SDFFE_PN0P_  (.CLK(clknet_leaf_222_clk_p2c),
    .RESET_B(net882),
    .D(_00386_),
    .Q_N(_06415_),
    .Q(\shift_storage.storage [1255]));
 sg13g2_dfrbp_1 \shift_storage.storage[1256]$_SDFFE_PN0P_  (.CLK(clknet_leaf_221_clk_p2c),
    .RESET_B(net883),
    .D(_00387_),
    .Q_N(_06414_),
    .Q(\shift_storage.storage [1256]));
 sg13g2_dfrbp_1 \shift_storage.storage[1257]$_SDFFE_PN0P_  (.CLK(clknet_leaf_221_clk_p2c),
    .RESET_B(net884),
    .D(_00388_),
    .Q_N(_06413_),
    .Q(\shift_storage.storage [1257]));
 sg13g2_dfrbp_1 \shift_storage.storage[1258]$_SDFFE_PN0P_  (.CLK(clknet_leaf_221_clk_p2c),
    .RESET_B(net885),
    .D(_00389_),
    .Q_N(_06412_),
    .Q(\shift_storage.storage [1258]));
 sg13g2_dfrbp_1 \shift_storage.storage[1259]$_SDFFE_PN0P_  (.CLK(clknet_leaf_221_clk_p2c),
    .RESET_B(net886),
    .D(_00390_),
    .Q_N(_06411_),
    .Q(\shift_storage.storage [1259]));
 sg13g2_dfrbp_1 \shift_storage.storage[125]$_SDFFE_PN0P_  (.CLK(clknet_leaf_221_clk_p2c),
    .RESET_B(net887),
    .D(_00391_),
    .Q_N(_06410_),
    .Q(\shift_storage.storage [125]));
 sg13g2_dfrbp_1 \shift_storage.storage[1260]$_SDFFE_PN0P_  (.CLK(clknet_leaf_220_clk_p2c),
    .RESET_B(net888),
    .D(_00392_),
    .Q_N(_06409_),
    .Q(\shift_storage.storage [1260]));
 sg13g2_dfrbp_1 \shift_storage.storage[1261]$_SDFFE_PN0P_  (.CLK(clknet_leaf_220_clk_p2c),
    .RESET_B(net889),
    .D(_00393_),
    .Q_N(_06408_),
    .Q(\shift_storage.storage [1261]));
 sg13g2_dfrbp_1 \shift_storage.storage[1262]$_SDFFE_PN0P_  (.CLK(clknet_leaf_219_clk_p2c),
    .RESET_B(net890),
    .D(_00394_),
    .Q_N(_06407_),
    .Q(\shift_storage.storage [1262]));
 sg13g2_dfrbp_1 \shift_storage.storage[1263]$_SDFFE_PN0P_  (.CLK(clknet_leaf_219_clk_p2c),
    .RESET_B(net891),
    .D(_00395_),
    .Q_N(_06406_),
    .Q(\shift_storage.storage [1263]));
 sg13g2_dfrbp_1 \shift_storage.storage[1264]$_SDFFE_PN0P_  (.CLK(clknet_leaf_219_clk_p2c),
    .RESET_B(net892),
    .D(_00396_),
    .Q_N(_06405_),
    .Q(\shift_storage.storage [1264]));
 sg13g2_dfrbp_1 \shift_storage.storage[1265]$_SDFFE_PN0P_  (.CLK(clknet_leaf_218_clk_p2c),
    .RESET_B(net893),
    .D(_00397_),
    .Q_N(_06404_),
    .Q(\shift_storage.storage [1265]));
 sg13g2_dfrbp_1 \shift_storage.storage[1266]$_SDFFE_PN0P_  (.CLK(clknet_leaf_218_clk_p2c),
    .RESET_B(net894),
    .D(_00398_),
    .Q_N(_06403_),
    .Q(\shift_storage.storage [1266]));
 sg13g2_dfrbp_1 \shift_storage.storage[1267]$_SDFFE_PN0P_  (.CLK(clknet_leaf_218_clk_p2c),
    .RESET_B(net895),
    .D(_00399_),
    .Q_N(_06402_),
    .Q(\shift_storage.storage [1267]));
 sg13g2_dfrbp_1 \shift_storage.storage[1268]$_SDFFE_PN0P_  (.CLK(clknet_leaf_218_clk_p2c),
    .RESET_B(net896),
    .D(_00400_),
    .Q_N(_06401_),
    .Q(\shift_storage.storage [1268]));
 sg13g2_dfrbp_1 \shift_storage.storage[1269]$_SDFFE_PN0P_  (.CLK(clknet_leaf_218_clk_p2c),
    .RESET_B(net897),
    .D(_00401_),
    .Q_N(_06400_),
    .Q(\shift_storage.storage [1269]));
 sg13g2_dfrbp_1 \shift_storage.storage[126]$_SDFFE_PN0P_  (.CLK(clknet_leaf_218_clk_p2c),
    .RESET_B(net898),
    .D(_00402_),
    .Q_N(_06399_),
    .Q(\shift_storage.storage [126]));
 sg13g2_dfrbp_1 \shift_storage.storage[1270]$_SDFFE_PN0P_  (.CLK(clknet_leaf_217_clk_p2c),
    .RESET_B(net899),
    .D(_00403_),
    .Q_N(_06398_),
    .Q(\shift_storage.storage [1270]));
 sg13g2_dfrbp_1 \shift_storage.storage[1271]$_SDFFE_PN0P_  (.CLK(clknet_leaf_217_clk_p2c),
    .RESET_B(net900),
    .D(_00404_),
    .Q_N(_06397_),
    .Q(\shift_storage.storage [1271]));
 sg13g2_dfrbp_1 \shift_storage.storage[1272]$_SDFFE_PN0P_  (.CLK(clknet_leaf_217_clk_p2c),
    .RESET_B(net901),
    .D(_00405_),
    .Q_N(_06396_),
    .Q(\shift_storage.storage [1272]));
 sg13g2_dfrbp_1 \shift_storage.storage[1273]$_SDFFE_PN0P_  (.CLK(clknet_leaf_217_clk_p2c),
    .RESET_B(net902),
    .D(_00406_),
    .Q_N(_06395_),
    .Q(\shift_storage.storage [1273]));
 sg13g2_dfrbp_1 \shift_storage.storage[1274]$_SDFFE_PN0P_  (.CLK(clknet_leaf_217_clk_p2c),
    .RESET_B(net903),
    .D(_00407_),
    .Q_N(_06394_),
    .Q(\shift_storage.storage [1274]));
 sg13g2_dfrbp_1 \shift_storage.storage[1275]$_SDFFE_PN0P_  (.CLK(clknet_leaf_216_clk_p2c),
    .RESET_B(net904),
    .D(_00408_),
    .Q_N(_06393_),
    .Q(\shift_storage.storage [1275]));
 sg13g2_dfrbp_1 \shift_storage.storage[1276]$_SDFFE_PN0P_  (.CLK(clknet_leaf_216_clk_p2c),
    .RESET_B(net905),
    .D(_00409_),
    .Q_N(_06392_),
    .Q(\shift_storage.storage [1276]));
 sg13g2_dfrbp_1 \shift_storage.storage[1277]$_SDFFE_PN0P_  (.CLK(clknet_leaf_216_clk_p2c),
    .RESET_B(net906),
    .D(_00410_),
    .Q_N(_06391_),
    .Q(\shift_storage.storage [1277]));
 sg13g2_dfrbp_1 \shift_storage.storage[1278]$_SDFFE_PN0P_  (.CLK(clknet_leaf_217_clk_p2c),
    .RESET_B(net907),
    .D(_00411_),
    .Q_N(_06390_),
    .Q(\shift_storage.storage [1278]));
 sg13g2_dfrbp_1 \shift_storage.storage[1279]$_SDFFE_PN0P_  (.CLK(clknet_leaf_216_clk_p2c),
    .RESET_B(net908),
    .D(_00412_),
    .Q_N(_06389_),
    .Q(\shift_storage.storage [1279]));
 sg13g2_dfrbp_1 \shift_storage.storage[127]$_SDFFE_PN0P_  (.CLK(clknet_leaf_207_clk_p2c),
    .RESET_B(net909),
    .D(_00413_),
    .Q_N(_06388_),
    .Q(\shift_storage.storage [127]));
 sg13g2_dfrbp_1 \shift_storage.storage[1280]$_SDFFE_PN0P_  (.CLK(clknet_leaf_207_clk_p2c),
    .RESET_B(net910),
    .D(_00414_),
    .Q_N(_06387_),
    .Q(\shift_storage.storage [1280]));
 sg13g2_dfrbp_1 \shift_storage.storage[1281]$_SDFFE_PN0P_  (.CLK(clknet_leaf_206_clk_p2c),
    .RESET_B(net911),
    .D(_00415_),
    .Q_N(_06386_),
    .Q(\shift_storage.storage [1281]));
 sg13g2_dfrbp_1 \shift_storage.storage[1282]$_SDFFE_PN0P_  (.CLK(clknet_leaf_206_clk_p2c),
    .RESET_B(net912),
    .D(_00416_),
    .Q_N(_06385_),
    .Q(\shift_storage.storage [1282]));
 sg13g2_dfrbp_1 \shift_storage.storage[1283]$_SDFFE_PN0P_  (.CLK(clknet_leaf_206_clk_p2c),
    .RESET_B(net913),
    .D(_00417_),
    .Q_N(_06384_),
    .Q(\shift_storage.storage [1283]));
 sg13g2_dfrbp_1 \shift_storage.storage[1284]$_SDFFE_PN0P_  (.CLK(clknet_leaf_205_clk_p2c),
    .RESET_B(net914),
    .D(_00418_),
    .Q_N(_06383_),
    .Q(\shift_storage.storage [1284]));
 sg13g2_dfrbp_1 \shift_storage.storage[1285]$_SDFFE_PN0P_  (.CLK(clknet_leaf_205_clk_p2c),
    .RESET_B(net915),
    .D(_00419_),
    .Q_N(_06382_),
    .Q(\shift_storage.storage [1285]));
 sg13g2_dfrbp_1 \shift_storage.storage[1286]$_SDFFE_PN0P_  (.CLK(clknet_leaf_205_clk_p2c),
    .RESET_B(net916),
    .D(_00420_),
    .Q_N(_06381_),
    .Q(\shift_storage.storage [1286]));
 sg13g2_dfrbp_1 \shift_storage.storage[1287]$_SDFFE_PN0P_  (.CLK(clknet_leaf_204_clk_p2c),
    .RESET_B(net917),
    .D(_00421_),
    .Q_N(_06380_),
    .Q(\shift_storage.storage [1287]));
 sg13g2_dfrbp_1 \shift_storage.storage[1288]$_SDFFE_PN0P_  (.CLK(clknet_leaf_203_clk_p2c),
    .RESET_B(net918),
    .D(_00422_),
    .Q_N(_06379_),
    .Q(\shift_storage.storage [1288]));
 sg13g2_dfrbp_1 \shift_storage.storage[1289]$_SDFFE_PN0P_  (.CLK(clknet_leaf_206_clk_p2c),
    .RESET_B(net919),
    .D(_00423_),
    .Q_N(_06378_),
    .Q(\shift_storage.storage [1289]));
 sg13g2_dfrbp_1 \shift_storage.storage[128]$_SDFFE_PN0P_  (.CLK(clknet_leaf_203_clk_p2c),
    .RESET_B(net920),
    .D(_00424_),
    .Q_N(_06377_),
    .Q(\shift_storage.storage [128]));
 sg13g2_dfrbp_1 \shift_storage.storage[1290]$_SDFFE_PN0P_  (.CLK(clknet_leaf_206_clk_p2c),
    .RESET_B(net921),
    .D(_00425_),
    .Q_N(_06376_),
    .Q(\shift_storage.storage [1290]));
 sg13g2_dfrbp_1 \shift_storage.storage[1291]$_SDFFE_PN0P_  (.CLK(clknet_leaf_203_clk_p2c),
    .RESET_B(net922),
    .D(_00426_),
    .Q_N(_06375_),
    .Q(\shift_storage.storage [1291]));
 sg13g2_dfrbp_1 \shift_storage.storage[1292]$_SDFFE_PN0P_  (.CLK(clknet_leaf_203_clk_p2c),
    .RESET_B(net923),
    .D(_00427_),
    .Q_N(_06374_),
    .Q(\shift_storage.storage [1292]));
 sg13g2_dfrbp_1 \shift_storage.storage[1293]$_SDFFE_PN0P_  (.CLK(clknet_leaf_202_clk_p2c),
    .RESET_B(net924),
    .D(_00428_),
    .Q_N(_06373_),
    .Q(\shift_storage.storage [1293]));
 sg13g2_dfrbp_1 \shift_storage.storage[1294]$_SDFFE_PN0P_  (.CLK(clknet_leaf_203_clk_p2c),
    .RESET_B(net925),
    .D(_00429_),
    .Q_N(_06372_),
    .Q(\shift_storage.storage [1294]));
 sg13g2_dfrbp_1 \shift_storage.storage[1295]$_SDFFE_PN0P_  (.CLK(clknet_leaf_199_clk_p2c),
    .RESET_B(net926),
    .D(_00430_),
    .Q_N(_06371_),
    .Q(\shift_storage.storage [1295]));
 sg13g2_dfrbp_1 \shift_storage.storage[1296]$_SDFFE_PN0P_  (.CLK(clknet_leaf_199_clk_p2c),
    .RESET_B(net927),
    .D(_00431_),
    .Q_N(_06370_),
    .Q(\shift_storage.storage [1296]));
 sg13g2_dfrbp_1 \shift_storage.storage[1297]$_SDFFE_PN0P_  (.CLK(clknet_leaf_200_clk_p2c),
    .RESET_B(net928),
    .D(_00432_),
    .Q_N(_06369_),
    .Q(\shift_storage.storage [1297]));
 sg13g2_dfrbp_1 \shift_storage.storage[1298]$_SDFFE_PN0P_  (.CLK(clknet_leaf_200_clk_p2c),
    .RESET_B(net929),
    .D(_00433_),
    .Q_N(_06368_),
    .Q(\shift_storage.storage [1298]));
 sg13g2_dfrbp_1 \shift_storage.storage[1299]$_SDFFE_PN0P_  (.CLK(clknet_leaf_200_clk_p2c),
    .RESET_B(net930),
    .D(_00434_),
    .Q_N(_06367_),
    .Q(\shift_storage.storage [1299]));
 sg13g2_dfrbp_1 \shift_storage.storage[129]$_SDFFE_PN0P_  (.CLK(clknet_leaf_199_clk_p2c),
    .RESET_B(net931),
    .D(_00435_),
    .Q_N(_06366_),
    .Q(\shift_storage.storage [129]));
 sg13g2_dfrbp_1 \shift_storage.storage[12]$_SDFFE_PN0P_  (.CLK(clknet_leaf_200_clk_p2c),
    .RESET_B(net932),
    .D(_00436_),
    .Q_N(_06365_),
    .Q(\shift_storage.storage [12]));
 sg13g2_dfrbp_1 \shift_storage.storage[1300]$_SDFFE_PN0P_  (.CLK(clknet_leaf_200_clk_p2c),
    .RESET_B(net933),
    .D(_00437_),
    .Q_N(_06364_),
    .Q(\shift_storage.storage [1300]));
 sg13g2_dfrbp_1 \shift_storage.storage[1301]$_SDFFE_PN0P_  (.CLK(clknet_leaf_199_clk_p2c),
    .RESET_B(net934),
    .D(_00438_),
    .Q_N(_06363_),
    .Q(\shift_storage.storage [1301]));
 sg13g2_dfrbp_1 \shift_storage.storage[1302]$_SDFFE_PN0P_  (.CLK(clknet_leaf_199_clk_p2c),
    .RESET_B(net935),
    .D(_00439_),
    .Q_N(_06362_),
    .Q(\shift_storage.storage [1302]));
 sg13g2_dfrbp_1 \shift_storage.storage[1303]$_SDFFE_PN0P_  (.CLK(clknet_leaf_199_clk_p2c),
    .RESET_B(net936),
    .D(_00440_),
    .Q_N(_06361_),
    .Q(\shift_storage.storage [1303]));
 sg13g2_dfrbp_1 \shift_storage.storage[1304]$_SDFFE_PN0P_  (.CLK(clknet_leaf_210_clk_p2c),
    .RESET_B(net937),
    .D(_00441_),
    .Q_N(_06360_),
    .Q(\shift_storage.storage [1304]));
 sg13g2_dfrbp_1 \shift_storage.storage[1305]$_SDFFE_PN0P_  (.CLK(clknet_leaf_210_clk_p2c),
    .RESET_B(net938),
    .D(_00442_),
    .Q_N(_06359_),
    .Q(\shift_storage.storage [1305]));
 sg13g2_dfrbp_1 \shift_storage.storage[1306]$_SDFFE_PN0P_  (.CLK(clknet_leaf_210_clk_p2c),
    .RESET_B(net939),
    .D(_00443_),
    .Q_N(_06358_),
    .Q(\shift_storage.storage [1306]));
 sg13g2_dfrbp_1 \shift_storage.storage[1307]$_SDFFE_PN0P_  (.CLK(clknet_leaf_210_clk_p2c),
    .RESET_B(net940),
    .D(_00444_),
    .Q_N(_06357_),
    .Q(\shift_storage.storage [1307]));
 sg13g2_dfrbp_1 \shift_storage.storage[1308]$_SDFFE_PN0P_  (.CLK(clknet_leaf_209_clk_p2c),
    .RESET_B(net941),
    .D(_00445_),
    .Q_N(_06356_),
    .Q(\shift_storage.storage [1308]));
 sg13g2_dfrbp_1 \shift_storage.storage[1309]$_SDFFE_PN0P_  (.CLK(clknet_leaf_210_clk_p2c),
    .RESET_B(net942),
    .D(_00446_),
    .Q_N(_06355_),
    .Q(\shift_storage.storage [1309]));
 sg13g2_dfrbp_1 \shift_storage.storage[130]$_SDFFE_PN0P_  (.CLK(clknet_leaf_209_clk_p2c),
    .RESET_B(net943),
    .D(_00447_),
    .Q_N(_06354_),
    .Q(\shift_storage.storage [130]));
 sg13g2_dfrbp_1 \shift_storage.storage[1310]$_SDFFE_PN0P_  (.CLK(clknet_leaf_210_clk_p2c),
    .RESET_B(net944),
    .D(_00448_),
    .Q_N(_06353_),
    .Q(\shift_storage.storage [1310]));
 sg13g2_dfrbp_1 \shift_storage.storage[1311]$_SDFFE_PN0P_  (.CLK(clknet_leaf_207_clk_p2c),
    .RESET_B(net945),
    .D(_00449_),
    .Q_N(_06352_),
    .Q(\shift_storage.storage [1311]));
 sg13g2_dfrbp_1 \shift_storage.storage[1312]$_SDFFE_PN0P_  (.CLK(clknet_leaf_207_clk_p2c),
    .RESET_B(net946),
    .D(_00450_),
    .Q_N(_06351_),
    .Q(\shift_storage.storage [1312]));
 sg13g2_dfrbp_1 \shift_storage.storage[1313]$_SDFFE_PN0P_  (.CLK(clknet_leaf_207_clk_p2c),
    .RESET_B(net947),
    .D(_00451_),
    .Q_N(_06350_),
    .Q(\shift_storage.storage [1313]));
 sg13g2_dfrbp_1 \shift_storage.storage[1314]$_SDFFE_PN0P_  (.CLK(clknet_leaf_209_clk_p2c),
    .RESET_B(net948),
    .D(_00452_),
    .Q_N(_06349_),
    .Q(\shift_storage.storage [1314]));
 sg13g2_dfrbp_1 \shift_storage.storage[1315]$_SDFFE_PN0P_  (.CLK(clknet_leaf_209_clk_p2c),
    .RESET_B(net949),
    .D(_00453_),
    .Q_N(_06348_),
    .Q(\shift_storage.storage [1315]));
 sg13g2_dfrbp_1 \shift_storage.storage[1316]$_SDFFE_PN0P_  (.CLK(clknet_leaf_208_clk_p2c),
    .RESET_B(net950),
    .D(_00454_),
    .Q_N(_06347_),
    .Q(\shift_storage.storage [1316]));
 sg13g2_dfrbp_1 \shift_storage.storage[1317]$_SDFFE_PN0P_  (.CLK(clknet_leaf_208_clk_p2c),
    .RESET_B(net951),
    .D(_00455_),
    .Q_N(_06346_),
    .Q(\shift_storage.storage [1317]));
 sg13g2_dfrbp_1 \shift_storage.storage[1318]$_SDFFE_PN0P_  (.CLK(clknet_leaf_207_clk_p2c),
    .RESET_B(net952),
    .D(_00456_),
    .Q_N(_06345_),
    .Q(\shift_storage.storage [1318]));
 sg13g2_dfrbp_1 \shift_storage.storage[1319]$_SDFFE_PN0P_  (.CLK(clknet_leaf_208_clk_p2c),
    .RESET_B(net953),
    .D(_00457_),
    .Q_N(_06344_),
    .Q(\shift_storage.storage [1319]));
 sg13g2_dfrbp_1 \shift_storage.storage[131]$_SDFFE_PN0P_  (.CLK(clknet_leaf_209_clk_p2c),
    .RESET_B(net954),
    .D(_00458_),
    .Q_N(_06343_),
    .Q(\shift_storage.storage [131]));
 sg13g2_dfrbp_1 \shift_storage.storage[1320]$_SDFFE_PN0P_  (.CLK(clknet_leaf_208_clk_p2c),
    .RESET_B(net955),
    .D(_00459_),
    .Q_N(_06342_),
    .Q(\shift_storage.storage [1320]));
 sg13g2_dfrbp_1 \shift_storage.storage[1321]$_SDFFE_PN0P_  (.CLK(clknet_leaf_216_clk_p2c),
    .RESET_B(net956),
    .D(_00460_),
    .Q_N(_06341_),
    .Q(\shift_storage.storage [1321]));
 sg13g2_dfrbp_1 \shift_storage.storage[1322]$_SDFFE_PN0P_  (.CLK(clknet_leaf_216_clk_p2c),
    .RESET_B(net957),
    .D(_00461_),
    .Q_N(_06340_),
    .Q(\shift_storage.storage [1322]));
 sg13g2_dfrbp_1 \shift_storage.storage[1323]$_SDFFE_PN0P_  (.CLK(clknet_leaf_216_clk_p2c),
    .RESET_B(net958),
    .D(_00462_),
    .Q_N(_06339_),
    .Q(\shift_storage.storage [1323]));
 sg13g2_dfrbp_1 \shift_storage.storage[1324]$_SDFFE_PN0P_  (.CLK(clknet_leaf_215_clk_p2c),
    .RESET_B(net959),
    .D(_00463_),
    .Q_N(_06338_),
    .Q(\shift_storage.storage [1324]));
 sg13g2_dfrbp_1 \shift_storage.storage[1325]$_SDFFE_PN0P_  (.CLK(clknet_leaf_215_clk_p2c),
    .RESET_B(net960),
    .D(_00464_),
    .Q_N(_06337_),
    .Q(\shift_storage.storage [1325]));
 sg13g2_dfrbp_1 \shift_storage.storage[1326]$_SDFFE_PN0P_  (.CLK(clknet_leaf_215_clk_p2c),
    .RESET_B(net961),
    .D(_00465_),
    .Q_N(_06336_),
    .Q(\shift_storage.storage [1326]));
 sg13g2_dfrbp_1 \shift_storage.storage[1327]$_SDFFE_PN0P_  (.CLK(clknet_leaf_215_clk_p2c),
    .RESET_B(net962),
    .D(_00466_),
    .Q_N(_06335_),
    .Q(\shift_storage.storage [1327]));
 sg13g2_dfrbp_1 \shift_storage.storage[1328]$_SDFFE_PN0P_  (.CLK(clknet_leaf_208_clk_p2c),
    .RESET_B(net963),
    .D(_00467_),
    .Q_N(_06334_),
    .Q(\shift_storage.storage [1328]));
 sg13g2_dfrbp_1 \shift_storage.storage[1329]$_SDFFE_PN0P_  (.CLK(clknet_leaf_208_clk_p2c),
    .RESET_B(net964),
    .D(_00468_),
    .Q_N(_06333_),
    .Q(\shift_storage.storage [1329]));
 sg13g2_dfrbp_1 \shift_storage.storage[132]$_SDFFE_PN0P_  (.CLK(clknet_leaf_213_clk_p2c),
    .RESET_B(net965),
    .D(_00469_),
    .Q_N(_06332_),
    .Q(\shift_storage.storage [132]));
 sg13g2_dfrbp_1 \shift_storage.storage[1330]$_SDFFE_PN0P_  (.CLK(clknet_leaf_213_clk_p2c),
    .RESET_B(net966),
    .D(_00470_),
    .Q_N(_06331_),
    .Q(\shift_storage.storage [1330]));
 sg13g2_dfrbp_1 \shift_storage.storage[1331]$_SDFFE_PN0P_  (.CLK(clknet_leaf_213_clk_p2c),
    .RESET_B(net967),
    .D(_00471_),
    .Q_N(_06330_),
    .Q(\shift_storage.storage [1331]));
 sg13g2_dfrbp_1 \shift_storage.storage[1332]$_SDFFE_PN0P_  (.CLK(clknet_leaf_214_clk_p2c),
    .RESET_B(net968),
    .D(_00472_),
    .Q_N(_06329_),
    .Q(\shift_storage.storage [1332]));
 sg13g2_dfrbp_1 \shift_storage.storage[1333]$_SDFFE_PN0P_  (.CLK(clknet_leaf_213_clk_p2c),
    .RESET_B(net969),
    .D(_00473_),
    .Q_N(_06328_),
    .Q(\shift_storage.storage [1333]));
 sg13g2_dfrbp_1 \shift_storage.storage[1334]$_SDFFE_PN0P_  (.CLK(clknet_leaf_214_clk_p2c),
    .RESET_B(net970),
    .D(_00474_),
    .Q_N(_06327_),
    .Q(\shift_storage.storage [1334]));
 sg13g2_dfrbp_1 \shift_storage.storage[1335]$_SDFFE_PN0P_  (.CLK(clknet_leaf_214_clk_p2c),
    .RESET_B(net971),
    .D(_00475_),
    .Q_N(_06326_),
    .Q(\shift_storage.storage [1335]));
 sg13g2_dfrbp_1 \shift_storage.storage[1336]$_SDFFE_PN0P_  (.CLK(clknet_leaf_214_clk_p2c),
    .RESET_B(net972),
    .D(_00476_),
    .Q_N(_06325_),
    .Q(\shift_storage.storage [1336]));
 sg13g2_dfrbp_1 \shift_storage.storage[1337]$_SDFFE_PN0P_  (.CLK(clknet_leaf_214_clk_p2c),
    .RESET_B(net973),
    .D(_00477_),
    .Q_N(_06324_),
    .Q(\shift_storage.storage [1337]));
 sg13g2_dfrbp_1 \shift_storage.storage[1338]$_SDFFE_PN0P_  (.CLK(clknet_leaf_212_clk_p2c),
    .RESET_B(net974),
    .D(_00478_),
    .Q_N(_06323_),
    .Q(\shift_storage.storage [1338]));
 sg13g2_dfrbp_1 \shift_storage.storage[1339]$_SDFFE_PN0P_  (.CLK(clknet_leaf_212_clk_p2c),
    .RESET_B(net975),
    .D(_00479_),
    .Q_N(_06322_),
    .Q(\shift_storage.storage [1339]));
 sg13g2_dfrbp_1 \shift_storage.storage[133]$_SDFFE_PN0P_  (.CLK(clknet_leaf_213_clk_p2c),
    .RESET_B(net976),
    .D(_00480_),
    .Q_N(_06321_),
    .Q(\shift_storage.storage [133]));
 sg13g2_dfrbp_1 \shift_storage.storage[1340]$_SDFFE_PN0P_  (.CLK(clknet_leaf_212_clk_p2c),
    .RESET_B(net977),
    .D(_00481_),
    .Q_N(_06320_),
    .Q(\shift_storage.storage [1340]));
 sg13g2_dfrbp_1 \shift_storage.storage[1341]$_SDFFE_PN0P_  (.CLK(clknet_leaf_178_clk_p2c),
    .RESET_B(net978),
    .D(_00482_),
    .Q_N(_06319_),
    .Q(\shift_storage.storage [1341]));
 sg13g2_dfrbp_1 \shift_storage.storage[1342]$_SDFFE_PN0P_  (.CLK(clknet_leaf_178_clk_p2c),
    .RESET_B(net979),
    .D(_00483_),
    .Q_N(_06318_),
    .Q(\shift_storage.storage [1342]));
 sg13g2_dfrbp_1 \shift_storage.storage[1343]$_SDFFE_PN0P_  (.CLK(clknet_leaf_212_clk_p2c),
    .RESET_B(net980),
    .D(_00484_),
    .Q_N(_06317_),
    .Q(\shift_storage.storage [1343]));
 sg13g2_dfrbp_1 \shift_storage.storage[1344]$_SDFFE_PN0P_  (.CLK(clknet_leaf_212_clk_p2c),
    .RESET_B(net981),
    .D(_00485_),
    .Q_N(_06316_),
    .Q(\shift_storage.storage [1344]));
 sg13g2_dfrbp_1 \shift_storage.storage[1345]$_SDFFE_PN0P_  (.CLK(clknet_leaf_212_clk_p2c),
    .RESET_B(net982),
    .D(_00486_),
    .Q_N(_06315_),
    .Q(\shift_storage.storage [1345]));
 sg13g2_dfrbp_1 \shift_storage.storage[1346]$_SDFFE_PN0P_  (.CLK(clknet_leaf_213_clk_p2c),
    .RESET_B(net983),
    .D(_00487_),
    .Q_N(_06314_),
    .Q(\shift_storage.storage [1346]));
 sg13g2_dfrbp_1 \shift_storage.storage[1347]$_SDFFE_PN0P_  (.CLK(clknet_leaf_213_clk_p2c),
    .RESET_B(net984),
    .D(_00488_),
    .Q_N(_06313_),
    .Q(\shift_storage.storage [1347]));
 sg13g2_dfrbp_1 \shift_storage.storage[1348]$_SDFFE_PN0P_  (.CLK(clknet_leaf_209_clk_p2c),
    .RESET_B(net985),
    .D(_00489_),
    .Q_N(_06312_),
    .Q(\shift_storage.storage [1348]));
 sg13g2_dfrbp_1 \shift_storage.storage[1349]$_SDFFE_PN0P_  (.CLK(clknet_leaf_211_clk_p2c),
    .RESET_B(net986),
    .D(_00490_),
    .Q_N(_06311_),
    .Q(\shift_storage.storage [1349]));
 sg13g2_dfrbp_1 \shift_storage.storage[134]$_SDFFE_PN0P_  (.CLK(clknet_leaf_212_clk_p2c),
    .RESET_B(net987),
    .D(_00491_),
    .Q_N(_06310_),
    .Q(\shift_storage.storage [134]));
 sg13g2_dfrbp_1 \shift_storage.storage[1350]$_SDFFE_PN0P_  (.CLK(clknet_leaf_211_clk_p2c),
    .RESET_B(net988),
    .D(_00492_),
    .Q_N(_06309_),
    .Q(\shift_storage.storage [1350]));
 sg13g2_dfrbp_1 \shift_storage.storage[1351]$_SDFFE_PN0P_  (.CLK(clknet_leaf_211_clk_p2c),
    .RESET_B(net989),
    .D(_00493_),
    .Q_N(_06308_),
    .Q(\shift_storage.storage [1351]));
 sg13g2_dfrbp_1 \shift_storage.storage[1352]$_SDFFE_PN0P_  (.CLK(clknet_leaf_211_clk_p2c),
    .RESET_B(net990),
    .D(_00494_),
    .Q_N(_06307_),
    .Q(\shift_storage.storage [1352]));
 sg13g2_dfrbp_1 \shift_storage.storage[1353]$_SDFFE_PN0P_  (.CLK(clknet_leaf_178_clk_p2c),
    .RESET_B(net991),
    .D(_00495_),
    .Q_N(_06306_),
    .Q(\shift_storage.storage [1353]));
 sg13g2_dfrbp_1 \shift_storage.storage[1354]$_SDFFE_PN0P_  (.CLK(clknet_leaf_178_clk_p2c),
    .RESET_B(net992),
    .D(_00496_),
    .Q_N(_06305_),
    .Q(\shift_storage.storage [1354]));
 sg13g2_dfrbp_1 \shift_storage.storage[1355]$_SDFFE_PN0P_  (.CLK(clknet_leaf_178_clk_p2c),
    .RESET_B(net993),
    .D(_00497_),
    .Q_N(_06304_),
    .Q(\shift_storage.storage [1355]));
 sg13g2_dfrbp_1 \shift_storage.storage[1356]$_SDFFE_PN0P_  (.CLK(clknet_leaf_178_clk_p2c),
    .RESET_B(net994),
    .D(_00498_),
    .Q_N(_06303_),
    .Q(\shift_storage.storage [1356]));
 sg13g2_dfrbp_1 \shift_storage.storage[1357]$_SDFFE_PN0P_  (.CLK(clknet_leaf_179_clk_p2c),
    .RESET_B(net995),
    .D(_00499_),
    .Q_N(_06302_),
    .Q(\shift_storage.storage [1357]));
 sg13g2_dfrbp_1 \shift_storage.storage[1358]$_SDFFE_PN0P_  (.CLK(clknet_leaf_179_clk_p2c),
    .RESET_B(net996),
    .D(_00500_),
    .Q_N(_06301_),
    .Q(\shift_storage.storage [1358]));
 sg13g2_dfrbp_1 \shift_storage.storage[1359]$_SDFFE_PN0P_  (.CLK(clknet_leaf_187_clk_p2c),
    .RESET_B(net997),
    .D(_00501_),
    .Q_N(_06300_),
    .Q(\shift_storage.storage [1359]));
 sg13g2_dfrbp_1 \shift_storage.storage[135]$_SDFFE_PN0P_  (.CLK(clknet_leaf_211_clk_p2c),
    .RESET_B(net998),
    .D(_00502_),
    .Q_N(_06299_),
    .Q(\shift_storage.storage [135]));
 sg13g2_dfrbp_1 \shift_storage.storage[1360]$_SDFFE_PN0P_  (.CLK(clknet_leaf_198_clk_p2c),
    .RESET_B(net999),
    .D(_00503_),
    .Q_N(_06298_),
    .Q(\shift_storage.storage [1360]));
 sg13g2_dfrbp_1 \shift_storage.storage[1361]$_SDFFE_PN0P_  (.CLK(clknet_leaf_198_clk_p2c),
    .RESET_B(net1000),
    .D(_00504_),
    .Q_N(_06297_),
    .Q(\shift_storage.storage [1361]));
 sg13g2_dfrbp_1 \shift_storage.storage[1362]$_SDFFE_PN0P_  (.CLK(clknet_leaf_211_clk_p2c),
    .RESET_B(net1001),
    .D(_00505_),
    .Q_N(_06296_),
    .Q(\shift_storage.storage [1362]));
 sg13g2_dfrbp_1 \shift_storage.storage[1363]$_SDFFE_PN0P_  (.CLK(clknet_leaf_211_clk_p2c),
    .RESET_B(net1002),
    .D(_00506_),
    .Q_N(_06295_),
    .Q(\shift_storage.storage [1363]));
 sg13g2_dfrbp_1 \shift_storage.storage[1364]$_SDFFE_PN0P_  (.CLK(clknet_leaf_198_clk_p2c),
    .RESET_B(net1003),
    .D(_00507_),
    .Q_N(_06294_),
    .Q(\shift_storage.storage [1364]));
 sg13g2_dfrbp_1 \shift_storage.storage[1365]$_SDFFE_PN0P_  (.CLK(clknet_leaf_198_clk_p2c),
    .RESET_B(net1004),
    .D(_00508_),
    .Q_N(_06293_),
    .Q(\shift_storage.storage [1365]));
 sg13g2_dfrbp_1 \shift_storage.storage[1366]$_SDFFE_PN0P_  (.CLK(clknet_leaf_199_clk_p2c),
    .RESET_B(net1005),
    .D(_00509_),
    .Q_N(_06292_),
    .Q(\shift_storage.storage [1366]));
 sg13g2_dfrbp_1 \shift_storage.storage[1367]$_SDFFE_PN0P_  (.CLK(clknet_leaf_198_clk_p2c),
    .RESET_B(net1006),
    .D(_00510_),
    .Q_N(_06291_),
    .Q(\shift_storage.storage [1367]));
 sg13g2_dfrbp_1 \shift_storage.storage[1368]$_SDFFE_PN0P_  (.CLK(clknet_leaf_197_clk_p2c),
    .RESET_B(net1007),
    .D(_00511_),
    .Q_N(_06290_),
    .Q(\shift_storage.storage [1368]));
 sg13g2_dfrbp_1 \shift_storage.storage[1369]$_SDFFE_PN0P_  (.CLK(clknet_leaf_197_clk_p2c),
    .RESET_B(net1008),
    .D(_00512_),
    .Q_N(_06289_),
    .Q(\shift_storage.storage [1369]));
 sg13g2_dfrbp_1 \shift_storage.storage[136]$_SDFFE_PN0P_  (.CLK(clknet_leaf_197_clk_p2c),
    .RESET_B(net1009),
    .D(_00513_),
    .Q_N(_06288_),
    .Q(\shift_storage.storage [136]));
 sg13g2_dfrbp_1 \shift_storage.storage[1370]$_SDFFE_PN0P_  (.CLK(clknet_leaf_196_clk_p2c),
    .RESET_B(net1010),
    .D(_00514_),
    .Q_N(_06287_),
    .Q(\shift_storage.storage [1370]));
 sg13g2_dfrbp_1 \shift_storage.storage[1371]$_SDFFE_PN0P_  (.CLK(clknet_leaf_196_clk_p2c),
    .RESET_B(net1011),
    .D(_00515_),
    .Q_N(_06286_),
    .Q(\shift_storage.storage [1371]));
 sg13g2_dfrbp_1 \shift_storage.storage[1372]$_SDFFE_PN0P_  (.CLK(clknet_leaf_197_clk_p2c),
    .RESET_B(net1012),
    .D(_00516_),
    .Q_N(_06285_),
    .Q(\shift_storage.storage [1372]));
 sg13g2_dfrbp_1 \shift_storage.storage[1373]$_SDFFE_PN0P_  (.CLK(clknet_leaf_197_clk_p2c),
    .RESET_B(net1013),
    .D(_00517_),
    .Q_N(_06284_),
    .Q(\shift_storage.storage [1373]));
 sg13g2_dfrbp_1 \shift_storage.storage[1374]$_SDFFE_PN0P_  (.CLK(clknet_leaf_198_clk_p2c),
    .RESET_B(net1014),
    .D(_00518_),
    .Q_N(_06283_),
    .Q(\shift_storage.storage [1374]));
 sg13g2_dfrbp_1 \shift_storage.storage[1375]$_SDFFE_PN0P_  (.CLK(clknet_leaf_188_clk_p2c),
    .RESET_B(net1015),
    .D(_00519_),
    .Q_N(_06282_),
    .Q(\shift_storage.storage [1375]));
 sg13g2_dfrbp_1 \shift_storage.storage[1376]$_SDFFE_PN0P_  (.CLK(clknet_leaf_188_clk_p2c),
    .RESET_B(net1016),
    .D(_00520_),
    .Q_N(_06281_),
    .Q(\shift_storage.storage [1376]));
 sg13g2_dfrbp_1 \shift_storage.storage[1377]$_SDFFE_PN0P_  (.CLK(clknet_leaf_188_clk_p2c),
    .RESET_B(net1017),
    .D(_00521_),
    .Q_N(_06280_),
    .Q(\shift_storage.storage [1377]));
 sg13g2_dfrbp_1 \shift_storage.storage[1378]$_SDFFE_PN0P_  (.CLK(clknet_leaf_188_clk_p2c),
    .RESET_B(net1018),
    .D(_00522_),
    .Q_N(_06279_),
    .Q(\shift_storage.storage [1378]));
 sg13g2_dfrbp_1 \shift_storage.storage[1379]$_SDFFE_PN0P_  (.CLK(clknet_leaf_188_clk_p2c),
    .RESET_B(net1019),
    .D(_00523_),
    .Q_N(_06278_),
    .Q(\shift_storage.storage [1379]));
 sg13g2_dfrbp_1 \shift_storage.storage[137]$_SDFFE_PN0P_  (.CLK(clknet_leaf_188_clk_p2c),
    .RESET_B(net1020),
    .D(_00524_),
    .Q_N(_06277_),
    .Q(\shift_storage.storage [137]));
 sg13g2_dfrbp_1 \shift_storage.storage[1380]$_SDFFE_PN0P_  (.CLK(clknet_leaf_187_clk_p2c),
    .RESET_B(net1021),
    .D(_00525_),
    .Q_N(_06276_),
    .Q(\shift_storage.storage [1380]));
 sg13g2_dfrbp_1 \shift_storage.storage[1381]$_SDFFE_PN0P_  (.CLK(clknet_leaf_187_clk_p2c),
    .RESET_B(net1022),
    .D(_00526_),
    .Q_N(_06275_),
    .Q(\shift_storage.storage [1381]));
 sg13g2_dfrbp_1 \shift_storage.storage[1382]$_SDFFE_PN0P_  (.CLK(clknet_leaf_187_clk_p2c),
    .RESET_B(net1023),
    .D(_00527_),
    .Q_N(_06274_),
    .Q(\shift_storage.storage [1382]));
 sg13g2_dfrbp_1 \shift_storage.storage[1383]$_SDFFE_PN0P_  (.CLK(clknet_leaf_187_clk_p2c),
    .RESET_B(net1024),
    .D(_00528_),
    .Q_N(_06273_),
    .Q(\shift_storage.storage [1383]));
 sg13g2_dfrbp_1 \shift_storage.storage[1384]$_SDFFE_PN0P_  (.CLK(clknet_leaf_187_clk_p2c),
    .RESET_B(net1025),
    .D(_00529_),
    .Q_N(_06272_),
    .Q(\shift_storage.storage [1384]));
 sg13g2_dfrbp_1 \shift_storage.storage[1385]$_SDFFE_PN0P_  (.CLK(clknet_leaf_186_clk_p2c),
    .RESET_B(net1026),
    .D(_00530_),
    .Q_N(_06271_),
    .Q(\shift_storage.storage [1385]));
 sg13g2_dfrbp_1 \shift_storage.storage[1386]$_SDFFE_PN0P_  (.CLK(clknet_leaf_179_clk_p2c),
    .RESET_B(net1027),
    .D(_00531_),
    .Q_N(_06270_),
    .Q(\shift_storage.storage [1386]));
 sg13g2_dfrbp_1 \shift_storage.storage[1387]$_SDFFE_PN0P_  (.CLK(clknet_leaf_186_clk_p2c),
    .RESET_B(net1028),
    .D(_00532_),
    .Q_N(_06269_),
    .Q(\shift_storage.storage [1387]));
 sg13g2_dfrbp_1 \shift_storage.storage[1388]$_SDFFE_PN0P_  (.CLK(clknet_leaf_185_clk_p2c),
    .RESET_B(net1029),
    .D(_00533_),
    .Q_N(_06268_),
    .Q(\shift_storage.storage [1388]));
 sg13g2_dfrbp_1 \shift_storage.storage[1389]$_SDFFE_PN0P_  (.CLK(clknet_leaf_186_clk_p2c),
    .RESET_B(net1030),
    .D(_00534_),
    .Q_N(_06267_),
    .Q(\shift_storage.storage [1389]));
 sg13g2_dfrbp_1 \shift_storage.storage[138]$_SDFFE_PN0P_  (.CLK(clknet_leaf_189_clk_p2c),
    .RESET_B(net1031),
    .D(_00535_),
    .Q_N(_06266_),
    .Q(\shift_storage.storage [138]));
 sg13g2_dfrbp_1 \shift_storage.storage[1390]$_SDFFE_PN0P_  (.CLK(clknet_leaf_186_clk_p2c),
    .RESET_B(net1032),
    .D(_00536_),
    .Q_N(_06265_),
    .Q(\shift_storage.storage [1390]));
 sg13g2_dfrbp_1 \shift_storage.storage[1391]$_SDFFE_PN0P_  (.CLK(clknet_leaf_186_clk_p2c),
    .RESET_B(net1033),
    .D(_00537_),
    .Q_N(_06264_),
    .Q(\shift_storage.storage [1391]));
 sg13g2_dfrbp_1 \shift_storage.storage[1392]$_SDFFE_PN0P_  (.CLK(clknet_leaf_186_clk_p2c),
    .RESET_B(net1034),
    .D(_00538_),
    .Q_N(_06263_),
    .Q(\shift_storage.storage [1392]));
 sg13g2_dfrbp_1 \shift_storage.storage[1393]$_SDFFE_PN0P_  (.CLK(clknet_leaf_183_clk_p2c),
    .RESET_B(net1035),
    .D(_00539_),
    .Q_N(_06262_),
    .Q(\shift_storage.storage [1393]));
 sg13g2_dfrbp_1 \shift_storage.storage[1394]$_SDFFE_PN0P_  (.CLK(clknet_leaf_183_clk_p2c),
    .RESET_B(net1036),
    .D(_00540_),
    .Q_N(_06261_),
    .Q(\shift_storage.storage [1394]));
 sg13g2_dfrbp_1 \shift_storage.storage[1395]$_SDFFE_PN0P_  (.CLK(clknet_leaf_184_clk_p2c),
    .RESET_B(net1037),
    .D(_00541_),
    .Q_N(_06260_),
    .Q(\shift_storage.storage [1395]));
 sg13g2_dfrbp_1 \shift_storage.storage[1396]$_SDFFE_PN0P_  (.CLK(clknet_leaf_184_clk_p2c),
    .RESET_B(net1038),
    .D(_00542_),
    .Q_N(_06259_),
    .Q(\shift_storage.storage [1396]));
 sg13g2_dfrbp_1 \shift_storage.storage[1397]$_SDFFE_PN0P_  (.CLK(clknet_leaf_185_clk_p2c),
    .RESET_B(net1039),
    .D(_00543_),
    .Q_N(_06258_),
    .Q(\shift_storage.storage [1397]));
 sg13g2_dfrbp_1 \shift_storage.storage[1398]$_SDFFE_PN0P_  (.CLK(clknet_leaf_185_clk_p2c),
    .RESET_B(net1040),
    .D(_00544_),
    .Q_N(_06257_),
    .Q(\shift_storage.storage [1398]));
 sg13g2_dfrbp_1 \shift_storage.storage[1399]$_SDFFE_PN0P_  (.CLK(clknet_leaf_185_clk_p2c),
    .RESET_B(net1041),
    .D(_00545_),
    .Q_N(_06256_),
    .Q(\shift_storage.storage [1399]));
 sg13g2_dfrbp_1 \shift_storage.storage[139]$_SDFFE_PN0P_  (.CLK(clknet_leaf_189_clk_p2c),
    .RESET_B(net1042),
    .D(_00546_),
    .Q_N(_06255_),
    .Q(\shift_storage.storage [139]));
 sg13g2_dfrbp_1 \shift_storage.storage[13]$_SDFFE_PN0P_  (.CLK(clknet_leaf_184_clk_p2c),
    .RESET_B(net1043),
    .D(_00547_),
    .Q_N(_06254_),
    .Q(\shift_storage.storage [13]));
 sg13g2_dfrbp_1 \shift_storage.storage[1400]$_SDFFE_PN0P_  (.CLK(clknet_leaf_185_clk_p2c),
    .RESET_B(net1044),
    .D(_00548_),
    .Q_N(_06253_),
    .Q(\shift_storage.storage [1400]));
 sg13g2_dfrbp_1 \shift_storage.storage[1401]$_SDFFE_PN0P_  (.CLK(clknet_leaf_190_clk_p2c),
    .RESET_B(net1045),
    .D(_00549_),
    .Q_N(_06252_),
    .Q(\shift_storage.storage [1401]));
 sg13g2_dfrbp_1 \shift_storage.storage[1402]$_SDFFE_PN0P_  (.CLK(clknet_leaf_190_clk_p2c),
    .RESET_B(net1046),
    .D(_00550_),
    .Q_N(_06251_),
    .Q(\shift_storage.storage [1402]));
 sg13g2_dfrbp_1 \shift_storage.storage[1403]$_SDFFE_PN0P_  (.CLK(clknet_leaf_185_clk_p2c),
    .RESET_B(net1047),
    .D(_00551_),
    .Q_N(_06250_),
    .Q(\shift_storage.storage [1403]));
 sg13g2_dfrbp_1 \shift_storage.storage[1404]$_SDFFE_PN0P_  (.CLK(clknet_leaf_185_clk_p2c),
    .RESET_B(net1048),
    .D(_00552_),
    .Q_N(_06249_),
    .Q(\shift_storage.storage [1404]));
 sg13g2_dfrbp_1 \shift_storage.storage[1405]$_SDFFE_PN0P_  (.CLK(clknet_leaf_190_clk_p2c),
    .RESET_B(net1049),
    .D(_00553_),
    .Q_N(_06248_),
    .Q(\shift_storage.storage [1405]));
 sg13g2_dfrbp_1 \shift_storage.storage[1406]$_SDFFE_PN0P_  (.CLK(clknet_leaf_190_clk_p2c),
    .RESET_B(net1050),
    .D(_00554_),
    .Q_N(_06247_),
    .Q(\shift_storage.storage [1406]));
 sg13g2_dfrbp_1 \shift_storage.storage[1407]$_SDFFE_PN0P_  (.CLK(clknet_leaf_190_clk_p2c),
    .RESET_B(net1051),
    .D(_00555_),
    .Q_N(_06246_),
    .Q(\shift_storage.storage [1407]));
 sg13g2_dfrbp_1 \shift_storage.storage[1408]$_SDFFE_PN0P_  (.CLK(clknet_leaf_190_clk_p2c),
    .RESET_B(net1052),
    .D(_00556_),
    .Q_N(_06245_),
    .Q(\shift_storage.storage [1408]));
 sg13g2_dfrbp_1 \shift_storage.storage[1409]$_SDFFE_PN0P_  (.CLK(clknet_leaf_190_clk_p2c),
    .RESET_B(net1053),
    .D(_00557_),
    .Q_N(_06244_),
    .Q(\shift_storage.storage [1409]));
 sg13g2_dfrbp_1 \shift_storage.storage[140]$_SDFFE_PN0P_  (.CLK(clknet_leaf_189_clk_p2c),
    .RESET_B(net1054),
    .D(_00558_),
    .Q_N(_06243_),
    .Q(\shift_storage.storage [140]));
 sg13g2_dfrbp_1 \shift_storage.storage[1410]$_SDFFE_PN0P_  (.CLK(clknet_leaf_191_clk_p2c),
    .RESET_B(net1055),
    .D(_00559_),
    .Q_N(_06242_),
    .Q(\shift_storage.storage [1410]));
 sg13g2_dfrbp_1 \shift_storage.storage[1411]$_SDFFE_PN0P_  (.CLK(clknet_leaf_191_clk_p2c),
    .RESET_B(net1056),
    .D(_00560_),
    .Q_N(_06241_),
    .Q(\shift_storage.storage [1411]));
 sg13g2_dfrbp_1 \shift_storage.storage[1412]$_SDFFE_PN0P_  (.CLK(clknet_leaf_189_clk_p2c),
    .RESET_B(net1057),
    .D(_00561_),
    .Q_N(_06240_),
    .Q(\shift_storage.storage [1412]));
 sg13g2_dfrbp_1 \shift_storage.storage[1413]$_SDFFE_PN0P_  (.CLK(clknet_leaf_189_clk_p2c),
    .RESET_B(net1058),
    .D(_00562_),
    .Q_N(_06239_),
    .Q(\shift_storage.storage [1413]));
 sg13g2_dfrbp_1 \shift_storage.storage[1414]$_SDFFE_PN0P_  (.CLK(clknet_leaf_192_clk_p2c),
    .RESET_B(net1059),
    .D(_00563_),
    .Q_N(_06238_),
    .Q(\shift_storage.storage [1414]));
 sg13g2_dfrbp_1 \shift_storage.storage[1415]$_SDFFE_PN0P_  (.CLK(clknet_leaf_192_clk_p2c),
    .RESET_B(net1060),
    .D(_00564_),
    .Q_N(_06237_),
    .Q(\shift_storage.storage [1415]));
 sg13g2_dfrbp_1 \shift_storage.storage[1416]$_SDFFE_PN0P_  (.CLK(clknet_leaf_189_clk_p2c),
    .RESET_B(net1061),
    .D(_00565_),
    .Q_N(_06236_),
    .Q(\shift_storage.storage [1416]));
 sg13g2_dfrbp_1 \shift_storage.storage[1417]$_SDFFE_PN0P_  (.CLK(clknet_leaf_188_clk_p2c),
    .RESET_B(net1062),
    .D(_00566_),
    .Q_N(_06235_),
    .Q(\shift_storage.storage [1417]));
 sg13g2_dfrbp_1 \shift_storage.storage[1418]$_SDFFE_PN0P_  (.CLK(clknet_leaf_195_clk_p2c),
    .RESET_B(net1063),
    .D(_00567_),
    .Q_N(_06234_),
    .Q(\shift_storage.storage [1418]));
 sg13g2_dfrbp_1 \shift_storage.storage[1419]$_SDFFE_PN0P_  (.CLK(clknet_leaf_197_clk_p2c),
    .RESET_B(net1064),
    .D(_00568_),
    .Q_N(_06233_),
    .Q(\shift_storage.storage [1419]));
 sg13g2_dfrbp_1 \shift_storage.storage[141]$_SDFFE_PN0P_  (.CLK(clknet_leaf_192_clk_p2c),
    .RESET_B(net1065),
    .D(_00569_),
    .Q_N(_06232_),
    .Q(\shift_storage.storage [141]));
 sg13g2_dfrbp_1 \shift_storage.storage[1420]$_SDFFE_PN0P_  (.CLK(clknet_leaf_194_clk_p2c),
    .RESET_B(net1066),
    .D(_00570_),
    .Q_N(_06231_),
    .Q(\shift_storage.storage [1420]));
 sg13g2_dfrbp_1 \shift_storage.storage[1421]$_SDFFE_PN0P_  (.CLK(clknet_leaf_194_clk_p2c),
    .RESET_B(net1067),
    .D(_00571_),
    .Q_N(_06230_),
    .Q(\shift_storage.storage [1421]));
 sg13g2_dfrbp_1 \shift_storage.storage[1422]$_SDFFE_PN0P_  (.CLK(clknet_leaf_192_clk_p2c),
    .RESET_B(net1068),
    .D(_00572_),
    .Q_N(_06229_),
    .Q(\shift_storage.storage [1422]));
 sg13g2_dfrbp_1 \shift_storage.storage[1423]$_SDFFE_PN0P_  (.CLK(clknet_leaf_194_clk_p2c),
    .RESET_B(net1069),
    .D(_00573_),
    .Q_N(_06228_),
    .Q(\shift_storage.storage [1423]));
 sg13g2_dfrbp_1 \shift_storage.storage[1424]$_SDFFE_PN0P_  (.CLK(clknet_leaf_193_clk_p2c),
    .RESET_B(net1070),
    .D(_00574_),
    .Q_N(_06227_),
    .Q(\shift_storage.storage [1424]));
 sg13g2_dfrbp_1 \shift_storage.storage[1425]$_SDFFE_PN0P_  (.CLK(clknet_leaf_193_clk_p2c),
    .RESET_B(net1071),
    .D(_00575_),
    .Q_N(_06226_),
    .Q(\shift_storage.storage [1425]));
 sg13g2_dfrbp_1 \shift_storage.storage[1426]$_SDFFE_PN0P_  (.CLK(clknet_leaf_193_clk_p2c),
    .RESET_B(net1072),
    .D(_00576_),
    .Q_N(_06225_),
    .Q(\shift_storage.storage [1426]));
 sg13g2_dfrbp_1 \shift_storage.storage[1427]$_SDFFE_PN0P_  (.CLK(clknet_leaf_193_clk_p2c),
    .RESET_B(net1073),
    .D(_00577_),
    .Q_N(_06224_),
    .Q(\shift_storage.storage [1427]));
 sg13g2_dfrbp_1 \shift_storage.storage[1428]$_SDFFE_PN0P_  (.CLK(clknet_leaf_192_clk_p2c),
    .RESET_B(net1074),
    .D(_00578_),
    .Q_N(_06223_),
    .Q(\shift_storage.storage [1428]));
 sg13g2_dfrbp_1 \shift_storage.storage[1429]$_SDFFE_PN0P_  (.CLK(clknet_leaf_192_clk_p2c),
    .RESET_B(net1075),
    .D(_00579_),
    .Q_N(_06222_),
    .Q(\shift_storage.storage [1429]));
 sg13g2_dfrbp_1 \shift_storage.storage[142]$_SDFFE_PN0P_  (.CLK(clknet_leaf_191_clk_p2c),
    .RESET_B(net1076),
    .D(_00580_),
    .Q_N(_06221_),
    .Q(\shift_storage.storage [142]));
 sg13g2_dfrbp_1 \shift_storage.storage[1430]$_SDFFE_PN0P_  (.CLK(clknet_leaf_125_clk_p2c),
    .RESET_B(net1077),
    .D(_00581_),
    .Q_N(_06220_),
    .Q(\shift_storage.storage [1430]));
 sg13g2_dfrbp_1 \shift_storage.storage[1431]$_SDFFE_PN0P_  (.CLK(clknet_leaf_125_clk_p2c),
    .RESET_B(net1078),
    .D(_00582_),
    .Q_N(_06219_),
    .Q(\shift_storage.storage [1431]));
 sg13g2_dfrbp_1 \shift_storage.storage[1432]$_SDFFE_PN0P_  (.CLK(clknet_leaf_125_clk_p2c),
    .RESET_B(net1079),
    .D(_00583_),
    .Q_N(_06218_),
    .Q(\shift_storage.storage [1432]));
 sg13g2_dfrbp_1 \shift_storage.storage[1433]$_SDFFE_PN0P_  (.CLK(clknet_leaf_126_clk_p2c),
    .RESET_B(net1080),
    .D(_00584_),
    .Q_N(_06217_),
    .Q(\shift_storage.storage [1433]));
 sg13g2_dfrbp_1 \shift_storage.storage[1434]$_SDFFE_PN0P_  (.CLK(clknet_leaf_126_clk_p2c),
    .RESET_B(net1081),
    .D(_00585_),
    .Q_N(_06216_),
    .Q(\shift_storage.storage [1434]));
 sg13g2_dfrbp_1 \shift_storage.storage[1435]$_SDFFE_PN0P_  (.CLK(clknet_leaf_127_clk_p2c),
    .RESET_B(net1082),
    .D(_00586_),
    .Q_N(_06215_),
    .Q(\shift_storage.storage [1435]));
 sg13g2_dfrbp_1 \shift_storage.storage[1436]$_SDFFE_PN0P_  (.CLK(clknet_leaf_191_clk_p2c),
    .RESET_B(net1083),
    .D(_00587_),
    .Q_N(_06214_),
    .Q(\shift_storage.storage [1436]));
 sg13g2_dfrbp_1 \shift_storage.storage[1437]$_SDFFE_PN0P_  (.CLK(clknet_leaf_191_clk_p2c),
    .RESET_B(net1084),
    .D(_00588_),
    .Q_N(_06213_),
    .Q(\shift_storage.storage [1437]));
 sg13g2_dfrbp_1 \shift_storage.storage[1438]$_SDFFE_PN0P_  (.CLK(clknet_leaf_127_clk_p2c),
    .RESET_B(net1085),
    .D(_00589_),
    .Q_N(_06212_),
    .Q(\shift_storage.storage [1438]));
 sg13g2_dfrbp_1 \shift_storage.storage[1439]$_SDFFE_PN0P_  (.CLK(clknet_leaf_191_clk_p2c),
    .RESET_B(net1086),
    .D(_00590_),
    .Q_N(_06211_),
    .Q(\shift_storage.storage [1439]));
 sg13g2_dfrbp_1 \shift_storage.storage[143]$_SDFFE_PN0P_  (.CLK(clknet_leaf_127_clk_p2c),
    .RESET_B(net1087),
    .D(_00591_),
    .Q_N(_06210_),
    .Q(\shift_storage.storage [143]));
 sg13g2_dfrbp_1 \shift_storage.storage[1440]$_SDFFE_PN0P_  (.CLK(clknet_leaf_127_clk_p2c),
    .RESET_B(net1088),
    .D(_00592_),
    .Q_N(_06209_),
    .Q(\shift_storage.storage [1440]));
 sg13g2_dfrbp_1 \shift_storage.storage[1441]$_SDFFE_PN0P_  (.CLK(clknet_leaf_128_clk_p2c),
    .RESET_B(net1089),
    .D(_00593_),
    .Q_N(_06208_),
    .Q(\shift_storage.storage [1441]));
 sg13g2_dfrbp_1 \shift_storage.storage[1442]$_SDFFE_PN0P_  (.CLK(clknet_leaf_127_clk_p2c),
    .RESET_B(net1090),
    .D(_00594_),
    .Q_N(_06207_),
    .Q(\shift_storage.storage [1442]));
 sg13g2_dfrbp_1 \shift_storage.storage[1443]$_SDFFE_PN0P_  (.CLK(clknet_leaf_128_clk_p2c),
    .RESET_B(net1091),
    .D(_00595_),
    .Q_N(_06206_),
    .Q(\shift_storage.storage [1443]));
 sg13g2_dfrbp_1 \shift_storage.storage[1444]$_SDFFE_PN0P_  (.CLK(clknet_leaf_133_clk_p2c),
    .RESET_B(net1092),
    .D(_00596_),
    .Q_N(_06205_),
    .Q(\shift_storage.storage [1444]));
 sg13g2_dfrbp_1 \shift_storage.storage[1445]$_SDFFE_PN0P_  (.CLK(clknet_leaf_128_clk_p2c),
    .RESET_B(net1093),
    .D(_00597_),
    .Q_N(_06204_),
    .Q(\shift_storage.storage [1445]));
 sg13g2_dfrbp_1 \shift_storage.storage[1446]$_SDFFE_PN0P_  (.CLK(clknet_leaf_128_clk_p2c),
    .RESET_B(net1094),
    .D(_00598_),
    .Q_N(_06203_),
    .Q(\shift_storage.storage [1446]));
 sg13g2_dfrbp_1 \shift_storage.storage[1447]$_SDFFE_PN0P_  (.CLK(clknet_leaf_128_clk_p2c),
    .RESET_B(net1095),
    .D(_00599_),
    .Q_N(_06202_),
    .Q(\shift_storage.storage [1447]));
 sg13g2_dfrbp_1 \shift_storage.storage[1448]$_SDFFE_PN0P_  (.CLK(clknet_leaf_129_clk_p2c),
    .RESET_B(net1096),
    .D(_00600_),
    .Q_N(_06201_),
    .Q(\shift_storage.storage [1448]));
 sg13g2_dfrbp_1 \shift_storage.storage[1449]$_SDFFE_PN0P_  (.CLK(clknet_leaf_129_clk_p2c),
    .RESET_B(net1097),
    .D(_00601_),
    .Q_N(_06200_),
    .Q(\shift_storage.storage [1449]));
 sg13g2_dfrbp_1 \shift_storage.storage[144]$_SDFFE_PN0P_  (.CLK(clknet_leaf_131_clk_p2c),
    .RESET_B(net1098),
    .D(_00602_),
    .Q_N(_06199_),
    .Q(\shift_storage.storage [144]));
 sg13g2_dfrbp_1 \shift_storage.storage[1450]$_SDFFE_PN0P_  (.CLK(clknet_leaf_126_clk_p2c),
    .RESET_B(net1099),
    .D(_00603_),
    .Q_N(_06198_),
    .Q(\shift_storage.storage [1450]));
 sg13g2_dfrbp_1 \shift_storage.storage[1451]$_SDFFE_PN0P_  (.CLK(clknet_leaf_129_clk_p2c),
    .RESET_B(net1100),
    .D(_00604_),
    .Q_N(_06197_),
    .Q(\shift_storage.storage [1451]));
 sg13g2_dfrbp_1 \shift_storage.storage[1452]$_SDFFE_PN0P_  (.CLK(clknet_leaf_126_clk_p2c),
    .RESET_B(net1101),
    .D(_00605_),
    .Q_N(_06196_),
    .Q(\shift_storage.storage [1452]));
 sg13g2_dfrbp_1 \shift_storage.storage[1453]$_SDFFE_PN0P_  (.CLK(clknet_leaf_129_clk_p2c),
    .RESET_B(net1102),
    .D(_00606_),
    .Q_N(_06195_),
    .Q(\shift_storage.storage [1453]));
 sg13g2_dfrbp_1 \shift_storage.storage[1454]$_SDFFE_PN0P_  (.CLK(clknet_leaf_129_clk_p2c),
    .RESET_B(net1103),
    .D(_00607_),
    .Q_N(_06194_),
    .Q(\shift_storage.storage [1454]));
 sg13g2_dfrbp_1 \shift_storage.storage[1455]$_SDFFE_PN0P_  (.CLK(clknet_leaf_130_clk_p2c),
    .RESET_B(net1104),
    .D(_00608_),
    .Q_N(_06193_),
    .Q(\shift_storage.storage [1455]));
 sg13g2_dfrbp_1 \shift_storage.storage[1456]$_SDFFE_PN0P_  (.CLK(clknet_leaf_129_clk_p2c),
    .RESET_B(net1105),
    .D(_00609_),
    .Q_N(_06192_),
    .Q(\shift_storage.storage [1456]));
 sg13g2_dfrbp_1 \shift_storage.storage[1457]$_SDFFE_PN0P_  (.CLK(clknet_leaf_130_clk_p2c),
    .RESET_B(net1106),
    .D(_00610_),
    .Q_N(_06191_),
    .Q(\shift_storage.storage [1457]));
 sg13g2_dfrbp_1 \shift_storage.storage[1458]$_SDFFE_PN0P_  (.CLK(clknet_leaf_130_clk_p2c),
    .RESET_B(net1107),
    .D(_00611_),
    .Q_N(_06190_),
    .Q(\shift_storage.storage [1458]));
 sg13g2_dfrbp_1 \shift_storage.storage[1459]$_SDFFE_PN0P_  (.CLK(clknet_leaf_130_clk_p2c),
    .RESET_B(net1108),
    .D(_00612_),
    .Q_N(_06189_),
    .Q(\shift_storage.storage [1459]));
 sg13g2_dfrbp_1 \shift_storage.storage[145]$_SDFFE_PN0P_  (.CLK(clknet_leaf_131_clk_p2c),
    .RESET_B(net1109),
    .D(_00613_),
    .Q_N(_06188_),
    .Q(\shift_storage.storage [145]));
 sg13g2_dfrbp_1 \shift_storage.storage[1460]$_SDFFE_PN0P_  (.CLK(clknet_leaf_130_clk_p2c),
    .RESET_B(net1110),
    .D(_00614_),
    .Q_N(_06187_),
    .Q(\shift_storage.storage [1460]));
 sg13g2_dfrbp_1 \shift_storage.storage[1461]$_SDFFE_PN0P_  (.CLK(clknet_leaf_119_clk_p2c),
    .RESET_B(net1111),
    .D(_00615_),
    .Q_N(_06186_),
    .Q(\shift_storage.storage [1461]));
 sg13g2_dfrbp_1 \shift_storage.storage[1462]$_SDFFE_PN0P_  (.CLK(clknet_leaf_119_clk_p2c),
    .RESET_B(net1112),
    .D(_00616_),
    .Q_N(_06185_),
    .Q(\shift_storage.storage [1462]));
 sg13g2_dfrbp_1 \shift_storage.storage[1463]$_SDFFE_PN0P_  (.CLK(clknet_leaf_119_clk_p2c),
    .RESET_B(net1113),
    .D(_00617_),
    .Q_N(_06184_),
    .Q(\shift_storage.storage [1463]));
 sg13g2_dfrbp_1 \shift_storage.storage[1464]$_SDFFE_PN0P_  (.CLK(clknet_leaf_118_clk_p2c),
    .RESET_B(net1114),
    .D(_00618_),
    .Q_N(_06183_),
    .Q(\shift_storage.storage [1464]));
 sg13g2_dfrbp_1 \shift_storage.storage[1465]$_SDFFE_PN0P_  (.CLK(clknet_leaf_118_clk_p2c),
    .RESET_B(net1115),
    .D(_00619_),
    .Q_N(_06182_),
    .Q(\shift_storage.storage [1465]));
 sg13g2_dfrbp_1 \shift_storage.storage[1466]$_SDFFE_PN0P_  (.CLK(clknet_leaf_118_clk_p2c),
    .RESET_B(net1116),
    .D(_00620_),
    .Q_N(_06181_),
    .Q(\shift_storage.storage [1466]));
 sg13g2_dfrbp_1 \shift_storage.storage[1467]$_SDFFE_PN0P_  (.CLK(clknet_leaf_119_clk_p2c),
    .RESET_B(net1117),
    .D(_00621_),
    .Q_N(_06180_),
    .Q(\shift_storage.storage [1467]));
 sg13g2_dfrbp_1 \shift_storage.storage[1468]$_SDFFE_PN0P_  (.CLK(clknet_leaf_130_clk_p2c),
    .RESET_B(net1118),
    .D(_00622_),
    .Q_N(_06179_),
    .Q(\shift_storage.storage [1468]));
 sg13g2_dfrbp_1 \shift_storage.storage[1469]$_SDFFE_PN0P_  (.CLK(clknet_leaf_131_clk_p2c),
    .RESET_B(net1119),
    .D(_00623_),
    .Q_N(_06178_),
    .Q(\shift_storage.storage [1469]));
 sg13g2_dfrbp_1 \shift_storage.storage[146]$_SDFFE_PN0P_  (.CLK(clknet_leaf_131_clk_p2c),
    .RESET_B(net1120),
    .D(_00624_),
    .Q_N(_06177_),
    .Q(\shift_storage.storage [146]));
 sg13g2_dfrbp_1 \shift_storage.storage[1470]$_SDFFE_PN0P_  (.CLK(clknet_leaf_131_clk_p2c),
    .RESET_B(net1121),
    .D(_00625_),
    .Q_N(_06176_),
    .Q(\shift_storage.storage [1470]));
 sg13g2_dfrbp_1 \shift_storage.storage[1471]$_SDFFE_PN0P_  (.CLK(clknet_leaf_142_clk_p2c),
    .RESET_B(net1122),
    .D(_00626_),
    .Q_N(_06175_),
    .Q(\shift_storage.storage [1471]));
 sg13g2_dfrbp_1 \shift_storage.storage[1472]$_SDFFE_PN0P_  (.CLK(clknet_leaf_142_clk_p2c),
    .RESET_B(net1123),
    .D(_00627_),
    .Q_N(_06174_),
    .Q(\shift_storage.storage [1472]));
 sg13g2_dfrbp_1 \shift_storage.storage[1473]$_SDFFE_PN0P_  (.CLK(clknet_leaf_142_clk_p2c),
    .RESET_B(net1124),
    .D(_00628_),
    .Q_N(_06173_),
    .Q(\shift_storage.storage [1473]));
 sg13g2_dfrbp_1 \shift_storage.storage[1474]$_SDFFE_PN0P_  (.CLK(clknet_leaf_141_clk_p2c),
    .RESET_B(net1125),
    .D(_00629_),
    .Q_N(_06172_),
    .Q(\shift_storage.storage [1474]));
 sg13g2_dfrbp_1 \shift_storage.storage[1475]$_SDFFE_PN0P_  (.CLK(clknet_leaf_141_clk_p2c),
    .RESET_B(net1126),
    .D(_00630_),
    .Q_N(_06171_),
    .Q(\shift_storage.storage [1475]));
 sg13g2_dfrbp_1 \shift_storage.storage[1476]$_SDFFE_PN0P_  (.CLK(clknet_leaf_141_clk_p2c),
    .RESET_B(net1127),
    .D(_00631_),
    .Q_N(_06170_),
    .Q(\shift_storage.storage [1476]));
 sg13g2_dfrbp_1 \shift_storage.storage[1477]$_SDFFE_PN0P_  (.CLK(clknet_leaf_141_clk_p2c),
    .RESET_B(net1128),
    .D(_00632_),
    .Q_N(_06169_),
    .Q(\shift_storage.storage [1477]));
 sg13g2_dfrbp_1 \shift_storage.storage[1478]$_SDFFE_PN0P_  (.CLK(clknet_leaf_140_clk_p2c),
    .RESET_B(net1129),
    .D(_00633_),
    .Q_N(_06168_),
    .Q(\shift_storage.storage [1478]));
 sg13g2_dfrbp_1 \shift_storage.storage[1479]$_SDFFE_PN0P_  (.CLK(clknet_leaf_140_clk_p2c),
    .RESET_B(net1130),
    .D(_00634_),
    .Q_N(_06167_),
    .Q(\shift_storage.storage [1479]));
 sg13g2_dfrbp_1 \shift_storage.storage[147]$_SDFFE_PN0P_  (.CLK(clknet_leaf_131_clk_p2c),
    .RESET_B(net1131),
    .D(_00635_),
    .Q_N(_06166_),
    .Q(\shift_storage.storage [147]));
 sg13g2_dfrbp_1 \shift_storage.storage[1480]$_SDFFE_PN0P_  (.CLK(clknet_leaf_140_clk_p2c),
    .RESET_B(net1132),
    .D(_00636_),
    .Q_N(_06165_),
    .Q(\shift_storage.storage [1480]));
 sg13g2_dfrbp_1 \shift_storage.storage[1481]$_SDFFE_PN0P_  (.CLK(clknet_leaf_141_clk_p2c),
    .RESET_B(net1133),
    .D(_00637_),
    .Q_N(_06164_),
    .Q(\shift_storage.storage [1481]));
 sg13g2_dfrbp_1 \shift_storage.storage[1482]$_SDFFE_PN0P_  (.CLK(clknet_leaf_139_clk_p2c),
    .RESET_B(net1134),
    .D(_00638_),
    .Q_N(_06163_),
    .Q(\shift_storage.storage [1482]));
 sg13g2_dfrbp_1 \shift_storage.storage[1483]$_SDFFE_PN0P_  (.CLK(clknet_leaf_140_clk_p2c),
    .RESET_B(net1135),
    .D(_00639_),
    .Q_N(_06162_),
    .Q(\shift_storage.storage [1483]));
 sg13g2_dfrbp_1 \shift_storage.storage[1484]$_SDFFE_PN0P_  (.CLK(clknet_leaf_137_clk_p2c),
    .RESET_B(net1136),
    .D(_00640_),
    .Q_N(_06161_),
    .Q(\shift_storage.storage [1484]));
 sg13g2_dfrbp_1 \shift_storage.storage[1485]$_SDFFE_PN0P_  (.CLK(clknet_leaf_140_clk_p2c),
    .RESET_B(net1137),
    .D(_00641_),
    .Q_N(_06160_),
    .Q(\shift_storage.storage [1485]));
 sg13g2_dfrbp_1 \shift_storage.storage[1486]$_SDFFE_PN0P_  (.CLK(clknet_leaf_140_clk_p2c),
    .RESET_B(net1138),
    .D(_00642_),
    .Q_N(_06159_),
    .Q(\shift_storage.storage [1486]));
 sg13g2_dfrbp_1 \shift_storage.storage[1487]$_SDFFE_PN0P_  (.CLK(clknet_leaf_137_clk_p2c),
    .RESET_B(net1139),
    .D(_00643_),
    .Q_N(_06158_),
    .Q(\shift_storage.storage [1487]));
 sg13g2_dfrbp_1 \shift_storage.storage[1488]$_SDFFE_PN0P_  (.CLK(clknet_leaf_134_clk_p2c),
    .RESET_B(net1140),
    .D(_00644_),
    .Q_N(_06157_),
    .Q(\shift_storage.storage [1488]));
 sg13g2_dfrbp_1 \shift_storage.storage[1489]$_SDFFE_PN0P_  (.CLK(clknet_leaf_132_clk_p2c),
    .RESET_B(net1141),
    .D(_00645_),
    .Q_N(_06156_),
    .Q(\shift_storage.storage [1489]));
 sg13g2_dfrbp_1 \shift_storage.storage[148]$_SDFFE_PN0P_  (.CLK(clknet_leaf_134_clk_p2c),
    .RESET_B(net1142),
    .D(_00646_),
    .Q_N(_06155_),
    .Q(\shift_storage.storage [148]));
 sg13g2_dfrbp_1 \shift_storage.storage[1490]$_SDFFE_PN0P_  (.CLK(clknet_leaf_132_clk_p2c),
    .RESET_B(net1143),
    .D(_00647_),
    .Q_N(_06154_),
    .Q(\shift_storage.storage [1490]));
 sg13g2_dfrbp_1 \shift_storage.storage[1491]$_SDFFE_PN0P_  (.CLK(clknet_leaf_131_clk_p2c),
    .RESET_B(net1144),
    .D(_00648_),
    .Q_N(_06153_),
    .Q(\shift_storage.storage [1491]));
 sg13g2_dfrbp_1 \shift_storage.storage[1492]$_SDFFE_PN0P_  (.CLK(clknet_leaf_132_clk_p2c),
    .RESET_B(net1145),
    .D(_00649_),
    .Q_N(_06152_),
    .Q(\shift_storage.storage [1492]));
 sg13g2_dfrbp_1 \shift_storage.storage[1493]$_SDFFE_PN0P_  (.CLK(clknet_leaf_132_clk_p2c),
    .RESET_B(net1146),
    .D(_00650_),
    .Q_N(_06151_),
    .Q(\shift_storage.storage [1493]));
 sg13g2_dfrbp_1 \shift_storage.storage[1494]$_SDFFE_PN0P_  (.CLK(clknet_leaf_132_clk_p2c),
    .RESET_B(net1147),
    .D(_00651_),
    .Q_N(_06150_),
    .Q(\shift_storage.storage [1494]));
 sg13g2_dfrbp_1 \shift_storage.storage[1495]$_SDFFE_PN0P_  (.CLK(clknet_leaf_133_clk_p2c),
    .RESET_B(net1148),
    .D(_00652_),
    .Q_N(_06149_),
    .Q(\shift_storage.storage [1495]));
 sg13g2_dfrbp_1 \shift_storage.storage[1496]$_SDFFE_PN0P_  (.CLK(clknet_leaf_134_clk_p2c),
    .RESET_B(net1149),
    .D(_00653_),
    .Q_N(_06148_),
    .Q(\shift_storage.storage [1496]));
 sg13g2_dfrbp_1 \shift_storage.storage[1497]$_SDFFE_PN0P_  (.CLK(clknet_leaf_133_clk_p2c),
    .RESET_B(net1150),
    .D(_00654_),
    .Q_N(_06147_),
    .Q(\shift_storage.storage [1497]));
 sg13g2_dfrbp_1 \shift_storage.storage[1498]$_SDFFE_PN0P_  (.CLK(clknet_leaf_133_clk_p2c),
    .RESET_B(net1151),
    .D(_00655_),
    .Q_N(_06146_),
    .Q(\shift_storage.storage [1498]));
 sg13g2_dfrbp_1 \shift_storage.storage[1499]$_SDFFE_PN0P_  (.CLK(clknet_leaf_133_clk_p2c),
    .RESET_B(net1152),
    .D(_00656_),
    .Q_N(_06145_),
    .Q(\shift_storage.storage [1499]));
 sg13g2_dfrbp_1 \shift_storage.storage[149]$_SDFFE_PN0P_  (.CLK(clknet_leaf_134_clk_p2c),
    .RESET_B(net1153),
    .D(_00657_),
    .Q_N(_06144_),
    .Q(\shift_storage.storage [149]));
 sg13g2_dfrbp_1 \shift_storage.storage[14]$_SDFFE_PN0P_  (.CLK(clknet_leaf_134_clk_p2c),
    .RESET_B(net1154),
    .D(_00658_),
    .Q_N(_06143_),
    .Q(\shift_storage.storage [14]));
 sg13g2_dfrbp_1 \shift_storage.storage[1500]$_SDFFE_PN0P_  (.CLK(clknet_leaf_184_clk_p2c),
    .RESET_B(net1155),
    .D(_00659_),
    .Q_N(_06142_),
    .Q(\shift_storage.storage [1500]));
 sg13g2_dfrbp_1 \shift_storage.storage[1501]$_SDFFE_PN0P_  (.CLK(clknet_leaf_184_clk_p2c),
    .RESET_B(net1156),
    .D(_00660_),
    .Q_N(_06141_),
    .Q(\shift_storage.storage [1501]));
 sg13g2_dfrbp_1 \shift_storage.storage[1502]$_SDFFE_PN0P_  (.CLK(clknet_leaf_133_clk_p2c),
    .RESET_B(net1157),
    .D(_00661_),
    .Q_N(_06140_),
    .Q(\shift_storage.storage [1502]));
 sg13g2_dfrbp_1 \shift_storage.storage[1503]$_SDFFE_PN0P_  (.CLK(clknet_leaf_134_clk_p2c),
    .RESET_B(net1158),
    .D(_00662_),
    .Q_N(_06139_),
    .Q(\shift_storage.storage [1503]));
 sg13g2_dfrbp_1 \shift_storage.storage[1504]$_SDFFE_PN0P_  (.CLK(clknet_leaf_184_clk_p2c),
    .RESET_B(net1159),
    .D(_00663_),
    .Q_N(_06138_),
    .Q(\shift_storage.storage [1504]));
 sg13g2_dfrbp_1 \shift_storage.storage[1505]$_SDFFE_PN0P_  (.CLK(clknet_leaf_183_clk_p2c),
    .RESET_B(net1160),
    .D(_00664_),
    .Q_N(_06137_),
    .Q(\shift_storage.storage [1505]));
 sg13g2_dfrbp_1 \shift_storage.storage[1506]$_SDFFE_PN0P_  (.CLK(clknet_leaf_184_clk_p2c),
    .RESET_B(net1161),
    .D(_00665_),
    .Q_N(_06136_),
    .Q(\shift_storage.storage [1506]));
 sg13g2_dfrbp_1 \shift_storage.storage[1507]$_SDFFE_PN0P_  (.CLK(clknet_leaf_183_clk_p2c),
    .RESET_B(net1162),
    .D(_00666_),
    .Q_N(_06135_),
    .Q(\shift_storage.storage [1507]));
 sg13g2_dfrbp_1 \shift_storage.storage[1508]$_SDFFE_PN0P_  (.CLK(clknet_leaf_183_clk_p2c),
    .RESET_B(net1163),
    .D(_00667_),
    .Q_N(_06134_),
    .Q(\shift_storage.storage [1508]));
 sg13g2_dfrbp_1 \shift_storage.storage[1509]$_SDFFE_PN0P_  (.CLK(clknet_leaf_183_clk_p2c),
    .RESET_B(net1164),
    .D(_00668_),
    .Q_N(_06133_),
    .Q(\shift_storage.storage [1509]));
 sg13g2_dfrbp_1 \shift_storage.storage[150]$_SDFFE_PN0P_  (.CLK(clknet_leaf_134_clk_p2c),
    .RESET_B(net1165),
    .D(_00669_),
    .Q_N(_06132_),
    .Q(\shift_storage.storage [150]));
 sg13g2_dfrbp_1 \shift_storage.storage[1510]$_SDFFE_PN0P_  (.CLK(clknet_leaf_182_clk_p2c),
    .RESET_B(net1166),
    .D(_00670_),
    .Q_N(_06131_),
    .Q(\shift_storage.storage [1510]));
 sg13g2_dfrbp_1 \shift_storage.storage[1511]$_SDFFE_PN0P_  (.CLK(clknet_leaf_135_clk_p2c),
    .RESET_B(net1167),
    .D(_00671_),
    .Q_N(_06130_),
    .Q(\shift_storage.storage [1511]));
 sg13g2_dfrbp_1 \shift_storage.storage[1512]$_SDFFE_PN0P_  (.CLK(clknet_leaf_135_clk_p2c),
    .RESET_B(net1168),
    .D(_00672_),
    .Q_N(_06129_),
    .Q(\shift_storage.storage [1512]));
 sg13g2_dfrbp_1 \shift_storage.storage[1513]$_SDFFE_PN0P_  (.CLK(clknet_leaf_135_clk_p2c),
    .RESET_B(net1169),
    .D(_00673_),
    .Q_N(_06128_),
    .Q(\shift_storage.storage [1513]));
 sg13g2_dfrbp_1 \shift_storage.storage[1514]$_SDFFE_PN0P_  (.CLK(clknet_leaf_136_clk_p2c),
    .RESET_B(net1170),
    .D(_00674_),
    .Q_N(_06127_),
    .Q(\shift_storage.storage [1514]));
 sg13g2_dfrbp_1 \shift_storage.storage[1515]$_SDFFE_PN0P_  (.CLK(clknet_leaf_135_clk_p2c),
    .RESET_B(net1171),
    .D(_00675_),
    .Q_N(_06126_),
    .Q(\shift_storage.storage [1515]));
 sg13g2_dfrbp_1 \shift_storage.storage[1516]$_SDFFE_PN0P_  (.CLK(clknet_leaf_182_clk_p2c),
    .RESET_B(net1172),
    .D(_00676_),
    .Q_N(_06125_),
    .Q(\shift_storage.storage [1516]));
 sg13g2_dfrbp_1 \shift_storage.storage[1517]$_SDFFE_PN0P_  (.CLK(clknet_leaf_135_clk_p2c),
    .RESET_B(net1173),
    .D(_00677_),
    .Q_N(_06124_),
    .Q(\shift_storage.storage [1517]));
 sg13g2_dfrbp_1 \shift_storage.storage[1518]$_SDFFE_PN0P_  (.CLK(clknet_leaf_135_clk_p2c),
    .RESET_B(net1174),
    .D(_00678_),
    .Q_N(_06123_),
    .Q(\shift_storage.storage [1518]));
 sg13g2_dfrbp_1 \shift_storage.storage[1519]$_SDFFE_PN0P_  (.CLK(clknet_leaf_136_clk_p2c),
    .RESET_B(net1175),
    .D(_00679_),
    .Q_N(_06122_),
    .Q(\shift_storage.storage [1519]));
 sg13g2_dfrbp_1 \shift_storage.storage[151]$_SDFFE_PN0P_  (.CLK(clknet_leaf_136_clk_p2c),
    .RESET_B(net1176),
    .D(_00680_),
    .Q_N(_06121_),
    .Q(\shift_storage.storage [151]));
 sg13g2_dfrbp_1 \shift_storage.storage[1520]$_SDFFE_PN0P_  (.CLK(clknet_leaf_160_clk_p2c),
    .RESET_B(net1177),
    .D(_00681_),
    .Q_N(_06120_),
    .Q(\shift_storage.storage [1520]));
 sg13g2_dfrbp_1 \shift_storage.storage[1521]$_SDFFE_PN0P_  (.CLK(clknet_leaf_159_clk_p2c),
    .RESET_B(net1178),
    .D(_00682_),
    .Q_N(_06119_),
    .Q(\shift_storage.storage [1521]));
 sg13g2_dfrbp_1 \shift_storage.storage[1522]$_SDFFE_PN0P_  (.CLK(clknet_leaf_159_clk_p2c),
    .RESET_B(net1179),
    .D(_00683_),
    .Q_N(_06118_),
    .Q(\shift_storage.storage [1522]));
 sg13g2_dfrbp_1 \shift_storage.storage[1523]$_SDFFE_PN0P_  (.CLK(clknet_leaf_159_clk_p2c),
    .RESET_B(net1180),
    .D(_00684_),
    .Q_N(_06117_),
    .Q(\shift_storage.storage [1523]));
 sg13g2_dfrbp_1 \shift_storage.storage[1524]$_SDFFE_PN0P_  (.CLK(clknet_leaf_136_clk_p2c),
    .RESET_B(net1181),
    .D(_00685_),
    .Q_N(_06116_),
    .Q(\shift_storage.storage [1524]));
 sg13g2_dfrbp_1 \shift_storage.storage[1525]$_SDFFE_PN0P_  (.CLK(clknet_leaf_136_clk_p2c),
    .RESET_B(net1182),
    .D(_00686_),
    .Q_N(_06115_),
    .Q(\shift_storage.storage [1525]));
 sg13g2_dfrbp_1 \shift_storage.storage[1526]$_SDFFE_PN0P_  (.CLK(clknet_leaf_136_clk_p2c),
    .RESET_B(net1183),
    .D(_00687_),
    .Q_N(_06114_),
    .Q(\shift_storage.storage [1526]));
 sg13g2_dfrbp_1 \shift_storage.storage[1527]$_SDFFE_PN0P_  (.CLK(clknet_leaf_136_clk_p2c),
    .RESET_B(net1184),
    .D(_00688_),
    .Q_N(_06113_),
    .Q(\shift_storage.storage [1527]));
 sg13g2_dfrbp_1 \shift_storage.storage[1528]$_SDFFE_PN0P_  (.CLK(clknet_leaf_137_clk_p2c),
    .RESET_B(net1185),
    .D(_00689_),
    .Q_N(_06112_),
    .Q(\shift_storage.storage [1528]));
 sg13g2_dfrbp_1 \shift_storage.storage[1529]$_SDFFE_PN0P_  (.CLK(clknet_leaf_137_clk_p2c),
    .RESET_B(net1186),
    .D(_00690_),
    .Q_N(_06111_),
    .Q(\shift_storage.storage [1529]));
 sg13g2_dfrbp_1 \shift_storage.storage[152]$_SDFFE_PN0P_  (.CLK(clknet_leaf_138_clk_p2c),
    .RESET_B(net1187),
    .D(_00691_),
    .Q_N(_06110_),
    .Q(\shift_storage.storage [152]));
 sg13g2_dfrbp_1 \shift_storage.storage[1530]$_SDFFE_PN0P_  (.CLK(clknet_leaf_138_clk_p2c),
    .RESET_B(net1188),
    .D(_00692_),
    .Q_N(_06109_),
    .Q(\shift_storage.storage [1530]));
 sg13g2_dfrbp_1 \shift_storage.storage[1531]$_SDFFE_PN0P_  (.CLK(clknet_leaf_137_clk_p2c),
    .RESET_B(net1189),
    .D(_00693_),
    .Q_N(_06108_),
    .Q(\shift_storage.storage [1531]));
 sg13g2_dfrbp_1 \shift_storage.storage[1532]$_SDFFE_PN0P_  (.CLK(clknet_leaf_137_clk_p2c),
    .RESET_B(net1190),
    .D(_00694_),
    .Q_N(_06107_),
    .Q(\shift_storage.storage [1532]));
 sg13g2_dfrbp_1 \shift_storage.storage[1533]$_SDFFE_PN0P_  (.CLK(clknet_leaf_138_clk_p2c),
    .RESET_B(net1191),
    .D(_00695_),
    .Q_N(_06106_),
    .Q(\shift_storage.storage [1533]));
 sg13g2_dfrbp_1 \shift_storage.storage[1534]$_SDFFE_PN0P_  (.CLK(clknet_leaf_138_clk_p2c),
    .RESET_B(net1192),
    .D(_00696_),
    .Q_N(_06105_),
    .Q(\shift_storage.storage [1534]));
 sg13g2_dfrbp_1 \shift_storage.storage[1535]$_SDFFE_PN0P_  (.CLK(clknet_leaf_138_clk_p2c),
    .RESET_B(net1193),
    .D(_00697_),
    .Q_N(_06104_),
    .Q(\shift_storage.storage [1535]));
 sg13g2_dfrbp_1 \shift_storage.storage[1536]$_SDFFE_PN0P_  (.CLK(clknet_leaf_157_clk_p2c),
    .RESET_B(net1194),
    .D(_00698_),
    .Q_N(_06103_),
    .Q(\shift_storage.storage [1536]));
 sg13g2_dfrbp_1 \shift_storage.storage[1537]$_SDFFE_PN0P_  (.CLK(clknet_leaf_157_clk_p2c),
    .RESET_B(net1195),
    .D(_00699_),
    .Q_N(_06102_),
    .Q(\shift_storage.storage [1537]));
 sg13g2_dfrbp_1 \shift_storage.storage[1538]$_SDFFE_PN0P_  (.CLK(clknet_leaf_158_clk_p2c),
    .RESET_B(net1196),
    .D(_00700_),
    .Q_N(_06101_),
    .Q(\shift_storage.storage [1538]));
 sg13g2_dfrbp_1 \shift_storage.storage[1539]$_SDFFE_PN0P_  (.CLK(clknet_leaf_156_clk_p2c),
    .RESET_B(net1197),
    .D(_00701_),
    .Q_N(_06100_),
    .Q(\shift_storage.storage [1539]));
 sg13g2_dfrbp_1 \shift_storage.storage[153]$_SDFFE_PN0P_  (.CLK(clknet_leaf_157_clk_p2c),
    .RESET_B(net1198),
    .D(_00702_),
    .Q_N(_06099_),
    .Q(\shift_storage.storage [153]));
 sg13g2_dfrbp_1 \shift_storage.storage[1540]$_SDFFE_PN0P_  (.CLK(clknet_leaf_157_clk_p2c),
    .RESET_B(net1199),
    .D(_00703_),
    .Q_N(_06098_),
    .Q(\shift_storage.storage [1540]));
 sg13g2_dfrbp_1 \shift_storage.storage[1541]$_SDFFE_PN0P_  (.CLK(clknet_leaf_156_clk_p2c),
    .RESET_B(net1200),
    .D(_00704_),
    .Q_N(_06097_),
    .Q(\shift_storage.storage [1541]));
 sg13g2_dfrbp_1 \shift_storage.storage[1542]$_SDFFE_PN0P_  (.CLK(clknet_leaf_156_clk_p2c),
    .RESET_B(net1201),
    .D(_00705_),
    .Q_N(_06096_),
    .Q(\shift_storage.storage [1542]));
 sg13g2_dfrbp_1 \shift_storage.storage[1543]$_SDFFE_PN0P_  (.CLK(clknet_leaf_156_clk_p2c),
    .RESET_B(net1202),
    .D(_00706_),
    .Q_N(_06095_),
    .Q(\shift_storage.storage [1543]));
 sg13g2_dfrbp_1 \shift_storage.storage[1544]$_SDFFE_PN0P_  (.CLK(clknet_leaf_156_clk_p2c),
    .RESET_B(net1203),
    .D(_00707_),
    .Q_N(_06094_),
    .Q(\shift_storage.storage [1544]));
 sg13g2_dfrbp_1 \shift_storage.storage[1545]$_SDFFE_PN0P_  (.CLK(clknet_leaf_156_clk_p2c),
    .RESET_B(net1204),
    .D(_00708_),
    .Q_N(_06093_),
    .Q(\shift_storage.storage [1545]));
 sg13g2_dfrbp_1 \shift_storage.storage[1546]$_SDFFE_PN0P_  (.CLK(clknet_leaf_155_clk_p2c),
    .RESET_B(net1205),
    .D(_00709_),
    .Q_N(_06092_),
    .Q(\shift_storage.storage [1546]));
 sg13g2_dfrbp_1 \shift_storage.storage[1547]$_SDFFE_PN0P_  (.CLK(clknet_leaf_155_clk_p2c),
    .RESET_B(net1206),
    .D(_00710_),
    .Q_N(_06091_),
    .Q(\shift_storage.storage [1547]));
 sg13g2_dfrbp_1 \shift_storage.storage[1548]$_SDFFE_PN0P_  (.CLK(clknet_leaf_155_clk_p2c),
    .RESET_B(net1207),
    .D(_00711_),
    .Q_N(_06090_),
    .Q(\shift_storage.storage [1548]));
 sg13g2_dfrbp_1 \shift_storage.storage[1549]$_SDFFE_PN0P_  (.CLK(clknet_leaf_158_clk_p2c),
    .RESET_B(net1208),
    .D(_00712_),
    .Q_N(_06089_),
    .Q(\shift_storage.storage [1549]));
 sg13g2_dfrbp_1 \shift_storage.storage[154]$_SDFFE_PN0P_  (.CLK(clknet_leaf_158_clk_p2c),
    .RESET_B(net1209),
    .D(_00713_),
    .Q_N(_06088_),
    .Q(\shift_storage.storage [154]));
 sg13g2_dfrbp_1 \shift_storage.storage[1550]$_SDFFE_PN0P_  (.CLK(clknet_leaf_158_clk_p2c),
    .RESET_B(net1210),
    .D(_00714_),
    .Q_N(_06087_),
    .Q(\shift_storage.storage [1550]));
 sg13g2_dfrbp_1 \shift_storage.storage[1551]$_SDFFE_PN0P_  (.CLK(clknet_leaf_159_clk_p2c),
    .RESET_B(net1211),
    .D(_00715_),
    .Q_N(_06086_),
    .Q(\shift_storage.storage [1551]));
 sg13g2_dfrbp_1 \shift_storage.storage[1552]$_SDFFE_PN0P_  (.CLK(clknet_leaf_159_clk_p2c),
    .RESET_B(net1212),
    .D(_00716_),
    .Q_N(_06085_),
    .Q(\shift_storage.storage [1552]));
 sg13g2_dfrbp_1 \shift_storage.storage[1553]$_SDFFE_PN0P_  (.CLK(clknet_leaf_158_clk_p2c),
    .RESET_B(net1213),
    .D(_00717_),
    .Q_N(_06084_),
    .Q(\shift_storage.storage [1553]));
 sg13g2_dfrbp_1 \shift_storage.storage[1554]$_SDFFE_PN0P_  (.CLK(clknet_leaf_158_clk_p2c),
    .RESET_B(net1214),
    .D(_00718_),
    .Q_N(_06083_),
    .Q(\shift_storage.storage [1554]));
 sg13g2_dfrbp_1 \shift_storage.storage[1555]$_SDFFE_PN0P_  (.CLK(clknet_leaf_161_clk_p2c),
    .RESET_B(net1215),
    .D(_00719_),
    .Q_N(_06082_),
    .Q(\shift_storage.storage [1555]));
 sg13g2_dfrbp_1 \shift_storage.storage[1556]$_SDFFE_PN0P_  (.CLK(clknet_leaf_161_clk_p2c),
    .RESET_B(net1216),
    .D(_00720_),
    .Q_N(_06081_),
    .Q(\shift_storage.storage [1556]));
 sg13g2_dfrbp_1 \shift_storage.storage[1557]$_SDFFE_PN0P_  (.CLK(clknet_leaf_161_clk_p2c),
    .RESET_B(net1217),
    .D(_00721_),
    .Q_N(_06080_),
    .Q(\shift_storage.storage [1557]));
 sg13g2_dfrbp_1 \shift_storage.storage[1558]$_SDFFE_PN0P_  (.CLK(clknet_leaf_161_clk_p2c),
    .RESET_B(net1218),
    .D(_00722_),
    .Q_N(_06079_),
    .Q(\shift_storage.storage [1558]));
 sg13g2_dfrbp_1 \shift_storage.storage[1559]$_SDFFE_PN0P_  (.CLK(clknet_leaf_164_clk_p2c),
    .RESET_B(net1219),
    .D(_00723_),
    .Q_N(_06078_),
    .Q(\shift_storage.storage [1559]));
 sg13g2_dfrbp_1 \shift_storage.storage[155]$_SDFFE_PN0P_  (.CLK(clknet_leaf_164_clk_p2c),
    .RESET_B(net1220),
    .D(_00724_),
    .Q_N(_06077_),
    .Q(\shift_storage.storage [155]));
 sg13g2_dfrbp_1 \shift_storage.storage[1560]$_SDFFE_PN0P_  (.CLK(clknet_leaf_164_clk_p2c),
    .RESET_B(net1221),
    .D(_00725_),
    .Q_N(_06076_),
    .Q(\shift_storage.storage [1560]));
 sg13g2_dfrbp_1 \shift_storage.storage[1561]$_SDFFE_PN0P_  (.CLK(clknet_leaf_164_clk_p2c),
    .RESET_B(net1222),
    .D(_00726_),
    .Q_N(_06075_),
    .Q(\shift_storage.storage [1561]));
 sg13g2_dfrbp_1 \shift_storage.storage[1562]$_SDFFE_PN0P_  (.CLK(clknet_leaf_164_clk_p2c),
    .RESET_B(net1223),
    .D(_00727_),
    .Q_N(_06074_),
    .Q(\shift_storage.storage [1562]));
 sg13g2_dfrbp_1 \shift_storage.storage[1563]$_SDFFE_PN0P_  (.CLK(clknet_leaf_162_clk_p2c),
    .RESET_B(net1224),
    .D(_00728_),
    .Q_N(_06073_),
    .Q(\shift_storage.storage [1563]));
 sg13g2_dfrbp_1 \shift_storage.storage[1564]$_SDFFE_PN0P_  (.CLK(clknet_leaf_162_clk_p2c),
    .RESET_B(net1225),
    .D(_00729_),
    .Q_N(_06072_),
    .Q(\shift_storage.storage [1564]));
 sg13g2_dfrbp_1 \shift_storage.storage[1565]$_SDFFE_PN0P_  (.CLK(clknet_leaf_163_clk_p2c),
    .RESET_B(net1226),
    .D(_00730_),
    .Q_N(_06071_),
    .Q(\shift_storage.storage [1565]));
 sg13g2_dfrbp_1 \shift_storage.storage[1566]$_SDFFE_PN0P_  (.CLK(clknet_leaf_163_clk_p2c),
    .RESET_B(net1227),
    .D(_00731_),
    .Q_N(_06070_),
    .Q(\shift_storage.storage [1566]));
 sg13g2_dfrbp_1 \shift_storage.storage[1567]$_SDFFE_PN0P_  (.CLK(clknet_leaf_163_clk_p2c),
    .RESET_B(net1228),
    .D(_00732_),
    .Q_N(_06069_),
    .Q(\shift_storage.storage [1567]));
 sg13g2_dfrbp_1 \shift_storage.storage[1568]$_SDFFE_PN0P_  (.CLK(clknet_leaf_163_clk_p2c),
    .RESET_B(net1229),
    .D(_00733_),
    .Q_N(_06068_),
    .Q(\shift_storage.storage [1568]));
 sg13g2_dfrbp_1 \shift_storage.storage[1569]$_SDFFE_PN0P_  (.CLK(clknet_leaf_168_clk_p2c),
    .RESET_B(net1230),
    .D(_00734_),
    .Q_N(_06067_),
    .Q(\shift_storage.storage [1569]));
 sg13g2_dfrbp_1 \shift_storage.storage[156]$_SDFFE_PN0P_  (.CLK(clknet_leaf_165_clk_p2c),
    .RESET_B(net1231),
    .D(_00735_),
    .Q_N(_06066_),
    .Q(\shift_storage.storage [156]));
 sg13g2_dfrbp_1 \shift_storage.storage[1570]$_SDFFE_PN0P_  (.CLK(clknet_leaf_163_clk_p2c),
    .RESET_B(net1232),
    .D(_00736_),
    .Q_N(_06065_),
    .Q(\shift_storage.storage [1570]));
 sg13g2_dfrbp_1 \shift_storage.storage[1571]$_SDFFE_PN0P_  (.CLK(clknet_leaf_163_clk_p2c),
    .RESET_B(net1233),
    .D(_00737_),
    .Q_N(_06064_),
    .Q(\shift_storage.storage [1571]));
 sg13g2_dfrbp_1 \shift_storage.storage[1572]$_SDFFE_PN0P_  (.CLK(clknet_leaf_165_clk_p2c),
    .RESET_B(net1234),
    .D(_00738_),
    .Q_N(_06063_),
    .Q(\shift_storage.storage [1572]));
 sg13g2_dfrbp_1 \shift_storage.storage[1573]$_SDFFE_PN0P_  (.CLK(clknet_leaf_165_clk_p2c),
    .RESET_B(net1235),
    .D(_00739_),
    .Q_N(_06062_),
    .Q(\shift_storage.storage [1573]));
 sg13g2_dfrbp_1 \shift_storage.storage[1574]$_SDFFE_PN0P_  (.CLK(clknet_leaf_165_clk_p2c),
    .RESET_B(net1236),
    .D(_00740_),
    .Q_N(_06061_),
    .Q(\shift_storage.storage [1574]));
 sg13g2_dfrbp_1 \shift_storage.storage[1575]$_SDFFE_PN0P_  (.CLK(clknet_leaf_167_clk_p2c),
    .RESET_B(net1237),
    .D(_00741_),
    .Q_N(_06060_),
    .Q(\shift_storage.storage [1575]));
 sg13g2_dfrbp_1 \shift_storage.storage[1576]$_SDFFE_PN0P_  (.CLK(clknet_leaf_167_clk_p2c),
    .RESET_B(net1238),
    .D(_00742_),
    .Q_N(_06059_),
    .Q(\shift_storage.storage [1576]));
 sg13g2_dfrbp_1 \shift_storage.storage[1577]$_SDFFE_PN0P_  (.CLK(clknet_leaf_167_clk_p2c),
    .RESET_B(net1239),
    .D(_00743_),
    .Q_N(_06058_),
    .Q(\shift_storage.storage [1577]));
 sg13g2_dfrbp_1 \shift_storage.storage[1578]$_SDFFE_PN0P_  (.CLK(clknet_leaf_167_clk_p2c),
    .RESET_B(net1240),
    .D(_00744_),
    .Q_N(_06057_),
    .Q(\shift_storage.storage [1578]));
 sg13g2_dfrbp_1 \shift_storage.storage[1579]$_SDFFE_PN0P_  (.CLK(clknet_leaf_167_clk_p2c),
    .RESET_B(net1241),
    .D(_00745_),
    .Q_N(_06056_),
    .Q(\shift_storage.storage [1579]));
 sg13g2_dfrbp_1 \shift_storage.storage[157]$_SDFFE_PN0P_  (.CLK(clknet_leaf_165_clk_p2c),
    .RESET_B(net1242),
    .D(_00746_),
    .Q_N(_06055_),
    .Q(\shift_storage.storage [157]));
 sg13g2_dfrbp_1 \shift_storage.storage[1580]$_SDFFE_PN0P_  (.CLK(clknet_leaf_166_clk_p2c),
    .RESET_B(net1243),
    .D(_00747_),
    .Q_N(_06054_),
    .Q(\shift_storage.storage [1580]));
 sg13g2_dfrbp_1 \shift_storage.storage[1581]$_SDFFE_PN0P_  (.CLK(clknet_leaf_166_clk_p2c),
    .RESET_B(net1244),
    .D(_00748_),
    .Q_N(_06053_),
    .Q(\shift_storage.storage [1581]));
 sg13g2_dfrbp_1 \shift_storage.storage[1582]$_SDFFE_PN0P_  (.CLK(clknet_leaf_166_clk_p2c),
    .RESET_B(net1245),
    .D(_00749_),
    .Q_N(_06052_),
    .Q(\shift_storage.storage [1582]));
 sg13g2_dfrbp_1 \shift_storage.storage[1583]$_SDFFE_PN0P_  (.CLK(clknet_leaf_166_clk_p2c),
    .RESET_B(net1246),
    .D(_00750_),
    .Q_N(_06051_),
    .Q(\shift_storage.storage [1583]));
 sg13g2_dfrbp_1 \shift_storage.storage[1584]$_SDFFE_PN0P_  (.CLK(clknet_leaf_166_clk_p2c),
    .RESET_B(net1247),
    .D(_00751_),
    .Q_N(_06050_),
    .Q(\shift_storage.storage [1584]));
 sg13g2_dfrbp_1 \shift_storage.storage[1585]$_SDFFE_PN0P_  (.CLK(clknet_leaf_166_clk_p2c),
    .RESET_B(net1248),
    .D(_00752_),
    .Q_N(_06049_),
    .Q(\shift_storage.storage [1585]));
 sg13g2_dfrbp_1 \shift_storage.storage[1586]$_SDFFE_PN0P_  (.CLK(clknet_leaf_154_clk_p2c),
    .RESET_B(net1249),
    .D(_00753_),
    .Q_N(_06048_),
    .Q(\shift_storage.storage [1586]));
 sg13g2_dfrbp_1 \shift_storage.storage[1587]$_SDFFE_PN0P_  (.CLK(clknet_leaf_154_clk_p2c),
    .RESET_B(net1250),
    .D(_00754_),
    .Q_N(_06047_),
    .Q(\shift_storage.storage [1587]));
 sg13g2_dfrbp_1 \shift_storage.storage[1588]$_SDFFE_PN0P_  (.CLK(clknet_leaf_154_clk_p2c),
    .RESET_B(net1251),
    .D(_00755_),
    .Q_N(_06046_),
    .Q(\shift_storage.storage [1588]));
 sg13g2_dfrbp_1 \shift_storage.storage[1589]$_SDFFE_PN0P_  (.CLK(clknet_leaf_154_clk_p2c),
    .RESET_B(net1252),
    .D(_00756_),
    .Q_N(_06045_),
    .Q(\shift_storage.storage [1589]));
 sg13g2_dfrbp_1 \shift_storage.storage[158]$_SDFFE_PN0P_  (.CLK(clknet_leaf_165_clk_p2c),
    .RESET_B(net1253),
    .D(_00757_),
    .Q_N(_06044_),
    .Q(\shift_storage.storage [158]));
 sg13g2_dfrbp_1 \shift_storage.storage[1590]$_SDFFE_PN0P_  (.CLK(clknet_leaf_155_clk_p2c),
    .RESET_B(net1254),
    .D(_00758_),
    .Q_N(_06043_),
    .Q(\shift_storage.storage [1590]));
 sg13g2_dfrbp_1 \shift_storage.storage[1591]$_SDFFE_PN0P_  (.CLK(clknet_leaf_155_clk_p2c),
    .RESET_B(net1255),
    .D(_00759_),
    .Q_N(_06042_),
    .Q(\shift_storage.storage [1591]));
 sg13g2_dfrbp_1 \shift_storage.storage[1592]$_SDFFE_PN0P_  (.CLK(clknet_leaf_154_clk_p2c),
    .RESET_B(net1256),
    .D(_00760_),
    .Q_N(_06041_),
    .Q(\shift_storage.storage [1592]));
 sg13g2_dfrbp_1 \shift_storage.storage[1593]$_SDFFE_PN0P_  (.CLK(clknet_leaf_153_clk_p2c),
    .RESET_B(net1257),
    .D(_00761_),
    .Q_N(_06040_),
    .Q(\shift_storage.storage [1593]));
 sg13g2_dfrbp_1 \shift_storage.storage[1594]$_SDFFE_PN0P_  (.CLK(clknet_leaf_153_clk_p2c),
    .RESET_B(net1258),
    .D(_00762_),
    .Q_N(_06039_),
    .Q(\shift_storage.storage [1594]));
 sg13g2_dfrbp_1 \shift_storage.storage[1595]$_SDFFE_PN0P_  (.CLK(clknet_leaf_153_clk_p2c),
    .RESET_B(net1259),
    .D(_00763_),
    .Q_N(_06038_),
    .Q(\shift_storage.storage [1595]));
 sg13g2_dfrbp_1 \shift_storage.storage[1596]$_SDFFE_PN0P_  (.CLK(clknet_leaf_152_clk_p2c),
    .RESET_B(net1260),
    .D(_00764_),
    .Q_N(_06037_),
    .Q(\shift_storage.storage [1596]));
 sg13g2_dfrbp_1 \shift_storage.storage[1597]$_SDFFE_PN0P_  (.CLK(clknet_leaf_152_clk_p2c),
    .RESET_B(net1261),
    .D(_00765_),
    .Q_N(_06036_),
    .Q(\shift_storage.storage [1597]));
 sg13g2_dfrbp_1 \shift_storage.storage[1598]$_SDFFE_PN0P_  (.CLK(clknet_leaf_153_clk_p2c),
    .RESET_B(net1262),
    .D(_00766_),
    .Q_N(_06035_),
    .Q(\shift_storage.storage [1598]));
 sg13g2_dfrbp_1 \shift_storage.storage[1599]$_SDFFE_PN0P_  (.CLK(clknet_leaf_153_clk_p2c),
    .RESET_B(net1263),
    .D(_00767_),
    .Q_N(_06034_),
    .Q(\shift_storage.shreg_out ));
 sg13g2_dfrbp_1 \shift_storage.storage[159]$_SDFFE_PN0P_  (.CLK(clknet_leaf_152_clk_p2c),
    .RESET_B(net1264),
    .D(_00768_),
    .Q_N(_06033_),
    .Q(\shift_storage.storage [159]));
 sg13g2_dfrbp_1 \shift_storage.storage[15]$_SDFFE_PN0P_  (.CLK(clknet_leaf_151_clk_p2c),
    .RESET_B(net1265),
    .D(_00769_),
    .Q_N(_06032_),
    .Q(\shift_storage.storage [15]));
 sg13g2_dfrbp_1 \shift_storage.storage[160]$_SDFFE_PN0P_  (.CLK(clknet_leaf_152_clk_p2c),
    .RESET_B(net1266),
    .D(_00770_),
    .Q_N(_06031_),
    .Q(\shift_storage.storage [160]));
 sg13g2_dfrbp_1 \shift_storage.storage[161]$_SDFFE_PN0P_  (.CLK(clknet_leaf_152_clk_p2c),
    .RESET_B(net1267),
    .D(_00771_),
    .Q_N(_06030_),
    .Q(\shift_storage.storage [161]));
 sg13g2_dfrbp_1 \shift_storage.storage[162]$_SDFFE_PN0P_  (.CLK(clknet_leaf_152_clk_p2c),
    .RESET_B(net1268),
    .D(_00772_),
    .Q_N(_06029_),
    .Q(\shift_storage.storage [162]));
 sg13g2_dfrbp_1 \shift_storage.storage[163]$_SDFFE_PN0P_  (.CLK(clknet_leaf_153_clk_p2c),
    .RESET_B(net1269),
    .D(_00773_),
    .Q_N(_06028_),
    .Q(\shift_storage.storage [163]));
 sg13g2_dfrbp_1 \shift_storage.storage[164]$_SDFFE_PN0P_  (.CLK(clknet_leaf_152_clk_p2c),
    .RESET_B(net1270),
    .D(_00774_),
    .Q_N(_06027_),
    .Q(\shift_storage.storage [164]));
 sg13g2_dfrbp_1 \shift_storage.storage[165]$_SDFFE_PN0P_  (.CLK(clknet_leaf_149_clk_p2c),
    .RESET_B(net1271),
    .D(_00775_),
    .Q_N(_06026_),
    .Q(\shift_storage.storage [165]));
 sg13g2_dfrbp_1 \shift_storage.storage[166]$_SDFFE_PN0P_  (.CLK(clknet_leaf_149_clk_p2c),
    .RESET_B(net1272),
    .D(_00776_),
    .Q_N(_06025_),
    .Q(\shift_storage.storage [166]));
 sg13g2_dfrbp_1 \shift_storage.storage[167]$_SDFFE_PN0P_  (.CLK(clknet_leaf_149_clk_p2c),
    .RESET_B(net1273),
    .D(_00777_),
    .Q_N(_06024_),
    .Q(\shift_storage.storage [167]));
 sg13g2_dfrbp_1 \shift_storage.storage[168]$_SDFFE_PN0P_  (.CLK(clknet_leaf_149_clk_p2c),
    .RESET_B(net1274),
    .D(_00778_),
    .Q_N(_06023_),
    .Q(\shift_storage.storage [168]));
 sg13g2_dfrbp_1 \shift_storage.storage[169]$_SDFFE_PN0P_  (.CLK(clknet_leaf_149_clk_p2c),
    .RESET_B(net1275),
    .D(_00779_),
    .Q_N(_06022_),
    .Q(\shift_storage.storage [169]));
 sg13g2_dfrbp_1 \shift_storage.storage[16]$_SDFFE_PN0P_  (.CLK(clknet_leaf_151_clk_p2c),
    .RESET_B(net1276),
    .D(_00780_),
    .Q_N(_06021_),
    .Q(\shift_storage.storage [16]));
 sg13g2_dfrbp_1 \shift_storage.storage[170]$_SDFFE_PN0P_  (.CLK(clknet_leaf_150_clk_p2c),
    .RESET_B(net1277),
    .D(_00781_),
    .Q_N(_06020_),
    .Q(\shift_storage.storage [170]));
 sg13g2_dfrbp_1 \shift_storage.storage[171]$_SDFFE_PN0P_  (.CLK(clknet_leaf_150_clk_p2c),
    .RESET_B(net1278),
    .D(_00782_),
    .Q_N(_06019_),
    .Q(\shift_storage.storage [171]));
 sg13g2_dfrbp_1 \shift_storage.storage[172]$_SDFFE_PN0P_  (.CLK(clknet_leaf_150_clk_p2c),
    .RESET_B(net1279),
    .D(_00783_),
    .Q_N(_06018_),
    .Q(\shift_storage.storage [172]));
 sg13g2_dfrbp_1 \shift_storage.storage[173]$_SDFFE_PN0P_  (.CLK(clknet_leaf_145_clk_p2c),
    .RESET_B(net1280),
    .D(_00784_),
    .Q_N(_06017_),
    .Q(\shift_storage.storage [173]));
 sg13g2_dfrbp_1 \shift_storage.storage[174]$_SDFFE_PN0P_  (.CLK(clknet_leaf_151_clk_p2c),
    .RESET_B(net1281),
    .D(_00785_),
    .Q_N(_06016_),
    .Q(\shift_storage.storage [174]));
 sg13g2_dfrbp_1 \shift_storage.storage[175]$_SDFFE_PN0P_  (.CLK(clknet_leaf_151_clk_p2c),
    .RESET_B(net1282),
    .D(_00786_),
    .Q_N(_06015_),
    .Q(\shift_storage.storage [175]));
 sg13g2_dfrbp_1 \shift_storage.storage[176]$_SDFFE_PN0P_  (.CLK(clknet_leaf_151_clk_p2c),
    .RESET_B(net1283),
    .D(_00787_),
    .Q_N(_06014_),
    .Q(\shift_storage.storage [176]));
 sg13g2_dfrbp_1 \shift_storage.storage[177]$_SDFFE_PN0P_  (.CLK(clknet_leaf_157_clk_p2c),
    .RESET_B(net1284),
    .D(_00788_),
    .Q_N(_06013_),
    .Q(\shift_storage.storage [177]));
 sg13g2_dfrbp_1 \shift_storage.storage[178]$_SDFFE_PN0P_  (.CLK(clknet_leaf_157_clk_p2c),
    .RESET_B(net1285),
    .D(_00789_),
    .Q_N(_06012_),
    .Q(\shift_storage.storage [178]));
 sg13g2_dfrbp_1 \shift_storage.storage[179]$_SDFFE_PN0P_  (.CLK(clknet_leaf_138_clk_p2c),
    .RESET_B(net1286),
    .D(_00790_),
    .Q_N(_06011_),
    .Q(\shift_storage.storage [179]));
 sg13g2_dfrbp_1 \shift_storage.storage[17]$_SDFFE_PN0P_  (.CLK(clknet_leaf_144_clk_p2c),
    .RESET_B(net1287),
    .D(_00791_),
    .Q_N(_06010_),
    .Q(\shift_storage.storage [17]));
 sg13g2_dfrbp_1 \shift_storage.storage[180]$_SDFFE_PN0P_  (.CLK(clknet_leaf_139_clk_p2c),
    .RESET_B(net1288),
    .D(_00792_),
    .Q_N(_06009_),
    .Q(\shift_storage.storage [180]));
 sg13g2_dfrbp_1 \shift_storage.storage[181]$_SDFFE_PN0P_  (.CLK(clknet_leaf_139_clk_p2c),
    .RESET_B(net1289),
    .D(_00793_),
    .Q_N(_06008_),
    .Q(\shift_storage.storage [181]));
 sg13g2_dfrbp_1 \shift_storage.storage[182]$_SDFFE_PN0P_  (.CLK(clknet_leaf_139_clk_p2c),
    .RESET_B(net1290),
    .D(_00794_),
    .Q_N(_06007_),
    .Q(\shift_storage.storage [182]));
 sg13g2_dfrbp_1 \shift_storage.storage[183]$_SDFFE_PN0P_  (.CLK(clknet_leaf_139_clk_p2c),
    .RESET_B(net1291),
    .D(_00795_),
    .Q_N(_06006_),
    .Q(\shift_storage.storage [183]));
 sg13g2_dfrbp_1 \shift_storage.storage[184]$_SDFFE_PN0P_  (.CLK(clknet_leaf_144_clk_p2c),
    .RESET_B(net1292),
    .D(_00796_),
    .Q_N(_06005_),
    .Q(\shift_storage.storage [184]));
 sg13g2_dfrbp_1 \shift_storage.storage[185]$_SDFFE_PN0P_  (.CLK(clknet_leaf_144_clk_p2c),
    .RESET_B(net1293),
    .D(_00797_),
    .Q_N(_06004_),
    .Q(\shift_storage.storage [185]));
 sg13g2_dfrbp_1 \shift_storage.storage[186]$_SDFFE_PN0P_  (.CLK(clknet_leaf_144_clk_p2c),
    .RESET_B(net1294),
    .D(_00798_),
    .Q_N(_06003_),
    .Q(\shift_storage.storage [186]));
 sg13g2_dfrbp_1 \shift_storage.storage[187]$_SDFFE_PN0P_  (.CLK(clknet_leaf_143_clk_p2c),
    .RESET_B(net1295),
    .D(_00799_),
    .Q_N(_06002_),
    .Q(\shift_storage.storage [187]));
 sg13g2_dfrbp_1 \shift_storage.storage[188]$_SDFFE_PN0P_  (.CLK(clknet_leaf_143_clk_p2c),
    .RESET_B(net1296),
    .D(_00800_),
    .Q_N(_06001_),
    .Q(\shift_storage.storage [188]));
 sg13g2_dfrbp_1 \shift_storage.storage[189]$_SDFFE_PN0P_  (.CLK(clknet_leaf_144_clk_p2c),
    .RESET_B(net1297),
    .D(_00801_),
    .Q_N(_06000_),
    .Q(\shift_storage.storage [189]));
 sg13g2_dfrbp_1 \shift_storage.storage[18]$_SDFFE_PN0P_  (.CLK(clknet_leaf_143_clk_p2c),
    .RESET_B(net1298),
    .D(_00802_),
    .Q_N(_05999_),
    .Q(\shift_storage.storage [18]));
 sg13g2_dfrbp_1 \shift_storage.storage[190]$_SDFFE_PN0P_  (.CLK(clknet_leaf_143_clk_p2c),
    .RESET_B(net1299),
    .D(_00803_),
    .Q_N(_05998_),
    .Q(\shift_storage.storage [190]));
 sg13g2_dfrbp_1 \shift_storage.storage[191]$_SDFFE_PN0P_  (.CLK(clknet_leaf_143_clk_p2c),
    .RESET_B(net1300),
    .D(_00804_),
    .Q_N(_05997_),
    .Q(\shift_storage.storage [191]));
 sg13g2_dfrbp_1 \shift_storage.storage[192]$_SDFFE_PN0P_  (.CLK(clknet_leaf_139_clk_p2c),
    .RESET_B(net1301),
    .D(_00805_),
    .Q_N(_05996_),
    .Q(\shift_storage.storage [192]));
 sg13g2_dfrbp_1 \shift_storage.storage[193]$_SDFFE_PN0P_  (.CLK(clknet_leaf_142_clk_p2c),
    .RESET_B(net1302),
    .D(_00806_),
    .Q_N(_05995_),
    .Q(\shift_storage.storage [193]));
 sg13g2_dfrbp_1 \shift_storage.storage[194]$_SDFFE_PN0P_  (.CLK(clknet_leaf_142_clk_p2c),
    .RESET_B(net1303),
    .D(_00807_),
    .Q_N(_05994_),
    .Q(\shift_storage.storage [194]));
 sg13g2_dfrbp_1 \shift_storage.storage[195]$_SDFFE_PN0P_  (.CLK(clknet_leaf_143_clk_p2c),
    .RESET_B(net1304),
    .D(_00808_),
    .Q_N(_05993_),
    .Q(\shift_storage.storage [195]));
 sg13g2_dfrbp_1 \shift_storage.storage[196]$_SDFFE_PN0P_  (.CLK(clknet_leaf_106_clk_p2c),
    .RESET_B(net1305),
    .D(_00809_),
    .Q_N(_05992_),
    .Q(\shift_storage.storage [196]));
 sg13g2_dfrbp_1 \shift_storage.storage[197]$_SDFFE_PN0P_  (.CLK(clknet_leaf_106_clk_p2c),
    .RESET_B(net1306),
    .D(_00810_),
    .Q_N(_05991_),
    .Q(\shift_storage.storage [197]));
 sg13g2_dfrbp_1 \shift_storage.storage[198]$_SDFFE_PN0P_  (.CLK(clknet_leaf_106_clk_p2c),
    .RESET_B(net1307),
    .D(_00811_),
    .Q_N(_05990_),
    .Q(\shift_storage.storage [198]));
 sg13g2_dfrbp_1 \shift_storage.storage[199]$_SDFFE_PN0P_  (.CLK(clknet_leaf_107_clk_p2c),
    .RESET_B(net1308),
    .D(_00812_),
    .Q_N(_05989_),
    .Q(\shift_storage.storage [199]));
 sg13g2_dfrbp_1 \shift_storage.storage[19]$_SDFFE_PN0P_  (.CLK(clknet_leaf_106_clk_p2c),
    .RESET_B(net1309),
    .D(_00813_),
    .Q_N(_05988_),
    .Q(\shift_storage.storage [19]));
 sg13g2_dfrbp_1 \shift_storage.storage[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_107_clk_p2c),
    .RESET_B(net1310),
    .D(_00814_),
    .Q_N(_05987_),
    .Q(\shift_storage.storage [1]));
 sg13g2_dfrbp_1 \shift_storage.storage[200]$_SDFFE_PN0P_  (.CLK(clknet_leaf_107_clk_p2c),
    .RESET_B(net1311),
    .D(_00815_),
    .Q_N(_05986_),
    .Q(\shift_storage.storage [200]));
 sg13g2_dfrbp_1 \shift_storage.storage[201]$_SDFFE_PN0P_  (.CLK(clknet_leaf_107_clk_p2c),
    .RESET_B(net1312),
    .D(_00816_),
    .Q_N(_05985_),
    .Q(\shift_storage.storage [201]));
 sg13g2_dfrbp_1 \shift_storage.storage[202]$_SDFFE_PN0P_  (.CLK(clknet_leaf_107_clk_p2c),
    .RESET_B(net1313),
    .D(_00817_),
    .Q_N(_05984_),
    .Q(\shift_storage.storage [202]));
 sg13g2_dfrbp_1 \shift_storage.storage[203]$_SDFFE_PN0P_  (.CLK(clknet_leaf_107_clk_p2c),
    .RESET_B(net1314),
    .D(_00818_),
    .Q_N(_05983_),
    .Q(\shift_storage.storage [203]));
 sg13g2_dfrbp_1 \shift_storage.storage[204]$_SDFFE_PN0P_  (.CLK(clknet_leaf_106_clk_p2c),
    .RESET_B(net1315),
    .D(_00819_),
    .Q_N(_05982_),
    .Q(\shift_storage.storage [204]));
 sg13g2_dfrbp_1 \shift_storage.storage[205]$_SDFFE_PN0P_  (.CLK(clknet_leaf_106_clk_p2c),
    .RESET_B(net1316),
    .D(_00820_),
    .Q_N(_05981_),
    .Q(\shift_storage.storage [205]));
 sg13g2_dfrbp_1 \shift_storage.storage[206]$_SDFFE_PN0P_  (.CLK(clknet_leaf_105_clk_p2c),
    .RESET_B(net1317),
    .D(_00821_),
    .Q_N(_05980_),
    .Q(\shift_storage.storage [206]));
 sg13g2_dfrbp_1 \shift_storage.storage[207]$_SDFFE_PN0P_  (.CLK(clknet_leaf_105_clk_p2c),
    .RESET_B(net1318),
    .D(_00822_),
    .Q_N(_05979_),
    .Q(\shift_storage.storage [207]));
 sg13g2_dfrbp_1 \shift_storage.storage[208]$_SDFFE_PN0P_  (.CLK(clknet_leaf_105_clk_p2c),
    .RESET_B(net1319),
    .D(_00823_),
    .Q_N(_05978_),
    .Q(\shift_storage.storage [208]));
 sg13g2_dfrbp_1 \shift_storage.storage[209]$_SDFFE_PN0P_  (.CLK(clknet_leaf_105_clk_p2c),
    .RESET_B(net1320),
    .D(_00824_),
    .Q_N(_05977_),
    .Q(\shift_storage.storage [209]));
 sg13g2_dfrbp_1 \shift_storage.storage[20]$_SDFFE_PN0P_  (.CLK(clknet_leaf_105_clk_p2c),
    .RESET_B(net1321),
    .D(_00825_),
    .Q_N(_05976_),
    .Q(\shift_storage.storage [20]));
 sg13g2_dfrbp_1 \shift_storage.storage[210]$_SDFFE_PN0P_  (.CLK(clknet_leaf_104_clk_p2c),
    .RESET_B(net1322),
    .D(_00826_),
    .Q_N(_05975_),
    .Q(\shift_storage.storage [210]));
 sg13g2_dfrbp_1 \shift_storage.storage[211]$_SDFFE_PN0P_  (.CLK(clknet_leaf_105_clk_p2c),
    .RESET_B(net1323),
    .D(_00827_),
    .Q_N(_05974_),
    .Q(\shift_storage.storage [211]));
 sg13g2_dfrbp_1 \shift_storage.storage[212]$_SDFFE_PN0P_  (.CLK(clknet_leaf_103_clk_p2c),
    .RESET_B(net1324),
    .D(_00828_),
    .Q_N(_05973_),
    .Q(\shift_storage.storage [212]));
 sg13g2_dfrbp_1 \shift_storage.storage[213]$_SDFFE_PN0P_  (.CLK(clknet_leaf_103_clk_p2c),
    .RESET_B(net1325),
    .D(_00829_),
    .Q_N(_05972_),
    .Q(\shift_storage.storage [213]));
 sg13g2_dfrbp_1 \shift_storage.storage[214]$_SDFFE_PN0P_  (.CLK(clknet_leaf_103_clk_p2c),
    .RESET_B(net1326),
    .D(_00830_),
    .Q_N(_05971_),
    .Q(\shift_storage.storage [214]));
 sg13g2_dfrbp_1 \shift_storage.storage[215]$_SDFFE_PN0P_  (.CLK(clknet_leaf_103_clk_p2c),
    .RESET_B(net1327),
    .D(_00831_),
    .Q_N(_05970_),
    .Q(\shift_storage.storage [215]));
 sg13g2_dfrbp_1 \shift_storage.storage[216]$_SDFFE_PN0P_  (.CLK(clknet_leaf_103_clk_p2c),
    .RESET_B(net1328),
    .D(_00832_),
    .Q_N(_05969_),
    .Q(\shift_storage.storage [216]));
 sg13g2_dfrbp_1 \shift_storage.storage[217]$_SDFFE_PN0P_  (.CLK(clknet_leaf_102_clk_p2c),
    .RESET_B(net1329),
    .D(_00833_),
    .Q_N(_05968_),
    .Q(\shift_storage.storage [217]));
 sg13g2_dfrbp_1 \shift_storage.storage[218]$_SDFFE_PN0P_  (.CLK(clknet_leaf_102_clk_p2c),
    .RESET_B(net1330),
    .D(_00834_),
    .Q_N(_05967_),
    .Q(\shift_storage.storage [218]));
 sg13g2_dfrbp_1 \shift_storage.storage[219]$_SDFFE_PN0P_  (.CLK(clknet_leaf_102_clk_p2c),
    .RESET_B(net1331),
    .D(_00835_),
    .Q_N(_05966_),
    .Q(\shift_storage.storage [219]));
 sg13g2_dfrbp_1 \shift_storage.storage[21]$_SDFFE_PN0P_  (.CLK(clknet_leaf_102_clk_p2c),
    .RESET_B(net1332),
    .D(_00836_),
    .Q_N(_05965_),
    .Q(\shift_storage.storage [21]));
 sg13g2_dfrbp_1 \shift_storage.storage[220]$_SDFFE_PN0P_  (.CLK(clknet_leaf_103_clk_p2c),
    .RESET_B(net1333),
    .D(_00837_),
    .Q_N(_05964_),
    .Q(\shift_storage.storage [220]));
 sg13g2_dfrbp_1 \shift_storage.storage[221]$_SDFFE_PN0P_  (.CLK(clknet_leaf_103_clk_p2c),
    .RESET_B(net1334),
    .D(_00838_),
    .Q_N(_05963_),
    .Q(\shift_storage.storage [221]));
 sg13g2_dfrbp_1 \shift_storage.storage[222]$_SDFFE_PN0P_  (.CLK(clknet_leaf_106_clk_p2c),
    .RESET_B(net1335),
    .D(_00839_),
    .Q_N(_05962_),
    .Q(\shift_storage.storage [222]));
 sg13g2_dfrbp_1 \shift_storage.storage[223]$_SDFFE_PN0P_  (.CLK(clknet_leaf_146_clk_p2c),
    .RESET_B(net1336),
    .D(_00840_),
    .Q_N(_05961_),
    .Q(\shift_storage.storage [223]));
 sg13g2_dfrbp_1 \shift_storage.storage[224]$_SDFFE_PN0P_  (.CLK(clknet_leaf_146_clk_p2c),
    .RESET_B(net1337),
    .D(_00841_),
    .Q_N(_05960_),
    .Q(\shift_storage.storage [224]));
 sg13g2_dfrbp_1 \shift_storage.storage[225]$_SDFFE_PN0P_  (.CLK(clknet_leaf_146_clk_p2c),
    .RESET_B(net1338),
    .D(_00842_),
    .Q_N(_05959_),
    .Q(\shift_storage.storage [225]));
 sg13g2_dfrbp_1 \shift_storage.storage[226]$_SDFFE_PN0P_  (.CLK(clknet_leaf_143_clk_p2c),
    .RESET_B(net1339),
    .D(_00843_),
    .Q_N(_05958_),
    .Q(\shift_storage.storage [226]));
 sg13g2_dfrbp_1 \shift_storage.storage[227]$_SDFFE_PN0P_  (.CLK(clknet_leaf_146_clk_p2c),
    .RESET_B(net1340),
    .D(_00844_),
    .Q_N(_05957_),
    .Q(\shift_storage.storage [227]));
 sg13g2_dfrbp_1 \shift_storage.storage[228]$_SDFFE_PN0P_  (.CLK(clknet_leaf_145_clk_p2c),
    .RESET_B(net1341),
    .D(_00845_),
    .Q_N(_05956_),
    .Q(\shift_storage.storage [228]));
 sg13g2_dfrbp_1 \shift_storage.storage[229]$_SDFFE_PN0P_  (.CLK(clknet_leaf_145_clk_p2c),
    .RESET_B(net1342),
    .D(_00846_),
    .Q_N(_05955_),
    .Q(\shift_storage.storage [229]));
 sg13g2_dfrbp_1 \shift_storage.storage[22]$_SDFFE_PN0P_  (.CLK(clknet_leaf_146_clk_p2c),
    .RESET_B(net1343),
    .D(_00847_),
    .Q_N(_05954_),
    .Q(\shift_storage.storage [22]));
 sg13g2_dfrbp_1 \shift_storage.storage[230]$_SDFFE_PN0P_  (.CLK(clknet_leaf_145_clk_p2c),
    .RESET_B(net1344),
    .D(_00848_),
    .Q_N(_05953_),
    .Q(\shift_storage.storage [230]));
 sg13g2_dfrbp_1 \shift_storage.storage[231]$_SDFFE_PN0P_  (.CLK(clknet_leaf_145_clk_p2c),
    .RESET_B(net1345),
    .D(_00849_),
    .Q_N(_05952_),
    .Q(\shift_storage.storage [231]));
 sg13g2_dfrbp_1 \shift_storage.storage[232]$_SDFFE_PN0P_  (.CLK(clknet_leaf_145_clk_p2c),
    .RESET_B(net1346),
    .D(_00850_),
    .Q_N(_05951_),
    .Q(\shift_storage.storage [232]));
 sg13g2_dfrbp_1 \shift_storage.storage[233]$_SDFFE_PN0P_  (.CLK(clknet_leaf_150_clk_p2c),
    .RESET_B(net1347),
    .D(_00851_),
    .Q_N(_05950_),
    .Q(\shift_storage.storage [233]));
 sg13g2_dfrbp_1 \shift_storage.storage[234]$_SDFFE_PN0P_  (.CLK(clknet_leaf_150_clk_p2c),
    .RESET_B(net1348),
    .D(_00852_),
    .Q_N(_05949_),
    .Q(\shift_storage.storage [234]));
 sg13g2_dfrbp_1 \shift_storage.storage[235]$_SDFFE_PN0P_  (.CLK(clknet_leaf_150_clk_p2c),
    .RESET_B(net1349),
    .D(_00853_),
    .Q_N(_05948_),
    .Q(\shift_storage.storage [235]));
 sg13g2_dfrbp_1 \shift_storage.storage[236]$_SDFFE_PN0P_  (.CLK(clknet_leaf_148_clk_p2c),
    .RESET_B(net1350),
    .D(_00854_),
    .Q_N(_05947_),
    .Q(\shift_storage.storage [236]));
 sg13g2_dfrbp_1 \shift_storage.storage[237]$_SDFFE_PN0P_  (.CLK(clknet_leaf_148_clk_p2c),
    .RESET_B(net1351),
    .D(_00855_),
    .Q_N(_05946_),
    .Q(\shift_storage.storage [237]));
 sg13g2_dfrbp_1 \shift_storage.storage[238]$_SDFFE_PN0P_  (.CLK(clknet_leaf_149_clk_p2c),
    .RESET_B(net1352),
    .D(_00856_),
    .Q_N(_05945_),
    .Q(\shift_storage.storage [238]));
 sg13g2_dfrbp_1 \shift_storage.storage[239]$_SDFFE_PN0P_  (.CLK(clknet_leaf_148_clk_p2c),
    .RESET_B(net1353),
    .D(_00857_),
    .Q_N(_05944_),
    .Q(\shift_storage.storage [239]));
 sg13g2_dfrbp_1 \shift_storage.storage[23]$_SDFFE_PN0P_  (.CLK(clknet_leaf_147_clk_p2c),
    .RESET_B(net1354),
    .D(_00858_),
    .Q_N(_05943_),
    .Q(\shift_storage.storage [23]));
 sg13g2_dfrbp_1 \shift_storage.storage[240]$_SDFFE_PN0P_  (.CLK(clknet_leaf_148_clk_p2c),
    .RESET_B(net1355),
    .D(_00859_),
    .Q_N(_05942_),
    .Q(\shift_storage.storage [240]));
 sg13g2_dfrbp_1 \shift_storage.storage[241]$_SDFFE_PN0P_  (.CLK(clknet_leaf_148_clk_p2c),
    .RESET_B(net1356),
    .D(_00860_),
    .Q_N(_05941_),
    .Q(\shift_storage.storage [241]));
 sg13g2_dfrbp_1 \shift_storage.storage[242]$_SDFFE_PN0P_  (.CLK(clknet_leaf_148_clk_p2c),
    .RESET_B(net1357),
    .D(_00861_),
    .Q_N(_05940_),
    .Q(\shift_storage.storage [242]));
 sg13g2_dfrbp_1 \shift_storage.storage[243]$_SDFFE_PN0P_  (.CLK(clknet_leaf_147_clk_p2c),
    .RESET_B(net1358),
    .D(_00862_),
    .Q_N(_05939_),
    .Q(\shift_storage.storage [243]));
 sg13g2_dfrbp_1 \shift_storage.storage[244]$_SDFFE_PN0P_  (.CLK(clknet_leaf_147_clk_p2c),
    .RESET_B(net1359),
    .D(_00863_),
    .Q_N(_05938_),
    .Q(\shift_storage.storage [244]));
 sg13g2_dfrbp_1 \shift_storage.storage[245]$_SDFFE_PN0P_  (.CLK(clknet_leaf_101_clk_p2c),
    .RESET_B(net1360),
    .D(_00864_),
    .Q_N(_05937_),
    .Q(\shift_storage.storage [245]));
 sg13g2_dfrbp_1 \shift_storage.storage[246]$_SDFFE_PN0P_  (.CLK(clknet_leaf_147_clk_p2c),
    .RESET_B(net1361),
    .D(_00865_),
    .Q_N(_05936_),
    .Q(\shift_storage.storage [246]));
 sg13g2_dfrbp_1 \shift_storage.storage[247]$_SDFFE_PN0P_  (.CLK(clknet_leaf_148_clk_p2c),
    .RESET_B(net1362),
    .D(_00866_),
    .Q_N(_05935_),
    .Q(\shift_storage.storage [247]));
 sg13g2_dfrbp_1 \shift_storage.storage[248]$_SDFFE_PN0P_  (.CLK(clknet_leaf_147_clk_p2c),
    .RESET_B(net1363),
    .D(_00867_),
    .Q_N(_05934_),
    .Q(\shift_storage.storage [248]));
 sg13g2_dfrbp_1 \shift_storage.storage[249]$_SDFFE_PN0P_  (.CLK(clknet_leaf_147_clk_p2c),
    .RESET_B(net1364),
    .D(_00868_),
    .Q_N(_05933_),
    .Q(\shift_storage.storage [249]));
 sg13g2_dfrbp_1 \shift_storage.storage[24]$_SDFFE_PN0P_  (.CLK(clknet_leaf_101_clk_p2c),
    .RESET_B(net1365),
    .D(_00869_),
    .Q_N(_05932_),
    .Q(\shift_storage.storage [24]));
 sg13g2_dfrbp_1 \shift_storage.storage[250]$_SDFFE_PN0P_  (.CLK(clknet_leaf_101_clk_p2c),
    .RESET_B(net1366),
    .D(_00870_),
    .Q_N(_05931_),
    .Q(\shift_storage.storage [250]));
 sg13g2_dfrbp_1 \shift_storage.storage[251]$_SDFFE_PN0P_  (.CLK(clknet_leaf_101_clk_p2c),
    .RESET_B(net1367),
    .D(_00871_),
    .Q_N(_05930_),
    .Q(\shift_storage.storage [251]));
 sg13g2_dfrbp_1 \shift_storage.storage[252]$_SDFFE_PN0P_  (.CLK(clknet_leaf_101_clk_p2c),
    .RESET_B(net1368),
    .D(_00872_),
    .Q_N(_05929_),
    .Q(\shift_storage.storage [252]));
 sg13g2_dfrbp_1 \shift_storage.storage[253]$_SDFFE_PN0P_  (.CLK(clknet_leaf_100_clk_p2c),
    .RESET_B(net1369),
    .D(_00873_),
    .Q_N(_05928_),
    .Q(\shift_storage.storage [253]));
 sg13g2_dfrbp_1 \shift_storage.storage[254]$_SDFFE_PN0P_  (.CLK(clknet_leaf_100_clk_p2c),
    .RESET_B(net1370),
    .D(_00874_),
    .Q_N(_05927_),
    .Q(\shift_storage.storage [254]));
 sg13g2_dfrbp_1 \shift_storage.storage[255]$_SDFFE_PN0P_  (.CLK(clknet_leaf_100_clk_p2c),
    .RESET_B(net1371),
    .D(_00875_),
    .Q_N(_05926_),
    .Q(\shift_storage.storage [255]));
 sg13g2_dfrbp_1 \shift_storage.storage[256]$_SDFFE_PN0P_  (.CLK(clknet_leaf_101_clk_p2c),
    .RESET_B(net1372),
    .D(_00876_),
    .Q_N(_05925_),
    .Q(\shift_storage.storage [256]));
 sg13g2_dfrbp_1 \shift_storage.storage[257]$_SDFFE_PN0P_  (.CLK(clknet_leaf_101_clk_p2c),
    .RESET_B(net1373),
    .D(_00877_),
    .Q_N(_05924_),
    .Q(\shift_storage.storage [257]));
 sg13g2_dfrbp_1 \shift_storage.storage[258]$_SDFFE_PN0P_  (.CLK(clknet_leaf_102_clk_p2c),
    .RESET_B(net1374),
    .D(_00878_),
    .Q_N(_05923_),
    .Q(\shift_storage.storage [258]));
 sg13g2_dfrbp_1 \shift_storage.storage[259]$_SDFFE_PN0P_  (.CLK(clknet_leaf_99_clk_p2c),
    .RESET_B(net1375),
    .D(_00879_),
    .Q_N(_05922_),
    .Q(\shift_storage.storage [259]));
 sg13g2_dfrbp_1 \shift_storage.storage[25]$_SDFFE_PN0P_  (.CLK(clknet_leaf_99_clk_p2c),
    .RESET_B(net1376),
    .D(_00880_),
    .Q_N(_05921_),
    .Q(\shift_storage.storage [25]));
 sg13g2_dfrbp_1 \shift_storage.storage[260]$_SDFFE_PN0P_  (.CLK(clknet_leaf_99_clk_p2c),
    .RESET_B(net1377),
    .D(_00881_),
    .Q_N(_05920_),
    .Q(\shift_storage.storage [260]));
 sg13g2_dfrbp_1 \shift_storage.storage[261]$_SDFFE_PN0P_  (.CLK(clknet_leaf_100_clk_p2c),
    .RESET_B(net1378),
    .D(_00882_),
    .Q_N(_05919_),
    .Q(\shift_storage.storage [261]));
 sg13g2_dfrbp_1 \shift_storage.storage[262]$_SDFFE_PN0P_  (.CLK(clknet_leaf_100_clk_p2c),
    .RESET_B(net1379),
    .D(_00883_),
    .Q_N(_05918_),
    .Q(\shift_storage.storage [262]));
 sg13g2_dfrbp_1 \shift_storage.storage[263]$_SDFFE_PN0P_  (.CLK(clknet_leaf_100_clk_p2c),
    .RESET_B(net1380),
    .D(_00884_),
    .Q_N(_05917_),
    .Q(\shift_storage.storage [263]));
 sg13g2_dfrbp_1 \shift_storage.storage[264]$_SDFFE_PN0P_  (.CLK(clknet_leaf_97_clk_p2c),
    .RESET_B(net1381),
    .D(_00885_),
    .Q_N(_05916_),
    .Q(\shift_storage.storage [264]));
 sg13g2_dfrbp_1 \shift_storage.storage[265]$_SDFFE_PN0P_  (.CLK(clknet_leaf_97_clk_p2c),
    .RESET_B(net1382),
    .D(_00886_),
    .Q_N(_05915_),
    .Q(\shift_storage.storage [265]));
 sg13g2_dfrbp_1 \shift_storage.storage[266]$_SDFFE_PN0P_  (.CLK(clknet_leaf_97_clk_p2c),
    .RESET_B(net1383),
    .D(_00887_),
    .Q_N(_05914_),
    .Q(\shift_storage.storage [266]));
 sg13g2_dfrbp_1 \shift_storage.storage[267]$_SDFFE_PN0P_  (.CLK(clknet_leaf_99_clk_p2c),
    .RESET_B(net1384),
    .D(_00888_),
    .Q_N(_05913_),
    .Q(\shift_storage.storage [267]));
 sg13g2_dfrbp_1 \shift_storage.storage[268]$_SDFFE_PN0P_  (.CLK(clknet_leaf_98_clk_p2c),
    .RESET_B(net1385),
    .D(_00889_),
    .Q_N(_05912_),
    .Q(\shift_storage.storage [268]));
 sg13g2_dfrbp_1 \shift_storage.storage[269]$_SDFFE_PN0P_  (.CLK(clknet_leaf_98_clk_p2c),
    .RESET_B(net1386),
    .D(_00890_),
    .Q_N(_05911_),
    .Q(\shift_storage.storage [269]));
 sg13g2_dfrbp_1 \shift_storage.storage[26]$_SDFFE_PN0P_  (.CLK(clknet_leaf_99_clk_p2c),
    .RESET_B(net1387),
    .D(_00891_),
    .Q_N(_05910_),
    .Q(\shift_storage.storage [26]));
 sg13g2_dfrbp_1 \shift_storage.storage[270]$_SDFFE_PN0P_  (.CLK(clknet_leaf_98_clk_p2c),
    .RESET_B(net1388),
    .D(_00892_),
    .Q_N(_05909_),
    .Q(\shift_storage.storage [270]));
 sg13g2_dfrbp_1 \shift_storage.storage[271]$_SDFFE_PN0P_  (.CLK(clknet_leaf_98_clk_p2c),
    .RESET_B(net1389),
    .D(_00893_),
    .Q_N(_05908_),
    .Q(\shift_storage.storage [271]));
 sg13g2_dfrbp_1 \shift_storage.storage[272]$_SDFFE_PN0P_  (.CLK(clknet_leaf_95_clk_p2c),
    .RESET_B(net1390),
    .D(_00894_),
    .Q_N(_05907_),
    .Q(\shift_storage.storage [272]));
 sg13g2_dfrbp_1 \shift_storage.storage[273]$_SDFFE_PN0P_  (.CLK(clknet_leaf_95_clk_p2c),
    .RESET_B(net1391),
    .D(_00895_),
    .Q_N(_05906_),
    .Q(\shift_storage.storage [273]));
 sg13g2_dfrbp_1 \shift_storage.storage[274]$_SDFFE_PN0P_  (.CLK(clknet_leaf_97_clk_p2c),
    .RESET_B(net1392),
    .D(_00896_),
    .Q_N(_05905_),
    .Q(\shift_storage.storage [274]));
 sg13g2_dfrbp_1 \shift_storage.storage[275]$_SDFFE_PN0P_  (.CLK(clknet_leaf_97_clk_p2c),
    .RESET_B(net1393),
    .D(_00897_),
    .Q_N(_05904_),
    .Q(\shift_storage.storage [275]));
 sg13g2_dfrbp_1 \shift_storage.storage[276]$_SDFFE_PN0P_  (.CLK(clknet_leaf_97_clk_p2c),
    .RESET_B(net1394),
    .D(_00898_),
    .Q_N(_05903_),
    .Q(\shift_storage.storage [276]));
 sg13g2_dfrbp_1 \shift_storage.storage[277]$_SDFFE_PN0P_  (.CLK(clknet_leaf_97_clk_p2c),
    .RESET_B(net1395),
    .D(_00899_),
    .Q_N(_05902_),
    .Q(\shift_storage.storage [277]));
 sg13g2_dfrbp_1 \shift_storage.storage[278]$_SDFFE_PN0P_  (.CLK(clknet_leaf_96_clk_p2c),
    .RESET_B(net1396),
    .D(_00900_),
    .Q_N(_05901_),
    .Q(\shift_storage.storage [278]));
 sg13g2_dfrbp_1 \shift_storage.storage[279]$_SDFFE_PN0P_  (.CLK(clknet_leaf_95_clk_p2c),
    .RESET_B(net1397),
    .D(_00901_),
    .Q_N(_05900_),
    .Q(\shift_storage.storage [279]));
 sg13g2_dfrbp_1 \shift_storage.storage[27]$_SDFFE_PN0P_  (.CLK(clknet_leaf_95_clk_p2c),
    .RESET_B(net1398),
    .D(_00902_),
    .Q_N(_05899_),
    .Q(\shift_storage.storage [27]));
 sg13g2_dfrbp_1 \shift_storage.storage[280]$_SDFFE_PN0P_  (.CLK(clknet_leaf_96_clk_p2c),
    .RESET_B(net1399),
    .D(_00903_),
    .Q_N(_05898_),
    .Q(\shift_storage.storage [280]));
 sg13g2_dfrbp_1 \shift_storage.storage[281]$_SDFFE_PN0P_  (.CLK(clknet_leaf_96_clk_p2c),
    .RESET_B(net1400),
    .D(_00904_),
    .Q_N(_05897_),
    .Q(\shift_storage.storage [281]));
 sg13g2_dfrbp_1 \shift_storage.storage[282]$_SDFFE_PN0P_  (.CLK(clknet_leaf_96_clk_p2c),
    .RESET_B(net1401),
    .D(_00905_),
    .Q_N(_05896_),
    .Q(\shift_storage.storage [282]));
 sg13g2_dfrbp_1 \shift_storage.storage[283]$_SDFFE_PN0P_  (.CLK(clknet_leaf_88_clk_p2c),
    .RESET_B(net1402),
    .D(_00906_),
    .Q_N(_05895_),
    .Q(\shift_storage.storage [283]));
 sg13g2_dfrbp_1 \shift_storage.storage[284]$_SDFFE_PN0P_  (.CLK(clknet_leaf_88_clk_p2c),
    .RESET_B(net1403),
    .D(_00907_),
    .Q_N(_05894_),
    .Q(\shift_storage.storage [284]));
 sg13g2_dfrbp_1 \shift_storage.storage[285]$_SDFFE_PN0P_  (.CLK(clknet_leaf_88_clk_p2c),
    .RESET_B(net1404),
    .D(_00908_),
    .Q_N(_05893_),
    .Q(\shift_storage.storage [285]));
 sg13g2_dfrbp_1 \shift_storage.storage[286]$_SDFFE_PN0P_  (.CLK(clknet_leaf_88_clk_p2c),
    .RESET_B(net1405),
    .D(_00909_),
    .Q_N(_05892_),
    .Q(\shift_storage.storage [286]));
 sg13g2_dfrbp_1 \shift_storage.storage[287]$_SDFFE_PN0P_  (.CLK(clknet_leaf_96_clk_p2c),
    .RESET_B(net1406),
    .D(_00910_),
    .Q_N(_05891_),
    .Q(\shift_storage.storage [287]));
 sg13g2_dfrbp_1 \shift_storage.storage[288]$_SDFFE_PN0P_  (.CLK(clknet_leaf_96_clk_p2c),
    .RESET_B(net1407),
    .D(_00911_),
    .Q_N(_05890_),
    .Q(\shift_storage.storage [288]));
 sg13g2_dfrbp_1 \shift_storage.storage[289]$_SDFFE_PN0P_  (.CLK(clknet_leaf_95_clk_p2c),
    .RESET_B(net1408),
    .D(_00912_),
    .Q_N(_05889_),
    .Q(\shift_storage.storage [289]));
 sg13g2_dfrbp_1 \shift_storage.storage[28]$_SDFFE_PN0P_  (.CLK(clknet_leaf_93_clk_p2c),
    .RESET_B(net1409),
    .D(_00913_),
    .Q_N(_05888_),
    .Q(\shift_storage.storage [28]));
 sg13g2_dfrbp_1 \shift_storage.storage[290]$_SDFFE_PN0P_  (.CLK(clknet_leaf_93_clk_p2c),
    .RESET_B(net1410),
    .D(_00914_),
    .Q_N(_05887_),
    .Q(\shift_storage.storage [290]));
 sg13g2_dfrbp_1 \shift_storage.storage[291]$_SDFFE_PN0P_  (.CLK(clknet_leaf_93_clk_p2c),
    .RESET_B(net1411),
    .D(_00915_),
    .Q_N(_05886_),
    .Q(\shift_storage.storage [291]));
 sg13g2_dfrbp_1 \shift_storage.storage[292]$_SDFFE_PN0P_  (.CLK(clknet_leaf_93_clk_p2c),
    .RESET_B(net1412),
    .D(_00916_),
    .Q_N(_05885_),
    .Q(\shift_storage.storage [292]));
 sg13g2_dfrbp_1 \shift_storage.storage[293]$_SDFFE_PN0P_  (.CLK(clknet_leaf_90_clk_p2c),
    .RESET_B(net1413),
    .D(_00917_),
    .Q_N(_05884_),
    .Q(\shift_storage.storage [293]));
 sg13g2_dfrbp_1 \shift_storage.storage[294]$_SDFFE_PN0P_  (.CLK(clknet_leaf_90_clk_p2c),
    .RESET_B(net1414),
    .D(_00918_),
    .Q_N(_05883_),
    .Q(\shift_storage.storage [294]));
 sg13g2_dfrbp_1 \shift_storage.storage[295]$_SDFFE_PN0P_  (.CLK(clknet_leaf_89_clk_p2c),
    .RESET_B(net1415),
    .D(_00919_),
    .Q_N(_05882_),
    .Q(\shift_storage.storage [295]));
 sg13g2_dfrbp_1 \shift_storage.storage[296]$_SDFFE_PN0P_  (.CLK(clknet_leaf_90_clk_p2c),
    .RESET_B(net1416),
    .D(_00920_),
    .Q_N(_05881_),
    .Q(\shift_storage.storage [296]));
 sg13g2_dfrbp_1 \shift_storage.storage[297]$_SDFFE_PN0P_  (.CLK(clknet_leaf_90_clk_p2c),
    .RESET_B(net1417),
    .D(_00921_),
    .Q_N(_05880_),
    .Q(\shift_storage.storage [297]));
 sg13g2_dfrbp_1 \shift_storage.storage[298]$_SDFFE_PN0P_  (.CLK(clknet_leaf_90_clk_p2c),
    .RESET_B(net1418),
    .D(_00922_),
    .Q_N(_05879_),
    .Q(\shift_storage.storage [298]));
 sg13g2_dfrbp_1 \shift_storage.storage[299]$_SDFFE_PN0P_  (.CLK(clknet_leaf_90_clk_p2c),
    .RESET_B(net1419),
    .D(_00923_),
    .Q_N(_05878_),
    .Q(\shift_storage.storage [299]));
 sg13g2_dfrbp_1 \shift_storage.storage[29]$_SDFFE_PN0P_  (.CLK(clknet_leaf_93_clk_p2c),
    .RESET_B(net1420),
    .D(_00924_),
    .Q_N(_05877_),
    .Q(\shift_storage.storage [29]));
 sg13g2_dfrbp_1 \shift_storage.storage[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_91_clk_p2c),
    .RESET_B(net1421),
    .D(_00925_),
    .Q_N(_05876_),
    .Q(\shift_storage.storage [2]));
 sg13g2_dfrbp_1 \shift_storage.storage[300]$_SDFFE_PN0P_  (.CLK(clknet_leaf_91_clk_p2c),
    .RESET_B(net1422),
    .D(_00926_),
    .Q_N(_05875_),
    .Q(\shift_storage.storage [300]));
 sg13g2_dfrbp_1 \shift_storage.storage[301]$_SDFFE_PN0P_  (.CLK(clknet_leaf_91_clk_p2c),
    .RESET_B(net1423),
    .D(_00927_),
    .Q_N(_05874_),
    .Q(\shift_storage.storage [301]));
 sg13g2_dfrbp_1 \shift_storage.storage[302]$_SDFFE_PN0P_  (.CLK(clknet_leaf_91_clk_p2c),
    .RESET_B(net1424),
    .D(_00928_),
    .Q_N(_05873_),
    .Q(\shift_storage.storage [302]));
 sg13g2_dfrbp_1 \shift_storage.storage[303]$_SDFFE_PN0P_  (.CLK(clknet_leaf_91_clk_p2c),
    .RESET_B(net1425),
    .D(_00929_),
    .Q_N(_05872_),
    .Q(\shift_storage.storage [303]));
 sg13g2_dfrbp_1 \shift_storage.storage[304]$_SDFFE_PN0P_  (.CLK(clknet_leaf_92_clk_p2c),
    .RESET_B(net1426),
    .D(_00930_),
    .Q_N(_05871_),
    .Q(\shift_storage.storage [304]));
 sg13g2_dfrbp_1 \shift_storage.storage[305]$_SDFFE_PN0P_  (.CLK(clknet_leaf_92_clk_p2c),
    .RESET_B(net1427),
    .D(_00931_),
    .Q_N(_05870_),
    .Q(\shift_storage.storage [305]));
 sg13g2_dfrbp_1 \shift_storage.storage[306]$_SDFFE_PN0P_  (.CLK(clknet_leaf_92_clk_p2c),
    .RESET_B(net1428),
    .D(_00932_),
    .Q_N(_05869_),
    .Q(\shift_storage.storage [306]));
 sg13g2_dfrbp_1 \shift_storage.storage[307]$_SDFFE_PN0P_  (.CLK(clknet_leaf_91_clk_p2c),
    .RESET_B(net1429),
    .D(_00933_),
    .Q_N(_05868_),
    .Q(\shift_storage.storage [307]));
 sg13g2_dfrbp_1 \shift_storage.storage[308]$_SDFFE_PN0P_  (.CLK(clknet_leaf_92_clk_p2c),
    .RESET_B(net1430),
    .D(_00934_),
    .Q_N(_05867_),
    .Q(\shift_storage.storage [308]));
 sg13g2_dfrbp_1 \shift_storage.storage[309]$_SDFFE_PN0P_  (.CLK(clknet_leaf_92_clk_p2c),
    .RESET_B(net1431),
    .D(_00935_),
    .Q_N(_05866_),
    .Q(\shift_storage.storage [309]));
 sg13g2_dfrbp_1 \shift_storage.storage[30]$_SDFFE_PN0P_  (.CLK(clknet_leaf_93_clk_p2c),
    .RESET_B(net1432),
    .D(_00936_),
    .Q_N(_05865_),
    .Q(\shift_storage.storage [30]));
 sg13g2_dfrbp_1 \shift_storage.storage[310]$_SDFFE_PN0P_  (.CLK(clknet_leaf_112_clk_p2c),
    .RESET_B(net1433),
    .D(_00937_),
    .Q_N(_05864_),
    .Q(\shift_storage.storage [310]));
 sg13g2_dfrbp_1 \shift_storage.storage[311]$_SDFFE_PN0P_  (.CLK(clknet_leaf_112_clk_p2c),
    .RESET_B(net1434),
    .D(_00938_),
    .Q_N(_05863_),
    .Q(\shift_storage.storage [311]));
 sg13g2_dfrbp_1 \shift_storage.storage[312]$_SDFFE_PN0P_  (.CLK(clknet_leaf_110_clk_p2c),
    .RESET_B(net1435),
    .D(_00939_),
    .Q_N(_05862_),
    .Q(\shift_storage.storage [312]));
 sg13g2_dfrbp_1 \shift_storage.storage[313]$_SDFFE_PN0P_  (.CLK(clknet_leaf_110_clk_p2c),
    .RESET_B(net1436),
    .D(_00940_),
    .Q_N(_05861_),
    .Q(\shift_storage.storage [313]));
 sg13g2_dfrbp_1 \shift_storage.storage[314]$_SDFFE_PN0P_  (.CLK(clknet_leaf_110_clk_p2c),
    .RESET_B(net1437),
    .D(_00941_),
    .Q_N(_05860_),
    .Q(\shift_storage.storage [314]));
 sg13g2_dfrbp_1 \shift_storage.storage[315]$_SDFFE_PN0P_  (.CLK(clknet_leaf_94_clk_p2c),
    .RESET_B(net1438),
    .D(_00942_),
    .Q_N(_05859_),
    .Q(\shift_storage.storage [315]));
 sg13g2_dfrbp_1 \shift_storage.storage[316]$_SDFFE_PN0P_  (.CLK(clknet_leaf_94_clk_p2c),
    .RESET_B(net1439),
    .D(_00943_),
    .Q_N(_05858_),
    .Q(\shift_storage.storage [316]));
 sg13g2_dfrbp_1 \shift_storage.storage[317]$_SDFFE_PN0P_  (.CLK(clknet_leaf_94_clk_p2c),
    .RESET_B(net1440),
    .D(_00944_),
    .Q_N(_05857_),
    .Q(\shift_storage.storage [317]));
 sg13g2_dfrbp_1 \shift_storage.storage[318]$_SDFFE_PN0P_  (.CLK(clknet_leaf_94_clk_p2c),
    .RESET_B(net1441),
    .D(_00945_),
    .Q_N(_05856_),
    .Q(\shift_storage.storage [318]));
 sg13g2_dfrbp_1 \shift_storage.storage[319]$_SDFFE_PN0P_  (.CLK(clknet_leaf_94_clk_p2c),
    .RESET_B(net1442),
    .D(_00946_),
    .Q_N(_05855_),
    .Q(\shift_storage.storage [319]));
 sg13g2_dfrbp_1 \shift_storage.storage[31]$_SDFFE_PN0P_  (.CLK(clknet_leaf_110_clk_p2c),
    .RESET_B(net1443),
    .D(_00947_),
    .Q_N(_05854_),
    .Q(\shift_storage.storage [31]));
 sg13g2_dfrbp_1 \shift_storage.storage[320]$_SDFFE_PN0P_  (.CLK(clknet_leaf_94_clk_p2c),
    .RESET_B(net1444),
    .D(_00948_),
    .Q_N(_05853_),
    .Q(\shift_storage.storage [320]));
 sg13g2_dfrbp_1 \shift_storage.storage[321]$_SDFFE_PN0P_  (.CLK(clknet_leaf_110_clk_p2c),
    .RESET_B(net1445),
    .D(_00949_),
    .Q_N(_05852_),
    .Q(\shift_storage.storage [321]));
 sg13g2_dfrbp_1 \shift_storage.storage[322]$_SDFFE_PN0P_  (.CLK(clknet_leaf_98_clk_p2c),
    .RESET_B(net1446),
    .D(_00950_),
    .Q_N(_05851_),
    .Q(\shift_storage.storage [322]));
 sg13g2_dfrbp_1 \shift_storage.storage[323]$_SDFFE_PN0P_  (.CLK(clknet_leaf_98_clk_p2c),
    .RESET_B(net1447),
    .D(_00951_),
    .Q_N(_05850_),
    .Q(\shift_storage.storage [323]));
 sg13g2_dfrbp_1 \shift_storage.storage[324]$_SDFFE_PN0P_  (.CLK(clknet_leaf_104_clk_p2c),
    .RESET_B(net1448),
    .D(_00952_),
    .Q_N(_05849_),
    .Q(\shift_storage.storage [324]));
 sg13g2_dfrbp_1 \shift_storage.storage[325]$_SDFFE_PN0P_  (.CLK(clknet_leaf_104_clk_p2c),
    .RESET_B(net1449),
    .D(_00953_),
    .Q_N(_05848_),
    .Q(\shift_storage.storage [325]));
 sg13g2_dfrbp_1 \shift_storage.storage[326]$_SDFFE_PN0P_  (.CLK(clknet_leaf_104_clk_p2c),
    .RESET_B(net1450),
    .D(_00954_),
    .Q_N(_05847_),
    .Q(\shift_storage.storage [326]));
 sg13g2_dfrbp_1 \shift_storage.storage[327]$_SDFFE_PN0P_  (.CLK(clknet_leaf_104_clk_p2c),
    .RESET_B(net1451),
    .D(_00955_),
    .Q_N(_05846_),
    .Q(\shift_storage.storage [327]));
 sg13g2_dfrbp_1 \shift_storage.storage[328]$_SDFFE_PN0P_  (.CLK(clknet_leaf_109_clk_p2c),
    .RESET_B(net1452),
    .D(_00956_),
    .Q_N(_05845_),
    .Q(\shift_storage.storage [328]));
 sg13g2_dfrbp_1 \shift_storage.storage[329]$_SDFFE_PN0P_  (.CLK(clknet_leaf_109_clk_p2c),
    .RESET_B(net1453),
    .D(_00957_),
    .Q_N(_05844_),
    .Q(\shift_storage.storage [329]));
 sg13g2_dfrbp_1 \shift_storage.storage[32]$_SDFFE_PN0P_  (.CLK(clknet_leaf_110_clk_p2c),
    .RESET_B(net1454),
    .D(_00958_),
    .Q_N(_05843_),
    .Q(\shift_storage.storage [32]));
 sg13g2_dfrbp_1 \shift_storage.storage[330]$_SDFFE_PN0P_  (.CLK(clknet_leaf_109_clk_p2c),
    .RESET_B(net1455),
    .D(_00959_),
    .Q_N(_05842_),
    .Q(\shift_storage.storage [330]));
 sg13g2_dfrbp_1 \shift_storage.storage[331]$_SDFFE_PN0P_  (.CLK(clknet_leaf_109_clk_p2c),
    .RESET_B(net1456),
    .D(_00960_),
    .Q_N(_05841_),
    .Q(\shift_storage.storage [331]));
 sg13g2_dfrbp_1 \shift_storage.storage[332]$_SDFFE_PN0P_  (.CLK(clknet_leaf_109_clk_p2c),
    .RESET_B(net1457),
    .D(_00961_),
    .Q_N(_05840_),
    .Q(\shift_storage.storage [332]));
 sg13g2_dfrbp_1 \shift_storage.storage[333]$_SDFFE_PN0P_  (.CLK(clknet_leaf_110_clk_p2c),
    .RESET_B(net1458),
    .D(_00962_),
    .Q_N(_05839_),
    .Q(\shift_storage.storage [333]));
 sg13g2_dfrbp_1 \shift_storage.storage[334]$_SDFFE_PN0P_  (.CLK(clknet_leaf_111_clk_p2c),
    .RESET_B(net1459),
    .D(_00963_),
    .Q_N(_05838_),
    .Q(\shift_storage.storage [334]));
 sg13g2_dfrbp_1 \shift_storage.storage[335]$_SDFFE_PN0P_  (.CLK(clknet_leaf_111_clk_p2c),
    .RESET_B(net1460),
    .D(_00964_),
    .Q_N(_05837_),
    .Q(\shift_storage.storage [335]));
 sg13g2_dfrbp_1 \shift_storage.storage[336]$_SDFFE_PN0P_  (.CLK(clknet_leaf_108_clk_p2c),
    .RESET_B(net1461),
    .D(_00965_),
    .Q_N(_05836_),
    .Q(\shift_storage.storage [336]));
 sg13g2_dfrbp_1 \shift_storage.storage[337]$_SDFFE_PN0P_  (.CLK(clknet_leaf_108_clk_p2c),
    .RESET_B(net1462),
    .D(_00966_),
    .Q_N(_05835_),
    .Q(\shift_storage.storage [337]));
 sg13g2_dfrbp_1 \shift_storage.storage[338]$_SDFFE_PN0P_  (.CLK(clknet_leaf_108_clk_p2c),
    .RESET_B(net1463),
    .D(_00967_),
    .Q_N(_05834_),
    .Q(\shift_storage.storage [338]));
 sg13g2_dfrbp_1 \shift_storage.storage[339]$_SDFFE_PN0P_  (.CLK(clknet_leaf_108_clk_p2c),
    .RESET_B(net1464),
    .D(_00968_),
    .Q_N(_05833_),
    .Q(\shift_storage.storage [339]));
 sg13g2_dfrbp_1 \shift_storage.storage[33]$_SDFFE_PN0P_  (.CLK(clknet_leaf_111_clk_p2c),
    .RESET_B(net1465),
    .D(_00969_),
    .Q_N(_05832_),
    .Q(\shift_storage.storage [33]));
 sg13g2_dfrbp_1 \shift_storage.storage[340]$_SDFFE_PN0P_  (.CLK(clknet_leaf_107_clk_p2c),
    .RESET_B(net1466),
    .D(_00970_),
    .Q_N(_05831_),
    .Q(\shift_storage.storage [340]));
 sg13g2_dfrbp_1 \shift_storage.storage[341]$_SDFFE_PN0P_  (.CLK(clknet_leaf_108_clk_p2c),
    .RESET_B(net1467),
    .D(_00971_),
    .Q_N(_05830_),
    .Q(\shift_storage.storage [341]));
 sg13g2_dfrbp_1 \shift_storage.storage[342]$_SDFFE_PN0P_  (.CLK(clknet_leaf_108_clk_p2c),
    .RESET_B(net1468),
    .D(_00972_),
    .Q_N(_05829_),
    .Q(\shift_storage.storage [342]));
 sg13g2_dfrbp_1 \shift_storage.storage[343]$_SDFFE_PN0P_  (.CLK(clknet_leaf_117_clk_p2c),
    .RESET_B(net1469),
    .D(_00973_),
    .Q_N(_05828_),
    .Q(\shift_storage.storage [343]));
 sg13g2_dfrbp_1 \shift_storage.storage[344]$_SDFFE_PN0P_  (.CLK(clknet_leaf_118_clk_p2c),
    .RESET_B(net1470),
    .D(_00974_),
    .Q_N(_05827_),
    .Q(\shift_storage.storage [344]));
 sg13g2_dfrbp_1 \shift_storage.storage[345]$_SDFFE_PN0P_  (.CLK(clknet_leaf_118_clk_p2c),
    .RESET_B(net1471),
    .D(_00975_),
    .Q_N(_05826_),
    .Q(\shift_storage.storage [345]));
 sg13g2_dfrbp_1 \shift_storage.storage[346]$_SDFFE_PN0P_  (.CLK(clknet_leaf_118_clk_p2c),
    .RESET_B(net1472),
    .D(_00976_),
    .Q_N(_05825_),
    .Q(\shift_storage.storage [346]));
 sg13g2_dfrbp_1 \shift_storage.storage[347]$_SDFFE_PN0P_  (.CLK(clknet_leaf_117_clk_p2c),
    .RESET_B(net1473),
    .D(_00977_),
    .Q_N(_05824_),
    .Q(\shift_storage.storage [347]));
 sg13g2_dfrbp_1 \shift_storage.storage[348]$_SDFFE_PN0P_  (.CLK(clknet_leaf_117_clk_p2c),
    .RESET_B(net1474),
    .D(_00978_),
    .Q_N(_05823_),
    .Q(\shift_storage.storage [348]));
 sg13g2_dfrbp_1 \shift_storage.storage[349]$_SDFFE_PN0P_  (.CLK(clknet_leaf_117_clk_p2c),
    .RESET_B(net1475),
    .D(_00979_),
    .Q_N(_05822_),
    .Q(\shift_storage.storage [349]));
 sg13g2_dfrbp_1 \shift_storage.storage[34]$_SDFFE_PN0P_  (.CLK(clknet_leaf_117_clk_p2c),
    .RESET_B(net1476),
    .D(_00980_),
    .Q_N(_05821_),
    .Q(\shift_storage.storage [34]));
 sg13g2_dfrbp_1 \shift_storage.storage[350]$_SDFFE_PN0P_  (.CLK(clknet_leaf_114_clk_p2c),
    .RESET_B(net1477),
    .D(_00981_),
    .Q_N(_05820_),
    .Q(\shift_storage.storage [350]));
 sg13g2_dfrbp_1 \shift_storage.storage[351]$_SDFFE_PN0P_  (.CLK(clknet_leaf_114_clk_p2c),
    .RESET_B(net1478),
    .D(_00982_),
    .Q_N(_05819_),
    .Q(\shift_storage.storage [351]));
 sg13g2_dfrbp_1 \shift_storage.storage[352]$_SDFFE_PN0P_  (.CLK(clknet_leaf_114_clk_p2c),
    .RESET_B(net1479),
    .D(_00983_),
    .Q_N(_05818_),
    .Q(\shift_storage.storage [352]));
 sg13g2_dfrbp_1 \shift_storage.storage[353]$_SDFFE_PN0P_  (.CLK(clknet_leaf_114_clk_p2c),
    .RESET_B(net1480),
    .D(_00984_),
    .Q_N(_05817_),
    .Q(\shift_storage.storage [353]));
 sg13g2_dfrbp_1 \shift_storage.storage[354]$_SDFFE_PN0P_  (.CLK(clknet_leaf_114_clk_p2c),
    .RESET_B(net1481),
    .D(_00985_),
    .Q_N(_05816_),
    .Q(\shift_storage.storage [354]));
 sg13g2_dfrbp_1 \shift_storage.storage[355]$_SDFFE_PN0P_  (.CLK(clknet_leaf_111_clk_p2c),
    .RESET_B(net1482),
    .D(_00986_),
    .Q_N(_05815_),
    .Q(\shift_storage.storage [355]));
 sg13g2_dfrbp_1 \shift_storage.storage[356]$_SDFFE_PN0P_  (.CLK(clknet_leaf_111_clk_p2c),
    .RESET_B(net1483),
    .D(_00987_),
    .Q_N(_05814_),
    .Q(\shift_storage.storage [356]));
 sg13g2_dfrbp_1 \shift_storage.storage[357]$_SDFFE_PN0P_  (.CLK(clknet_leaf_111_clk_p2c),
    .RESET_B(net1484),
    .D(_00988_),
    .Q_N(_05813_),
    .Q(\shift_storage.storage [357]));
 sg13g2_dfrbp_1 \shift_storage.storage[358]$_SDFFE_PN0P_  (.CLK(clknet_leaf_112_clk_p2c),
    .RESET_B(net1485),
    .D(_00989_),
    .Q_N(_05812_),
    .Q(\shift_storage.storage [358]));
 sg13g2_dfrbp_1 \shift_storage.storage[359]$_SDFFE_PN0P_  (.CLK(clknet_leaf_112_clk_p2c),
    .RESET_B(net1486),
    .D(_00990_),
    .Q_N(_05811_),
    .Q(\shift_storage.storage [359]));
 sg13g2_dfrbp_1 \shift_storage.storage[35]$_SDFFE_PN0P_  (.CLK(clknet_leaf_113_clk_p2c),
    .RESET_B(net1487),
    .D(_00991_),
    .Q_N(_05810_),
    .Q(\shift_storage.storage [35]));
 sg13g2_dfrbp_1 \shift_storage.storage[360]$_SDFFE_PN0P_  (.CLK(clknet_leaf_112_clk_p2c),
    .RESET_B(net1488),
    .D(_00992_),
    .Q_N(_05809_),
    .Q(\shift_storage.storage [360]));
 sg13g2_dfrbp_1 \shift_storage.storage[361]$_SDFFE_PN0P_  (.CLK(clknet_leaf_112_clk_p2c),
    .RESET_B(net1489),
    .D(_00993_),
    .Q_N(_05808_),
    .Q(\shift_storage.storage [361]));
 sg13g2_dfrbp_1 \shift_storage.storage[362]$_SDFFE_PN0P_  (.CLK(clknet_leaf_113_clk_p2c),
    .RESET_B(net1490),
    .D(_00994_),
    .Q_N(_05807_),
    .Q(\shift_storage.storage [362]));
 sg13g2_dfrbp_1 \shift_storage.storage[363]$_SDFFE_PN0P_  (.CLK(clknet_leaf_113_clk_p2c),
    .RESET_B(net1491),
    .D(_00995_),
    .Q_N(_05806_),
    .Q(\shift_storage.storage [363]));
 sg13g2_dfrbp_1 \shift_storage.storage[364]$_SDFFE_PN0P_  (.CLK(clknet_leaf_113_clk_p2c),
    .RESET_B(net1492),
    .D(_00996_),
    .Q_N(_05805_),
    .Q(\shift_storage.storage [364]));
 sg13g2_dfrbp_1 \shift_storage.storage[365]$_SDFFE_PN0P_  (.CLK(clknet_leaf_113_clk_p2c),
    .RESET_B(net1493),
    .D(_00997_),
    .Q_N(_05804_),
    .Q(\shift_storage.storage [365]));
 sg13g2_dfrbp_1 \shift_storage.storage[366]$_SDFFE_PN0P_  (.CLK(clknet_leaf_114_clk_p2c),
    .RESET_B(net1494),
    .D(_00998_),
    .Q_N(_05803_),
    .Q(\shift_storage.storage [366]));
 sg13g2_dfrbp_1 \shift_storage.storage[367]$_SDFFE_PN0P_  (.CLK(clknet_leaf_58_clk_p2c),
    .RESET_B(net1495),
    .D(_00999_),
    .Q_N(_05802_),
    .Q(\shift_storage.storage [367]));
 sg13g2_dfrbp_1 \shift_storage.storage[368]$_SDFFE_PN0P_  (.CLK(clknet_leaf_58_clk_p2c),
    .RESET_B(net1496),
    .D(_01000_),
    .Q_N(_05801_),
    .Q(\shift_storage.storage [368]));
 sg13g2_dfrbp_1 \shift_storage.storage[369]$_SDFFE_PN0P_  (.CLK(clknet_leaf_58_clk_p2c),
    .RESET_B(net1497),
    .D(_01001_),
    .Q_N(_05800_),
    .Q(\shift_storage.storage [369]));
 sg13g2_dfrbp_1 \shift_storage.storage[36]$_SDFFE_PN0P_  (.CLK(clknet_leaf_58_clk_p2c),
    .RESET_B(net1498),
    .D(_01002_),
    .Q_N(_05799_),
    .Q(\shift_storage.storage [36]));
 sg13g2_dfrbp_1 \shift_storage.storage[370]$_SDFFE_PN0P_  (.CLK(clknet_leaf_57_clk_p2c),
    .RESET_B(net1499),
    .D(_01003_),
    .Q_N(_05798_),
    .Q(\shift_storage.storage [370]));
 sg13g2_dfrbp_1 \shift_storage.storage[371]$_SDFFE_PN0P_  (.CLK(clknet_leaf_56_clk_p2c),
    .RESET_B(net1500),
    .D(_01004_),
    .Q_N(_05797_),
    .Q(\shift_storage.storage [371]));
 sg13g2_dfrbp_1 \shift_storage.storage[372]$_SDFFE_PN0P_  (.CLK(clknet_leaf_115_clk_p2c),
    .RESET_B(net1501),
    .D(_01005_),
    .Q_N(_05796_),
    .Q(\shift_storage.storage [372]));
 sg13g2_dfrbp_1 \shift_storage.storage[373]$_SDFFE_PN0P_  (.CLK(clknet_leaf_115_clk_p2c),
    .RESET_B(net1502),
    .D(_01006_),
    .Q_N(_05795_),
    .Q(\shift_storage.storage [373]));
 sg13g2_dfrbp_1 \shift_storage.storage[374]$_SDFFE_PN0P_  (.CLK(clknet_leaf_115_clk_p2c),
    .RESET_B(net1503),
    .D(_01007_),
    .Q_N(_05794_),
    .Q(\shift_storage.storage [374]));
 sg13g2_dfrbp_1 \shift_storage.storage[375]$_SDFFE_PN0P_  (.CLK(clknet_leaf_116_clk_p2c),
    .RESET_B(net1504),
    .D(_01008_),
    .Q_N(_05793_),
    .Q(\shift_storage.storage [375]));
 sg13g2_dfrbp_1 \shift_storage.storage[376]$_SDFFE_PN0P_  (.CLK(clknet_leaf_115_clk_p2c),
    .RESET_B(net1505),
    .D(_01009_),
    .Q_N(_05792_),
    .Q(\shift_storage.storage [376]));
 sg13g2_dfrbp_1 \shift_storage.storage[377]$_SDFFE_PN0P_  (.CLK(clknet_leaf_115_clk_p2c),
    .RESET_B(net1506),
    .D(_01010_),
    .Q_N(_05791_),
    .Q(\shift_storage.storage [377]));
 sg13g2_dfrbp_1 \shift_storage.storage[378]$_SDFFE_PN0P_  (.CLK(clknet_leaf_56_clk_p2c),
    .RESET_B(net1507),
    .D(_01011_),
    .Q_N(_05790_),
    .Q(\shift_storage.storage [378]));
 sg13g2_dfrbp_1 \shift_storage.storage[379]$_SDFFE_PN0P_  (.CLK(clknet_leaf_56_clk_p2c),
    .RESET_B(net1508),
    .D(_01012_),
    .Q_N(_05789_),
    .Q(\shift_storage.storage [379]));
 sg13g2_dfrbp_1 \shift_storage.storage[37]$_SDFFE_PN0P_  (.CLK(clknet_leaf_57_clk_p2c),
    .RESET_B(net1509),
    .D(_01013_),
    .Q_N(_05788_),
    .Q(\shift_storage.storage [37]));
 sg13g2_dfrbp_1 \shift_storage.storage[380]$_SDFFE_PN0P_  (.CLK(clknet_leaf_57_clk_p2c),
    .RESET_B(net1510),
    .D(_01014_),
    .Q_N(_05787_),
    .Q(\shift_storage.storage [380]));
 sg13g2_dfrbp_1 \shift_storage.storage[381]$_SDFFE_PN0P_  (.CLK(clknet_leaf_57_clk_p2c),
    .RESET_B(net1511),
    .D(_01015_),
    .Q_N(_05786_),
    .Q(\shift_storage.storage [381]));
 sg13g2_dfrbp_1 \shift_storage.storage[382]$_SDFFE_PN0P_  (.CLK(clknet_leaf_57_clk_p2c),
    .RESET_B(net1512),
    .D(_01016_),
    .Q_N(_05785_),
    .Q(\shift_storage.storage [382]));
 sg13g2_dfrbp_1 \shift_storage.storage[383]$_SDFFE_PN0P_  (.CLK(clknet_leaf_55_clk_p2c),
    .RESET_B(net1513),
    .D(_01017_),
    .Q_N(_05784_),
    .Q(\shift_storage.storage [383]));
 sg13g2_dfrbp_1 \shift_storage.storage[384]$_SDFFE_PN0P_  (.CLK(clknet_leaf_55_clk_p2c),
    .RESET_B(net1514),
    .D(_01018_),
    .Q_N(_05783_),
    .Q(\shift_storage.storage [384]));
 sg13g2_dfrbp_1 \shift_storage.storage[385]$_SDFFE_PN0P_  (.CLK(clknet_leaf_54_clk_p2c),
    .RESET_B(net1515),
    .D(_01019_),
    .Q_N(_05782_),
    .Q(\shift_storage.storage [385]));
 sg13g2_dfrbp_1 \shift_storage.storage[386]$_SDFFE_PN0P_  (.CLK(clknet_leaf_54_clk_p2c),
    .RESET_B(net1516),
    .D(_01020_),
    .Q_N(_05781_),
    .Q(\shift_storage.storage [386]));
 sg13g2_dfrbp_1 \shift_storage.storage[387]$_SDFFE_PN0P_  (.CLK(clknet_leaf_54_clk_p2c),
    .RESET_B(net1517),
    .D(_01021_),
    .Q_N(_05780_),
    .Q(\shift_storage.storage [387]));
 sg13g2_dfrbp_1 \shift_storage.storage[388]$_SDFFE_PN0P_  (.CLK(clknet_leaf_54_clk_p2c),
    .RESET_B(net1518),
    .D(_01022_),
    .Q_N(_05779_),
    .Q(\shift_storage.storage [388]));
 sg13g2_dfrbp_1 \shift_storage.storage[389]$_SDFFE_PN0P_  (.CLK(clknet_leaf_54_clk_p2c),
    .RESET_B(net1519),
    .D(_01023_),
    .Q_N(_05778_),
    .Q(\shift_storage.storage [389]));
 sg13g2_dfrbp_1 \shift_storage.storage[38]$_SDFFE_PN0P_  (.CLK(clknet_leaf_57_clk_p2c),
    .RESET_B(net1520),
    .D(_01024_),
    .Q_N(_05777_),
    .Q(\shift_storage.storage [38]));
 sg13g2_dfrbp_1 \shift_storage.storage[390]$_SDFFE_PN0P_  (.CLK(clknet_leaf_54_clk_p2c),
    .RESET_B(net1521),
    .D(_01025_),
    .Q_N(_05776_),
    .Q(\shift_storage.storage [390]));
 sg13g2_dfrbp_1 \shift_storage.storage[391]$_SDFFE_PN0P_  (.CLK(clknet_leaf_54_clk_p2c),
    .RESET_B(net1522),
    .D(_01026_),
    .Q_N(_05775_),
    .Q(\shift_storage.storage [391]));
 sg13g2_dfrbp_1 \shift_storage.storage[392]$_SDFFE_PN0P_  (.CLK(clknet_leaf_52_clk_p2c),
    .RESET_B(net1523),
    .D(_01027_),
    .Q_N(_05774_),
    .Q(\shift_storage.storage [392]));
 sg13g2_dfrbp_1 \shift_storage.storage[393]$_SDFFE_PN0P_  (.CLK(clknet_leaf_53_clk_p2c),
    .RESET_B(net1524),
    .D(_01028_),
    .Q_N(_05773_),
    .Q(\shift_storage.storage [393]));
 sg13g2_dfrbp_1 \shift_storage.storage[394]$_SDFFE_PN0P_  (.CLK(clknet_leaf_64_clk_p2c),
    .RESET_B(net1525),
    .D(_01029_),
    .Q_N(_05772_),
    .Q(\shift_storage.storage [394]));
 sg13g2_dfrbp_1 \shift_storage.storage[395]$_SDFFE_PN0P_  (.CLK(clknet_leaf_64_clk_p2c),
    .RESET_B(net1526),
    .D(_01030_),
    .Q_N(_05771_),
    .Q(\shift_storage.storage [395]));
 sg13g2_dfrbp_1 \shift_storage.storage[396]$_SDFFE_PN0P_  (.CLK(clknet_leaf_64_clk_p2c),
    .RESET_B(net1527),
    .D(_01031_),
    .Q_N(_05770_),
    .Q(\shift_storage.storage [396]));
 sg13g2_dfrbp_1 \shift_storage.storage[397]$_SDFFE_PN0P_  (.CLK(clknet_leaf_64_clk_p2c),
    .RESET_B(net1528),
    .D(_01032_),
    .Q_N(_05769_),
    .Q(\shift_storage.storage [397]));
 sg13g2_dfrbp_1 \shift_storage.storage[398]$_SDFFE_PN0P_  (.CLK(clknet_leaf_63_clk_p2c),
    .RESET_B(net1529),
    .D(_01033_),
    .Q_N(_05768_),
    .Q(\shift_storage.storage [398]));
 sg13g2_dfrbp_1 \shift_storage.storage[399]$_SDFFE_PN0P_  (.CLK(clknet_leaf_63_clk_p2c),
    .RESET_B(net1530),
    .D(_01034_),
    .Q_N(_05767_),
    .Q(\shift_storage.storage [399]));
 sg13g2_dfrbp_1 \shift_storage.storage[39]$_SDFFE_PN0P_  (.CLK(clknet_leaf_60_clk_p2c),
    .RESET_B(net1531),
    .D(_01035_),
    .Q_N(_05766_),
    .Q(\shift_storage.storage [39]));
 sg13g2_dfrbp_1 \shift_storage.storage[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_64_clk_p2c),
    .RESET_B(net1532),
    .D(_01036_),
    .Q_N(_05765_),
    .Q(\shift_storage.storage [3]));
 sg13g2_dfrbp_1 \shift_storage.storage[400]$_SDFFE_PN0P_  (.CLK(clknet_leaf_63_clk_p2c),
    .RESET_B(net1533),
    .D(_01037_),
    .Q_N(_05764_),
    .Q(\shift_storage.storage [400]));
 sg13g2_dfrbp_1 \shift_storage.storage[401]$_SDFFE_PN0P_  (.CLK(clknet_leaf_63_clk_p2c),
    .RESET_B(net1534),
    .D(_01038_),
    .Q_N(_05763_),
    .Q(\shift_storage.storage [401]));
 sg13g2_dfrbp_1 \shift_storage.storage[402]$_SDFFE_PN0P_  (.CLK(clknet_leaf_61_clk_p2c),
    .RESET_B(net1535),
    .D(_01039_),
    .Q_N(_05762_),
    .Q(\shift_storage.storage [402]));
 sg13g2_dfrbp_1 \shift_storage.storage[403]$_SDFFE_PN0P_  (.CLK(clknet_leaf_63_clk_p2c),
    .RESET_B(net1536),
    .D(_01040_),
    .Q_N(_05761_),
    .Q(\shift_storage.storage [403]));
 sg13g2_dfrbp_1 \shift_storage.storage[404]$_SDFFE_PN0P_  (.CLK(clknet_leaf_63_clk_p2c),
    .RESET_B(net1537),
    .D(_01041_),
    .Q_N(_05760_),
    .Q(\shift_storage.storage [404]));
 sg13g2_dfrbp_1 \shift_storage.storage[405]$_SDFFE_PN0P_  (.CLK(clknet_leaf_62_clk_p2c),
    .RESET_B(net1538),
    .D(_01042_),
    .Q_N(_05759_),
    .Q(\shift_storage.storage [405]));
 sg13g2_dfrbp_1 \shift_storage.storage[406]$_SDFFE_PN0P_  (.CLK(clknet_leaf_62_clk_p2c),
    .RESET_B(net1539),
    .D(_01043_),
    .Q_N(_05758_),
    .Q(\shift_storage.storage [406]));
 sg13g2_dfrbp_1 \shift_storage.storage[407]$_SDFFE_PN0P_  (.CLK(clknet_leaf_62_clk_p2c),
    .RESET_B(net1540),
    .D(_01044_),
    .Q_N(_05757_),
    .Q(\shift_storage.storage [407]));
 sg13g2_dfrbp_1 \shift_storage.storage[408]$_SDFFE_PN0P_  (.CLK(clknet_leaf_62_clk_p2c),
    .RESET_B(net1541),
    .D(_01045_),
    .Q_N(_05756_),
    .Q(\shift_storage.storage [408]));
 sg13g2_dfrbp_1 \shift_storage.storage[409]$_SDFFE_PN0P_  (.CLK(clknet_leaf_78_clk_p2c),
    .RESET_B(net1542),
    .D(_01046_),
    .Q_N(_05755_),
    .Q(\shift_storage.storage [409]));
 sg13g2_dfrbp_1 \shift_storage.storage[40]$_SDFFE_PN0P_  (.CLK(clknet_leaf_61_clk_p2c),
    .RESET_B(net1543),
    .D(_01047_),
    .Q_N(_05754_),
    .Q(\shift_storage.storage [40]));
 sg13g2_dfrbp_1 \shift_storage.storage[410]$_SDFFE_PN0P_  (.CLK(clknet_leaf_78_clk_p2c),
    .RESET_B(net1544),
    .D(_01048_),
    .Q_N(_05753_),
    .Q(\shift_storage.storage [410]));
 sg13g2_dfrbp_1 \shift_storage.storage[411]$_SDFFE_PN0P_  (.CLK(clknet_leaf_79_clk_p2c),
    .RESET_B(net1545),
    .D(_01049_),
    .Q_N(_05752_),
    .Q(\shift_storage.storage [411]));
 sg13g2_dfrbp_1 \shift_storage.storage[412]$_SDFFE_PN0P_  (.CLK(clknet_leaf_61_clk_p2c),
    .RESET_B(net1546),
    .D(_01050_),
    .Q_N(_05751_),
    .Q(\shift_storage.storage [412]));
 sg13g2_dfrbp_1 \shift_storage.storage[413]$_SDFFE_PN0P_  (.CLK(clknet_leaf_61_clk_p2c),
    .RESET_B(net1547),
    .D(_01051_),
    .Q_N(_05750_),
    .Q(\shift_storage.storage [413]));
 sg13g2_dfrbp_1 \shift_storage.storage[414]$_SDFFE_PN0P_  (.CLK(clknet_leaf_61_clk_p2c),
    .RESET_B(net1548),
    .D(_01052_),
    .Q_N(_05749_),
    .Q(\shift_storage.storage [414]));
 sg13g2_dfrbp_1 \shift_storage.storage[415]$_SDFFE_PN0P_  (.CLK(clknet_leaf_60_clk_p2c),
    .RESET_B(net1549),
    .D(_01053_),
    .Q_N(_05748_),
    .Q(\shift_storage.storage [415]));
 sg13g2_dfrbp_1 \shift_storage.storage[416]$_SDFFE_PN0P_  (.CLK(clknet_leaf_60_clk_p2c),
    .RESET_B(net1550),
    .D(_01054_),
    .Q_N(_05747_),
    .Q(\shift_storage.storage [416]));
 sg13g2_dfrbp_1 \shift_storage.storage[417]$_SDFFE_PN0P_  (.CLK(clknet_leaf_60_clk_p2c),
    .RESET_B(net1551),
    .D(_01055_),
    .Q_N(_05746_),
    .Q(\shift_storage.storage [417]));
 sg13g2_dfrbp_1 \shift_storage.storage[418]$_SDFFE_PN0P_  (.CLK(clknet_leaf_60_clk_p2c),
    .RESET_B(net1552),
    .D(_01056_),
    .Q_N(_05745_),
    .Q(\shift_storage.storage [418]));
 sg13g2_dfrbp_1 \shift_storage.storage[419]$_SDFFE_PN0P_  (.CLK(clknet_leaf_60_clk_p2c),
    .RESET_B(net1553),
    .D(_01057_),
    .Q_N(_05744_),
    .Q(\shift_storage.storage [419]));
 sg13g2_dfrbp_1 \shift_storage.storage[41]$_SDFFE_PN0P_  (.CLK(clknet_leaf_61_clk_p2c),
    .RESET_B(net1554),
    .D(_01058_),
    .Q_N(_05743_),
    .Q(\shift_storage.storage [41]));
 sg13g2_dfrbp_1 \shift_storage.storage[420]$_SDFFE_PN0P_  (.CLK(clknet_leaf_59_clk_p2c),
    .RESET_B(net1555),
    .D(_01059_),
    .Q_N(_05742_),
    .Q(\shift_storage.storage [420]));
 sg13g2_dfrbp_1 \shift_storage.storage[421]$_SDFFE_PN0P_  (.CLK(clknet_leaf_59_clk_p2c),
    .RESET_B(net1556),
    .D(_01060_),
    .Q_N(_05741_),
    .Q(\shift_storage.storage [421]));
 sg13g2_dfrbp_1 \shift_storage.storage[422]$_SDFFE_PN0P_  (.CLK(clknet_leaf_59_clk_p2c),
    .RESET_B(net1557),
    .D(_01061_),
    .Q_N(_05740_),
    .Q(\shift_storage.storage [422]));
 sg13g2_dfrbp_1 \shift_storage.storage[423]$_SDFFE_PN0P_  (.CLK(clknet_leaf_58_clk_p2c),
    .RESET_B(net1558),
    .D(_01062_),
    .Q_N(_05739_),
    .Q(\shift_storage.storage [423]));
 sg13g2_dfrbp_1 \shift_storage.storage[424]$_SDFFE_PN0P_  (.CLK(clknet_leaf_59_clk_p2c),
    .RESET_B(net1559),
    .D(_01063_),
    .Q_N(_05738_),
    .Q(\shift_storage.storage [424]));
 sg13g2_dfrbp_1 \shift_storage.storage[425]$_SDFFE_PN0P_  (.CLK(clknet_leaf_59_clk_p2c),
    .RESET_B(net1560),
    .D(_01064_),
    .Q_N(_05737_),
    .Q(\shift_storage.storage [425]));
 sg13g2_dfrbp_1 \shift_storage.storage[426]$_SDFFE_PN0P_  (.CLK(clknet_leaf_81_clk_p2c),
    .RESET_B(net1561),
    .D(_01065_),
    .Q_N(_05736_),
    .Q(\shift_storage.storage [426]));
 sg13g2_dfrbp_1 \shift_storage.storage[427]$_SDFFE_PN0P_  (.CLK(clknet_leaf_81_clk_p2c),
    .RESET_B(net1562),
    .D(_01066_),
    .Q_N(_05735_),
    .Q(\shift_storage.storage [427]));
 sg13g2_dfrbp_1 \shift_storage.storage[428]$_SDFFE_PN0P_  (.CLK(clknet_leaf_59_clk_p2c),
    .RESET_B(net1563),
    .D(_01067_),
    .Q_N(_05734_),
    .Q(\shift_storage.storage [428]));
 sg13g2_dfrbp_1 \shift_storage.storage[429]$_SDFFE_PN0P_  (.CLK(clknet_leaf_59_clk_p2c),
    .RESET_B(net1564),
    .D(_01068_),
    .Q_N(_05733_),
    .Q(\shift_storage.storage [429]));
 sg13g2_dfrbp_1 \shift_storage.storage[42]$_SDFFE_PN0P_  (.CLK(clknet_leaf_81_clk_p2c),
    .RESET_B(net1565),
    .D(_01069_),
    .Q_N(_05732_),
    .Q(\shift_storage.storage [42]));
 sg13g2_dfrbp_1 \shift_storage.storage[430]$_SDFFE_PN0P_  (.CLK(clknet_leaf_81_clk_p2c),
    .RESET_B(net1566),
    .D(_01070_),
    .Q_N(_05731_),
    .Q(\shift_storage.storage [430]));
 sg13g2_dfrbp_1 \shift_storage.storage[431]$_SDFFE_PN0P_  (.CLK(clknet_leaf_80_clk_p2c),
    .RESET_B(net1567),
    .D(_01071_),
    .Q_N(_05730_),
    .Q(\shift_storage.storage [431]));
 sg13g2_dfrbp_1 \shift_storage.storage[432]$_SDFFE_PN0P_  (.CLK(clknet_leaf_81_clk_p2c),
    .RESET_B(net1568),
    .D(_01072_),
    .Q_N(_05729_),
    .Q(\shift_storage.storage [432]));
 sg13g2_dfrbp_1 \shift_storage.storage[433]$_SDFFE_PN0P_  (.CLK(clknet_leaf_80_clk_p2c),
    .RESET_B(net1569),
    .D(_01073_),
    .Q_N(_05728_),
    .Q(\shift_storage.storage [433]));
 sg13g2_dfrbp_1 \shift_storage.storage[434]$_SDFFE_PN0P_  (.CLK(clknet_leaf_80_clk_p2c),
    .RESET_B(net1570),
    .D(_01074_),
    .Q_N(_05727_),
    .Q(\shift_storage.storage [434]));
 sg13g2_dfrbp_1 \shift_storage.storage[435]$_SDFFE_PN0P_  (.CLK(clknet_leaf_82_clk_p2c),
    .RESET_B(net1571),
    .D(_01075_),
    .Q_N(_05726_),
    .Q(\shift_storage.storage [435]));
 sg13g2_dfrbp_1 \shift_storage.storage[436]$_SDFFE_PN0P_  (.CLK(clknet_leaf_81_clk_p2c),
    .RESET_B(net1572),
    .D(_01076_),
    .Q_N(_05725_),
    .Q(\shift_storage.storage [436]));
 sg13g2_dfrbp_1 \shift_storage.storage[437]$_SDFFE_PN0P_  (.CLK(clknet_leaf_82_clk_p2c),
    .RESET_B(net1573),
    .D(_01077_),
    .Q_N(_05724_),
    .Q(\shift_storage.storage [437]));
 sg13g2_dfrbp_1 \shift_storage.storage[438]$_SDFFE_PN0P_  (.CLK(clknet_leaf_82_clk_p2c),
    .RESET_B(net1574),
    .D(_01078_),
    .Q_N(_05723_),
    .Q(\shift_storage.storage [438]));
 sg13g2_dfrbp_1 \shift_storage.storage[439]$_SDFFE_PN0P_  (.CLK(clknet_leaf_82_clk_p2c),
    .RESET_B(net1575),
    .D(_01079_),
    .Q_N(_05722_),
    .Q(\shift_storage.storage [439]));
 sg13g2_dfrbp_1 \shift_storage.storage[43]$_SDFFE_PN0P_  (.CLK(clknet_leaf_79_clk_p2c),
    .RESET_B(net1576),
    .D(_01080_),
    .Q_N(_05721_),
    .Q(\shift_storage.storage [43]));
 sg13g2_dfrbp_1 \shift_storage.storage[440]$_SDFFE_PN0P_  (.CLK(clknet_leaf_82_clk_p2c),
    .RESET_B(net1577),
    .D(_01081_),
    .Q_N(_05720_),
    .Q(\shift_storage.storage [440]));
 sg13g2_dfrbp_1 \shift_storage.storage[441]$_SDFFE_PN0P_  (.CLK(clknet_leaf_82_clk_p2c),
    .RESET_B(net1578),
    .D(_01082_),
    .Q_N(_05719_),
    .Q(\shift_storage.storage [441]));
 sg13g2_dfrbp_1 \shift_storage.storage[442]$_SDFFE_PN0P_  (.CLK(clknet_leaf_84_clk_p2c),
    .RESET_B(net1579),
    .D(_01083_),
    .Q_N(_05718_),
    .Q(\shift_storage.storage [442]));
 sg13g2_dfrbp_1 \shift_storage.storage[443]$_SDFFE_PN0P_  (.CLK(clknet_leaf_77_clk_p2c),
    .RESET_B(net1580),
    .D(_01084_),
    .Q_N(_05717_),
    .Q(\shift_storage.storage [443]));
 sg13g2_dfrbp_1 \shift_storage.storage[444]$_SDFFE_PN0P_  (.CLK(clknet_leaf_77_clk_p2c),
    .RESET_B(net1581),
    .D(_01085_),
    .Q_N(_05716_),
    .Q(\shift_storage.storage [444]));
 sg13g2_dfrbp_1 \shift_storage.storage[445]$_SDFFE_PN0P_  (.CLK(clknet_leaf_80_clk_p2c),
    .RESET_B(net1582),
    .D(_01086_),
    .Q_N(_05715_),
    .Q(\shift_storage.storage [445]));
 sg13g2_dfrbp_1 \shift_storage.storage[446]$_SDFFE_PN0P_  (.CLK(clknet_leaf_80_clk_p2c),
    .RESET_B(net1583),
    .D(_01087_),
    .Q_N(_05714_),
    .Q(\shift_storage.storage [446]));
 sg13g2_dfrbp_1 \shift_storage.storage[447]$_SDFFE_PN0P_  (.CLK(clknet_leaf_79_clk_p2c),
    .RESET_B(net1584),
    .D(_01088_),
    .Q_N(_05713_),
    .Q(\shift_storage.storage [447]));
 sg13g2_dfrbp_1 \shift_storage.storage[448]$_SDFFE_PN0P_  (.CLK(clknet_leaf_79_clk_p2c),
    .RESET_B(net1585),
    .D(_01089_),
    .Q_N(_05712_),
    .Q(\shift_storage.storage [448]));
 sg13g2_dfrbp_1 \shift_storage.storage[449]$_SDFFE_PN0P_  (.CLK(clknet_leaf_77_clk_p2c),
    .RESET_B(net1586),
    .D(_01090_),
    .Q_N(_05711_),
    .Q(\shift_storage.storage [449]));
 sg13g2_dfrbp_1 \shift_storage.storage[44]$_SDFFE_PN0P_  (.CLK(clknet_leaf_79_clk_p2c),
    .RESET_B(net1587),
    .D(_01091_),
    .Q_N(_05710_),
    .Q(\shift_storage.storage [44]));
 sg13g2_dfrbp_1 \shift_storage.storage[450]$_SDFFE_PN0P_  (.CLK(clknet_leaf_77_clk_p2c),
    .RESET_B(net1588),
    .D(_01092_),
    .Q_N(_05709_),
    .Q(\shift_storage.storage [450]));
 sg13g2_dfrbp_1 \shift_storage.storage[451]$_SDFFE_PN0P_  (.CLK(clknet_leaf_77_clk_p2c),
    .RESET_B(net1589),
    .D(_01093_),
    .Q_N(_05708_),
    .Q(\shift_storage.storage [451]));
 sg13g2_dfrbp_1 \shift_storage.storage[452]$_SDFFE_PN0P_  (.CLK(clknet_leaf_77_clk_p2c),
    .RESET_B(net1590),
    .D(_01094_),
    .Q_N(_05707_),
    .Q(\shift_storage.storage [452]));
 sg13g2_dfrbp_1 \shift_storage.storage[453]$_SDFFE_PN0P_  (.CLK(clknet_leaf_78_clk_p2c),
    .RESET_B(net1591),
    .D(_01095_),
    .Q_N(_05706_),
    .Q(\shift_storage.storage [453]));
 sg13g2_dfrbp_1 \shift_storage.storage[454]$_SDFFE_PN0P_  (.CLK(clknet_leaf_78_clk_p2c),
    .RESET_B(net1592),
    .D(_01096_),
    .Q_N(_05705_),
    .Q(\shift_storage.storage [454]));
 sg13g2_dfrbp_1 \shift_storage.storage[455]$_SDFFE_PN0P_  (.CLK(clknet_leaf_79_clk_p2c),
    .RESET_B(net1593),
    .D(_01097_),
    .Q_N(_05704_),
    .Q(\shift_storage.storage [455]));
 sg13g2_dfrbp_1 \shift_storage.storage[456]$_SDFFE_PN0P_  (.CLK(clknet_leaf_78_clk_p2c),
    .RESET_B(net1594),
    .D(_01098_),
    .Q_N(_05703_),
    .Q(\shift_storage.storage [456]));
 sg13g2_dfrbp_1 \shift_storage.storage[457]$_SDFFE_PN0P_  (.CLK(clknet_leaf_75_clk_p2c),
    .RESET_B(net1595),
    .D(_01099_),
    .Q_N(_05702_),
    .Q(\shift_storage.storage [457]));
 sg13g2_dfrbp_1 \shift_storage.storage[458]$_SDFFE_PN0P_  (.CLK(clknet_leaf_75_clk_p2c),
    .RESET_B(net1596),
    .D(_01100_),
    .Q_N(_05701_),
    .Q(\shift_storage.storage [458]));
 sg13g2_dfrbp_1 \shift_storage.storage[459]$_SDFFE_PN0P_  (.CLK(clknet_leaf_75_clk_p2c),
    .RESET_B(net1597),
    .D(_01101_),
    .Q_N(_05700_),
    .Q(\shift_storage.storage [459]));
 sg13g2_dfrbp_1 \shift_storage.storage[45]$_SDFFE_PN0P_  (.CLK(clknet_leaf_74_clk_p2c),
    .RESET_B(net1598),
    .D(_01102_),
    .Q_N(_05699_),
    .Q(\shift_storage.storage [45]));
 sg13g2_dfrbp_1 \shift_storage.storage[460]$_SDFFE_PN0P_  (.CLK(clknet_leaf_74_clk_p2c),
    .RESET_B(net1599),
    .D(_01103_),
    .Q_N(_05698_),
    .Q(\shift_storage.storage [460]));
 sg13g2_dfrbp_1 \shift_storage.storage[461]$_SDFFE_PN0P_  (.CLK(clknet_leaf_76_clk_p2c),
    .RESET_B(net1600),
    .D(_01104_),
    .Q_N(_05697_),
    .Q(\shift_storage.storage [461]));
 sg13g2_dfrbp_1 \shift_storage.storage[462]$_SDFFE_PN0P_  (.CLK(clknet_leaf_76_clk_p2c),
    .RESET_B(net1601),
    .D(_01105_),
    .Q_N(_05696_),
    .Q(\shift_storage.storage [462]));
 sg13g2_dfrbp_1 \shift_storage.storage[463]$_SDFFE_PN0P_  (.CLK(clknet_leaf_75_clk_p2c),
    .RESET_B(net1602),
    .D(_01106_),
    .Q_N(_05695_),
    .Q(\shift_storage.storage [463]));
 sg13g2_dfrbp_1 \shift_storage.storage[464]$_SDFFE_PN0P_  (.CLK(clknet_leaf_76_clk_p2c),
    .RESET_B(net1603),
    .D(_01107_),
    .Q_N(_05694_),
    .Q(\shift_storage.storage [464]));
 sg13g2_dfrbp_1 \shift_storage.storage[465]$_SDFFE_PN0P_  (.CLK(clknet_leaf_77_clk_p2c),
    .RESET_B(net1604),
    .D(_01108_),
    .Q_N(_05693_),
    .Q(\shift_storage.storage [465]));
 sg13g2_dfrbp_1 \shift_storage.storage[466]$_SDFFE_PN0P_  (.CLK(clknet_leaf_76_clk_p2c),
    .RESET_B(net1605),
    .D(_01109_),
    .Q_N(_05692_),
    .Q(\shift_storage.storage [466]));
 sg13g2_dfrbp_1 \shift_storage.storage[467]$_SDFFE_PN0P_  (.CLK(clknet_leaf_76_clk_p2c),
    .RESET_B(net1606),
    .D(_01110_),
    .Q_N(_05691_),
    .Q(\shift_storage.storage [467]));
 sg13g2_dfrbp_1 \shift_storage.storage[468]$_SDFFE_PN0P_  (.CLK(clknet_leaf_76_clk_p2c),
    .RESET_B(net1607),
    .D(_01111_),
    .Q_N(_05690_),
    .Q(\shift_storage.storage [468]));
 sg13g2_dfrbp_1 \shift_storage.storage[469]$_SDFFE_PN0P_  (.CLK(clknet_leaf_76_clk_p2c),
    .RESET_B(net1608),
    .D(_01112_),
    .Q_N(_05689_),
    .Q(\shift_storage.storage [469]));
 sg13g2_dfrbp_1 \shift_storage.storage[46]$_SDFFE_PN0P_  (.CLK(clknet_leaf_74_clk_p2c),
    .RESET_B(net1609),
    .D(_01113_),
    .Q_N(_05688_),
    .Q(\shift_storage.storage [46]));
 sg13g2_dfrbp_1 \shift_storage.storage[470]$_SDFFE_PN0P_  (.CLK(clknet_leaf_73_clk_p2c),
    .RESET_B(net1610),
    .D(_01114_),
    .Q_N(_05687_),
    .Q(\shift_storage.storage [470]));
 sg13g2_dfrbp_1 \shift_storage.storage[471]$_SDFFE_PN0P_  (.CLK(clknet_leaf_73_clk_p2c),
    .RESET_B(net1611),
    .D(_01115_),
    .Q_N(_05686_),
    .Q(\shift_storage.storage [471]));
 sg13g2_dfrbp_1 \shift_storage.storage[472]$_SDFFE_PN0P_  (.CLK(clknet_leaf_73_clk_p2c),
    .RESET_B(net1612),
    .D(_01116_),
    .Q_N(_05685_),
    .Q(\shift_storage.storage [472]));
 sg13g2_dfrbp_1 \shift_storage.storage[473]$_SDFFE_PN0P_  (.CLK(clknet_leaf_73_clk_p2c),
    .RESET_B(net1613),
    .D(_01117_),
    .Q_N(_05684_),
    .Q(\shift_storage.storage [473]));
 sg13g2_dfrbp_1 \shift_storage.storage[474]$_SDFFE_PN0P_  (.CLK(clknet_leaf_74_clk_p2c),
    .RESET_B(net1614),
    .D(_01118_),
    .Q_N(_05683_),
    .Q(\shift_storage.storage [474]));
 sg13g2_dfrbp_1 \shift_storage.storage[475]$_SDFFE_PN0P_  (.CLK(clknet_leaf_74_clk_p2c),
    .RESET_B(net1615),
    .D(_01119_),
    .Q_N(_05682_),
    .Q(\shift_storage.storage [475]));
 sg13g2_dfrbp_1 \shift_storage.storage[476]$_SDFFE_PN0P_  (.CLK(clknet_leaf_74_clk_p2c),
    .RESET_B(net1616),
    .D(_01120_),
    .Q_N(_05681_),
    .Q(\shift_storage.storage [476]));
 sg13g2_dfrbp_1 \shift_storage.storage[477]$_SDFFE_PN0P_  (.CLK(clknet_leaf_69_clk_p2c),
    .RESET_B(net1617),
    .D(_01121_),
    .Q_N(_05680_),
    .Q(\shift_storage.storage [477]));
 sg13g2_dfrbp_1 \shift_storage.storage[478]$_SDFFE_PN0P_  (.CLK(clknet_leaf_69_clk_p2c),
    .RESET_B(net1618),
    .D(_01122_),
    .Q_N(_05679_),
    .Q(\shift_storage.storage [478]));
 sg13g2_dfrbp_1 \shift_storage.storage[479]$_SDFFE_PN0P_  (.CLK(clknet_leaf_69_clk_p2c),
    .RESET_B(net1619),
    .D(_01123_),
    .Q_N(_05678_),
    .Q(\shift_storage.storage [479]));
 sg13g2_dfrbp_1 \shift_storage.storage[47]$_SDFFE_PN0P_  (.CLK(clknet_leaf_69_clk_p2c),
    .RESET_B(net1620),
    .D(_01124_),
    .Q_N(_05677_),
    .Q(\shift_storage.storage [47]));
 sg13g2_dfrbp_1 \shift_storage.storage[480]$_SDFFE_PN0P_  (.CLK(clknet_leaf_75_clk_p2c),
    .RESET_B(net1621),
    .D(_01125_),
    .Q_N(_05676_),
    .Q(\shift_storage.storage [480]));
 sg13g2_dfrbp_1 \shift_storage.storage[481]$_SDFFE_PN0P_  (.CLK(clknet_leaf_75_clk_p2c),
    .RESET_B(net1622),
    .D(_01126_),
    .Q_N(_05675_),
    .Q(\shift_storage.storage [481]));
 sg13g2_dfrbp_1 \shift_storage.storage[482]$_SDFFE_PN0P_  (.CLK(clknet_leaf_78_clk_p2c),
    .RESET_B(net1623),
    .D(_01127_),
    .Q_N(_05674_),
    .Q(\shift_storage.storage [482]));
 sg13g2_dfrbp_1 \shift_storage.storage[483]$_SDFFE_PN0P_  (.CLK(clknet_leaf_68_clk_p2c),
    .RESET_B(net1624),
    .D(_01128_),
    .Q_N(_05673_),
    .Q(\shift_storage.storage [483]));
 sg13g2_dfrbp_1 \shift_storage.storage[484]$_SDFFE_PN0P_  (.CLK(clknet_leaf_68_clk_p2c),
    .RESET_B(net1625),
    .D(_01129_),
    .Q_N(_05672_),
    .Q(\shift_storage.storage [484]));
 sg13g2_dfrbp_1 \shift_storage.storage[485]$_SDFFE_PN0P_  (.CLK(clknet_leaf_69_clk_p2c),
    .RESET_B(net1626),
    .D(_01130_),
    .Q_N(_05671_),
    .Q(\shift_storage.storage [485]));
 sg13g2_dfrbp_1 \shift_storage.storage[486]$_SDFFE_PN0P_  (.CLK(clknet_leaf_68_clk_p2c),
    .RESET_B(net1627),
    .D(_01131_),
    .Q_N(_05670_),
    .Q(\shift_storage.storage [486]));
 sg13g2_dfrbp_1 \shift_storage.storage[487]$_SDFFE_PN0P_  (.CLK(clknet_leaf_68_clk_p2c),
    .RESET_B(net1628),
    .D(_01132_),
    .Q_N(_05669_),
    .Q(\shift_storage.storage [487]));
 sg13g2_dfrbp_1 \shift_storage.storage[488]$_SDFFE_PN0P_  (.CLK(clknet_leaf_68_clk_p2c),
    .RESET_B(net1629),
    .D(_01133_),
    .Q_N(_05668_),
    .Q(\shift_storage.storage [488]));
 sg13g2_dfrbp_1 \shift_storage.storage[489]$_SDFFE_PN0P_  (.CLK(clknet_leaf_62_clk_p2c),
    .RESET_B(net1630),
    .D(_01134_),
    .Q_N(_05667_),
    .Q(\shift_storage.storage [489]));
 sg13g2_dfrbp_1 \shift_storage.storage[48]$_SDFFE_PN0P_  (.CLK(clknet_leaf_67_clk_p2c),
    .RESET_B(net1631),
    .D(_01135_),
    .Q_N(_05666_),
    .Q(\shift_storage.storage [48]));
 sg13g2_dfrbp_1 \shift_storage.storage[490]$_SDFFE_PN0P_  (.CLK(clknet_leaf_62_clk_p2c),
    .RESET_B(net1632),
    .D(_01136_),
    .Q_N(_05665_),
    .Q(\shift_storage.storage [490]));
 sg13g2_dfrbp_1 \shift_storage.storage[491]$_SDFFE_PN0P_  (.CLK(clknet_leaf_64_clk_p2c),
    .RESET_B(net1633),
    .D(_01137_),
    .Q_N(_05664_),
    .Q(\shift_storage.storage [491]));
 sg13g2_dfrbp_1 \shift_storage.storage[492]$_SDFFE_PN0P_  (.CLK(clknet_leaf_67_clk_p2c),
    .RESET_B(net1634),
    .D(_01138_),
    .Q_N(_05663_),
    .Q(\shift_storage.storage [492]));
 sg13g2_dfrbp_1 \shift_storage.storage[493]$_SDFFE_PN0P_  (.CLK(clknet_leaf_67_clk_p2c),
    .RESET_B(net1635),
    .D(_01139_),
    .Q_N(_05662_),
    .Q(\shift_storage.storage [493]));
 sg13g2_dfrbp_1 \shift_storage.storage[494]$_SDFFE_PN0P_  (.CLK(clknet_leaf_66_clk_p2c),
    .RESET_B(net1636),
    .D(_01140_),
    .Q_N(_05661_),
    .Q(\shift_storage.storage [494]));
 sg13g2_dfrbp_1 \shift_storage.storage[495]$_SDFFE_PN0P_  (.CLK(clknet_leaf_66_clk_p2c),
    .RESET_B(net1637),
    .D(_01141_),
    .Q_N(_05660_),
    .Q(\shift_storage.storage [495]));
 sg13g2_dfrbp_1 \shift_storage.storage[496]$_SDFFE_PN0P_  (.CLK(clknet_leaf_65_clk_p2c),
    .RESET_B(net1638),
    .D(_01142_),
    .Q_N(_05659_),
    .Q(\shift_storage.storage [496]));
 sg13g2_dfrbp_1 \shift_storage.storage[497]$_SDFFE_PN0P_  (.CLK(clknet_leaf_65_clk_p2c),
    .RESET_B(net1639),
    .D(_01143_),
    .Q_N(_05658_),
    .Q(\shift_storage.storage [497]));
 sg13g2_dfrbp_1 \shift_storage.storage[498]$_SDFFE_PN0P_  (.CLK(clknet_leaf_65_clk_p2c),
    .RESET_B(net1640),
    .D(_01144_),
    .Q_N(_05657_),
    .Q(\shift_storage.storage [498]));
 sg13g2_dfrbp_1 \shift_storage.storage[499]$_SDFFE_PN0P_  (.CLK(clknet_leaf_66_clk_p2c),
    .RESET_B(net1641),
    .D(_01145_),
    .Q_N(_05656_),
    .Q(\shift_storage.storage [499]));
 sg13g2_dfrbp_1 \shift_storage.storage[49]$_SDFFE_PN0P_  (.CLK(clknet_leaf_67_clk_p2c),
    .RESET_B(net1642),
    .D(_01146_),
    .Q_N(_05655_),
    .Q(\shift_storage.storage [49]));
 sg13g2_dfrbp_1 \shift_storage.storage[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_65_clk_p2c),
    .RESET_B(net1643),
    .D(_01147_),
    .Q_N(_05654_),
    .Q(\shift_storage.storage [4]));
 sg13g2_dfrbp_1 \shift_storage.storage[500]$_SDFFE_PN0P_  (.CLK(clknet_leaf_66_clk_p2c),
    .RESET_B(net1644),
    .D(_01148_),
    .Q_N(_05653_),
    .Q(\shift_storage.storage [500]));
 sg13g2_dfrbp_1 \shift_storage.storage[501]$_SDFFE_PN0P_  (.CLK(clknet_leaf_66_clk_p2c),
    .RESET_B(net1645),
    .D(_01149_),
    .Q_N(_05652_),
    .Q(\shift_storage.storage [501]));
 sg13g2_dfrbp_1 \shift_storage.storage[502]$_SDFFE_PN0P_  (.CLK(clknet_leaf_66_clk_p2c),
    .RESET_B(net1646),
    .D(_01150_),
    .Q_N(_05651_),
    .Q(\shift_storage.storage [502]));
 sg13g2_dfrbp_1 \shift_storage.storage[503]$_SDFFE_PN0P_  (.CLK(clknet_leaf_70_clk_p2c),
    .RESET_B(net1647),
    .D(_01151_),
    .Q_N(_05650_),
    .Q(\shift_storage.storage [503]));
 sg13g2_dfrbp_1 \shift_storage.storage[504]$_SDFFE_PN0P_  (.CLK(clknet_leaf_67_clk_p2c),
    .RESET_B(net1648),
    .D(_01152_),
    .Q_N(_05649_),
    .Q(\shift_storage.storage [504]));
 sg13g2_dfrbp_1 \shift_storage.storage[505]$_SDFFE_PN0P_  (.CLK(clknet_leaf_70_clk_p2c),
    .RESET_B(net1649),
    .D(_01153_),
    .Q_N(_05648_),
    .Q(\shift_storage.storage [505]));
 sg13g2_dfrbp_1 \shift_storage.storage[506]$_SDFFE_PN0P_  (.CLK(clknet_leaf_70_clk_p2c),
    .RESET_B(net1650),
    .D(_01154_),
    .Q_N(_05647_),
    .Q(\shift_storage.storage [506]));
 sg13g2_dfrbp_1 \shift_storage.storage[507]$_SDFFE_PN0P_  (.CLK(clknet_leaf_70_clk_p2c),
    .RESET_B(net1651),
    .D(_01155_),
    .Q_N(_05646_),
    .Q(\shift_storage.storage [507]));
 sg13g2_dfrbp_1 \shift_storage.storage[508]$_SDFFE_PN0P_  (.CLK(clknet_leaf_69_clk_p2c),
    .RESET_B(net1652),
    .D(_01156_),
    .Q_N(_05645_),
    .Q(\shift_storage.storage [508]));
 sg13g2_dfrbp_1 \shift_storage.storage[509]$_SDFFE_PN0P_  (.CLK(clknet_leaf_70_clk_p2c),
    .RESET_B(net1653),
    .D(_01157_),
    .Q_N(_05644_),
    .Q(\shift_storage.storage [509]));
 sg13g2_dfrbp_1 \shift_storage.storage[50]$_SDFFE_PN0P_  (.CLK(clknet_leaf_70_clk_p2c),
    .RESET_B(net1654),
    .D(_01158_),
    .Q_N(_05643_),
    .Q(\shift_storage.storage [50]));
 sg13g2_dfrbp_1 \shift_storage.storage[510]$_SDFFE_PN0P_  (.CLK(clknet_leaf_71_clk_p2c),
    .RESET_B(net1655),
    .D(_01159_),
    .Q_N(_05642_),
    .Q(\shift_storage.storage [510]));
 sg13g2_dfrbp_1 \shift_storage.storage[511]$_SDFFE_PN0P_  (.CLK(clknet_leaf_71_clk_p2c),
    .RESET_B(net1656),
    .D(_01160_),
    .Q_N(_05641_),
    .Q(\shift_storage.storage [511]));
 sg13g2_dfrbp_1 \shift_storage.storage[512]$_SDFFE_PN0P_  (.CLK(clknet_leaf_71_clk_p2c),
    .RESET_B(net1657),
    .D(_01161_),
    .Q_N(_05640_),
    .Q(\shift_storage.storage [512]));
 sg13g2_dfrbp_1 \shift_storage.storage[513]$_SDFFE_PN0P_  (.CLK(clknet_leaf_73_clk_p2c),
    .RESET_B(net1658),
    .D(_01162_),
    .Q_N(_05639_),
    .Q(\shift_storage.storage [513]));
 sg13g2_dfrbp_1 \shift_storage.storage[514]$_SDFFE_PN0P_  (.CLK(clknet_leaf_73_clk_p2c),
    .RESET_B(net1659),
    .D(_01163_),
    .Q_N(_05638_),
    .Q(\shift_storage.storage [514]));
 sg13g2_dfrbp_1 \shift_storage.storage[515]$_SDFFE_PN0P_  (.CLK(clknet_leaf_72_clk_p2c),
    .RESET_B(net1660),
    .D(_01164_),
    .Q_N(_05637_),
    .Q(\shift_storage.storage [515]));
 sg13g2_dfrbp_1 \shift_storage.storage[516]$_SDFFE_PN0P_  (.CLK(clknet_leaf_72_clk_p2c),
    .RESET_B(net1661),
    .D(_01165_),
    .Q_N(_05636_),
    .Q(\shift_storage.storage [516]));
 sg13g2_dfrbp_1 \shift_storage.storage[517]$_SDFFE_PN0P_  (.CLK(clknet_leaf_72_clk_p2c),
    .RESET_B(net1662),
    .D(_01166_),
    .Q_N(_05635_),
    .Q(\shift_storage.storage [517]));
 sg13g2_dfrbp_1 \shift_storage.storage[518]$_SDFFE_PN0P_  (.CLK(clknet_leaf_72_clk_p2c),
    .RESET_B(net1663),
    .D(_01167_),
    .Q_N(_05634_),
    .Q(\shift_storage.storage [518]));
 sg13g2_dfrbp_1 \shift_storage.storage[519]$_SDFFE_PN0P_  (.CLK(clknet_leaf_72_clk_p2c),
    .RESET_B(net1664),
    .D(_01168_),
    .Q_N(_05633_),
    .Q(\shift_storage.storage [519]));
 sg13g2_dfrbp_1 \shift_storage.storage[51]$_SDFFE_PN0P_  (.CLK(clknet_leaf_71_clk_p2c),
    .RESET_B(net1665),
    .D(_01169_),
    .Q_N(_05632_),
    .Q(\shift_storage.storage [51]));
 sg13g2_dfrbp_1 \shift_storage.storage[520]$_SDFFE_PN0P_  (.CLK(clknet_leaf_72_clk_p2c),
    .RESET_B(net1666),
    .D(_01170_),
    .Q_N(_05631_),
    .Q(\shift_storage.storage [520]));
 sg13g2_dfrbp_1 \shift_storage.storage[521]$_SDFFE_PN0P_  (.CLK(clknet_leaf_71_clk_p2c),
    .RESET_B(net1667),
    .D(_01171_),
    .Q_N(_05630_),
    .Q(\shift_storage.storage [521]));
 sg13g2_dfrbp_1 \shift_storage.storage[522]$_SDFFE_PN0P_  (.CLK(clknet_leaf_71_clk_p2c),
    .RESET_B(net1668),
    .D(_01172_),
    .Q_N(_05629_),
    .Q(\shift_storage.storage [522]));
 sg13g2_dfrbp_1 \shift_storage.storage[523]$_SDFFE_PN0P_  (.CLK(clknet_leaf_24_clk_p2c),
    .RESET_B(net1669),
    .D(_01173_),
    .Q_N(_05628_),
    .Q(\shift_storage.storage [523]));
 sg13g2_dfrbp_1 \shift_storage.storage[524]$_SDFFE_PN0P_  (.CLK(clknet_leaf_24_clk_p2c),
    .RESET_B(net1670),
    .D(_01174_),
    .Q_N(_05627_),
    .Q(\shift_storage.storage [524]));
 sg13g2_dfrbp_1 \shift_storage.storage[525]$_SDFFE_PN0P_  (.CLK(clknet_leaf_23_clk_p2c),
    .RESET_B(net1671),
    .D(_01175_),
    .Q_N(_05626_),
    .Q(\shift_storage.storage [525]));
 sg13g2_dfrbp_1 \shift_storage.storage[526]$_SDFFE_PN0P_  (.CLK(clknet_leaf_23_clk_p2c),
    .RESET_B(net1672),
    .D(_01176_),
    .Q_N(_05625_),
    .Q(\shift_storage.storage [526]));
 sg13g2_dfrbp_1 \shift_storage.storage[527]$_SDFFE_PN0P_  (.CLK(clknet_leaf_24_clk_p2c),
    .RESET_B(net1673),
    .D(_01177_),
    .Q_N(_05624_),
    .Q(\shift_storage.storage [527]));
 sg13g2_dfrbp_1 \shift_storage.storage[528]$_SDFFE_PN0P_  (.CLK(clknet_leaf_24_clk_p2c),
    .RESET_B(net1674),
    .D(_01178_),
    .Q_N(_05623_),
    .Q(\shift_storage.storage [528]));
 sg13g2_dfrbp_1 \shift_storage.storage[529]$_SDFFE_PN0P_  (.CLK(clknet_leaf_25_clk_p2c),
    .RESET_B(net1675),
    .D(_01179_),
    .Q_N(_05622_),
    .Q(\shift_storage.storage [529]));
 sg13g2_dfrbp_1 \shift_storage.storage[52]$_SDFFE_PN0P_  (.CLK(clknet_leaf_25_clk_p2c),
    .RESET_B(net1676),
    .D(_01180_),
    .Q_N(_05621_),
    .Q(\shift_storage.storage [52]));
 sg13g2_dfrbp_1 \shift_storage.storage[530]$_SDFFE_PN0P_  (.CLK(clknet_leaf_25_clk_p2c),
    .RESET_B(net1677),
    .D(_01181_),
    .Q_N(_05620_),
    .Q(\shift_storage.storage [530]));
 sg13g2_dfrbp_1 \shift_storage.storage[531]$_SDFFE_PN0P_  (.CLK(clknet_leaf_25_clk_p2c),
    .RESET_B(net1678),
    .D(_01182_),
    .Q_N(_05619_),
    .Q(\shift_storage.storage [531]));
 sg13g2_dfrbp_1 \shift_storage.storage[532]$_SDFFE_PN0P_  (.CLK(clknet_leaf_25_clk_p2c),
    .RESET_B(net1679),
    .D(_01183_),
    .Q_N(_05618_),
    .Q(\shift_storage.storage [532]));
 sg13g2_dfrbp_1 \shift_storage.storage[533]$_SDFFE_PN0P_  (.CLK(clknet_leaf_26_clk_p2c),
    .RESET_B(net1680),
    .D(_01184_),
    .Q_N(_05617_),
    .Q(\shift_storage.storage [533]));
 sg13g2_dfrbp_1 \shift_storage.storage[534]$_SDFFE_PN0P_  (.CLK(clknet_leaf_25_clk_p2c),
    .RESET_B(net1681),
    .D(_01185_),
    .Q_N(_05616_),
    .Q(\shift_storage.storage [534]));
 sg13g2_dfrbp_1 \shift_storage.storage[535]$_SDFFE_PN0P_  (.CLK(clknet_leaf_25_clk_p2c),
    .RESET_B(net1682),
    .D(_01186_),
    .Q_N(_05615_),
    .Q(\shift_storage.storage [535]));
 sg13g2_dfrbp_1 \shift_storage.storage[536]$_SDFFE_PN0P_  (.CLK(clknet_leaf_28_clk_p2c),
    .RESET_B(net1683),
    .D(_01187_),
    .Q_N(_05614_),
    .Q(\shift_storage.storage [536]));
 sg13g2_dfrbp_1 \shift_storage.storage[537]$_SDFFE_PN0P_  (.CLK(clknet_leaf_28_clk_p2c),
    .RESET_B(net1684),
    .D(_01188_),
    .Q_N(_05613_),
    .Q(\shift_storage.storage [537]));
 sg13g2_dfrbp_1 \shift_storage.storage[538]$_SDFFE_PN0P_  (.CLK(clknet_leaf_29_clk_p2c),
    .RESET_B(net1685),
    .D(_01189_),
    .Q_N(_05612_),
    .Q(\shift_storage.storage [538]));
 sg13g2_dfrbp_1 \shift_storage.storage[539]$_SDFFE_PN0P_  (.CLK(clknet_leaf_29_clk_p2c),
    .RESET_B(net1686),
    .D(_01190_),
    .Q_N(_05611_),
    .Q(\shift_storage.storage [539]));
 sg13g2_dfrbp_1 \shift_storage.storage[53]$_SDFFE_PN0P_  (.CLK(clknet_leaf_28_clk_p2c),
    .RESET_B(net1687),
    .D(_01191_),
    .Q_N(_05610_),
    .Q(\shift_storage.storage [53]));
 sg13g2_dfrbp_1 \shift_storage.storage[540]$_SDFFE_PN0P_  (.CLK(clknet_leaf_29_clk_p2c),
    .RESET_B(net1688),
    .D(_01192_),
    .Q_N(_05609_),
    .Q(\shift_storage.storage [540]));
 sg13g2_dfrbp_1 \shift_storage.storage[541]$_SDFFE_PN0P_  (.CLK(clknet_leaf_28_clk_p2c),
    .RESET_B(net1689),
    .D(_01193_),
    .Q_N(_05608_),
    .Q(\shift_storage.storage [541]));
 sg13g2_dfrbp_1 \shift_storage.storage[542]$_SDFFE_PN0P_  (.CLK(clknet_leaf_28_clk_p2c),
    .RESET_B(net1690),
    .D(_01194_),
    .Q_N(_05607_),
    .Q(\shift_storage.storage [542]));
 sg13g2_dfrbp_1 \shift_storage.storage[543]$_SDFFE_PN0P_  (.CLK(clknet_leaf_28_clk_p2c),
    .RESET_B(net1691),
    .D(_01195_),
    .Q_N(_05606_),
    .Q(\shift_storage.storage [543]));
 sg13g2_dfrbp_1 \shift_storage.storage[544]$_SDFFE_PN0P_  (.CLK(clknet_leaf_32_clk_p2c),
    .RESET_B(net1692),
    .D(_01196_),
    .Q_N(_05605_),
    .Q(\shift_storage.storage [544]));
 sg13g2_dfrbp_1 \shift_storage.storage[545]$_SDFFE_PN0P_  (.CLK(clknet_leaf_33_clk_p2c),
    .RESET_B(net1693),
    .D(_01197_),
    .Q_N(_05604_),
    .Q(\shift_storage.storage [545]));
 sg13g2_dfrbp_1 \shift_storage.storage[546]$_SDFFE_PN0P_  (.CLK(clknet_leaf_33_clk_p2c),
    .RESET_B(net1694),
    .D(_01198_),
    .Q_N(_05603_),
    .Q(\shift_storage.storage [546]));
 sg13g2_dfrbp_1 \shift_storage.storage[547]$_SDFFE_PN0P_  (.CLK(clknet_leaf_27_clk_p2c),
    .RESET_B(net1695),
    .D(_01199_),
    .Q_N(_05602_),
    .Q(\shift_storage.storage [547]));
 sg13g2_dfrbp_1 \shift_storage.storage[548]$_SDFFE_PN0P_  (.CLK(clknet_leaf_27_clk_p2c),
    .RESET_B(net1696),
    .D(_01200_),
    .Q_N(_05601_),
    .Q(\shift_storage.storage [548]));
 sg13g2_dfrbp_1 \shift_storage.storage[549]$_SDFFE_PN0P_  (.CLK(clknet_leaf_27_clk_p2c),
    .RESET_B(net1697),
    .D(_01201_),
    .Q_N(_05600_),
    .Q(\shift_storage.storage [549]));
 sg13g2_dfrbp_1 \shift_storage.storage[54]$_SDFFE_PN0P_  (.CLK(clknet_leaf_27_clk_p2c),
    .RESET_B(net1698),
    .D(_01202_),
    .Q_N(_05599_),
    .Q(\shift_storage.storage [54]));
 sg13g2_dfrbp_1 \shift_storage.storage[550]$_SDFFE_PN0P_  (.CLK(clknet_leaf_26_clk_p2c),
    .RESET_B(net1699),
    .D(_01203_),
    .Q_N(_05598_),
    .Q(\shift_storage.storage [550]));
 sg13g2_dfrbp_1 \shift_storage.storage[551]$_SDFFE_PN0P_  (.CLK(clknet_leaf_26_clk_p2c),
    .RESET_B(net1700),
    .D(_01204_),
    .Q_N(_05597_),
    .Q(\shift_storage.storage [551]));
 sg13g2_dfrbp_1 \shift_storage.storage[552]$_SDFFE_PN0P_  (.CLK(clknet_leaf_26_clk_p2c),
    .RESET_B(net1701),
    .D(_01205_),
    .Q_N(_05596_),
    .Q(\shift_storage.storage [552]));
 sg13g2_dfrbp_1 \shift_storage.storage[553]$_SDFFE_PN0P_  (.CLK(clknet_leaf_27_clk_p2c),
    .RESET_B(net1702),
    .D(_01206_),
    .Q_N(_05595_),
    .Q(\shift_storage.storage [553]));
 sg13g2_dfrbp_1 \shift_storage.storage[554]$_SDFFE_PN0P_  (.CLK(clknet_leaf_26_clk_p2c),
    .RESET_B(net1703),
    .D(_01207_),
    .Q_N(_05594_),
    .Q(\shift_storage.storage [554]));
 sg13g2_dfrbp_1 \shift_storage.storage[555]$_SDFFE_PN0P_  (.CLK(clknet_leaf_21_clk_p2c),
    .RESET_B(net1704),
    .D(_01208_),
    .Q_N(_05593_),
    .Q(\shift_storage.storage [555]));
 sg13g2_dfrbp_1 \shift_storage.storage[556]$_SDFFE_PN0P_  (.CLK(clknet_leaf_21_clk_p2c),
    .RESET_B(net1705),
    .D(_01209_),
    .Q_N(_05592_),
    .Q(\shift_storage.storage [556]));
 sg13g2_dfrbp_1 \shift_storage.storage[557]$_SDFFE_PN0P_  (.CLK(clknet_leaf_21_clk_p2c),
    .RESET_B(net1706),
    .D(_01210_),
    .Q_N(_05591_),
    .Q(\shift_storage.storage [557]));
 sg13g2_dfrbp_1 \shift_storage.storage[558]$_SDFFE_PN0P_  (.CLK(clknet_leaf_23_clk_p2c),
    .RESET_B(net1707),
    .D(_01211_),
    .Q_N(_05590_),
    .Q(\shift_storage.storage [558]));
 sg13g2_dfrbp_1 \shift_storage.storage[559]$_SDFFE_PN0P_  (.CLK(clknet_leaf_21_clk_p2c),
    .RESET_B(net1708),
    .D(_01212_),
    .Q_N(_05589_),
    .Q(\shift_storage.storage [559]));
 sg13g2_dfrbp_1 \shift_storage.storage[55]$_SDFFE_PN0P_  (.CLK(clknet_leaf_20_clk_p2c),
    .RESET_B(net1709),
    .D(_01213_),
    .Q_N(_05588_),
    .Q(\shift_storage.storage [55]));
 sg13g2_dfrbp_1 \shift_storage.storage[560]$_SDFFE_PN0P_  (.CLK(clknet_leaf_24_clk_p2c),
    .RESET_B(net1710),
    .D(_01214_),
    .Q_N(_05587_),
    .Q(\shift_storage.storage [560]));
 sg13g2_dfrbp_1 \shift_storage.storage[561]$_SDFFE_PN0P_  (.CLK(clknet_leaf_23_clk_p2c),
    .RESET_B(net1711),
    .D(_01215_),
    .Q_N(_05586_),
    .Q(\shift_storage.storage [561]));
 sg13g2_dfrbp_1 \shift_storage.storage[562]$_SDFFE_PN0P_  (.CLK(clknet_leaf_23_clk_p2c),
    .RESET_B(net1712),
    .D(_01216_),
    .Q_N(_05585_),
    .Q(\shift_storage.storage [562]));
 sg13g2_dfrbp_1 \shift_storage.storage[563]$_SDFFE_PN0P_  (.CLK(clknet_leaf_22_clk_p2c),
    .RESET_B(net1713),
    .D(_01217_),
    .Q_N(_05584_),
    .Q(\shift_storage.storage [563]));
 sg13g2_dfrbp_1 \shift_storage.storage[564]$_SDFFE_PN0P_  (.CLK(clknet_leaf_22_clk_p2c),
    .RESET_B(net1714),
    .D(_01218_),
    .Q_N(_05583_),
    .Q(\shift_storage.storage [564]));
 sg13g2_dfrbp_1 \shift_storage.storage[565]$_SDFFE_PN0P_  (.CLK(clknet_leaf_22_clk_p2c),
    .RESET_B(net1715),
    .D(_01219_),
    .Q_N(_05582_),
    .Q(\shift_storage.storage [565]));
 sg13g2_dfrbp_1 \shift_storage.storage[566]$_SDFFE_PN0P_  (.CLK(clknet_leaf_22_clk_p2c),
    .RESET_B(net1716),
    .D(_01220_),
    .Q_N(_05581_),
    .Q(\shift_storage.storage [566]));
 sg13g2_dfrbp_1 \shift_storage.storage[567]$_SDFFE_PN0P_  (.CLK(clknet_leaf_22_clk_p2c),
    .RESET_B(net1717),
    .D(_01221_),
    .Q_N(_05580_),
    .Q(\shift_storage.storage [567]));
 sg13g2_dfrbp_1 \shift_storage.storage[568]$_SDFFE_PN0P_  (.CLK(clknet_leaf_22_clk_p2c),
    .RESET_B(net1718),
    .D(_01222_),
    .Q_N(_05579_),
    .Q(\shift_storage.storage [568]));
 sg13g2_dfrbp_1 \shift_storage.storage[569]$_SDFFE_PN0P_  (.CLK(clknet_leaf_19_clk_p2c),
    .RESET_B(net1719),
    .D(_01223_),
    .Q_N(_05578_),
    .Q(\shift_storage.storage [569]));
 sg13g2_dfrbp_1 \shift_storage.storage[56]$_SDFFE_PN0P_  (.CLK(clknet_leaf_20_clk_p2c),
    .RESET_B(net1720),
    .D(_01224_),
    .Q_N(_05577_),
    .Q(\shift_storage.storage [56]));
 sg13g2_dfrbp_1 \shift_storage.storage[570]$_SDFFE_PN0P_  (.CLK(clknet_leaf_19_clk_p2c),
    .RESET_B(net1721),
    .D(_01225_),
    .Q_N(_05576_),
    .Q(\shift_storage.storage [570]));
 sg13g2_dfrbp_1 \shift_storage.storage[571]$_SDFFE_PN0P_  (.CLK(clknet_leaf_19_clk_p2c),
    .RESET_B(net1722),
    .D(_01226_),
    .Q_N(_05575_),
    .Q(\shift_storage.storage [571]));
 sg13g2_dfrbp_1 \shift_storage.storage[572]$_SDFFE_PN0P_  (.CLK(clknet_leaf_19_clk_p2c),
    .RESET_B(net1723),
    .D(_01227_),
    .Q_N(_05574_),
    .Q(\shift_storage.storage [572]));
 sg13g2_dfrbp_1 \shift_storage.storage[573]$_SDFFE_PN0P_  (.CLK(clknet_leaf_19_clk_p2c),
    .RESET_B(net1724),
    .D(_01228_),
    .Q_N(_05573_),
    .Q(\shift_storage.storage [573]));
 sg13g2_dfrbp_1 \shift_storage.storage[574]$_SDFFE_PN0P_  (.CLK(clknet_leaf_20_clk_p2c),
    .RESET_B(net1725),
    .D(_01229_),
    .Q_N(_05572_),
    .Q(\shift_storage.storage [574]));
 sg13g2_dfrbp_1 \shift_storage.storage[575]$_SDFFE_PN0P_  (.CLK(clknet_leaf_19_clk_p2c),
    .RESET_B(net1726),
    .D(_01230_),
    .Q_N(_05571_),
    .Q(\shift_storage.storage [575]));
 sg13g2_dfrbp_1 \shift_storage.storage[576]$_SDFFE_PN0P_  (.CLK(clknet_leaf_20_clk_p2c),
    .RESET_B(net1727),
    .D(_01231_),
    .Q_N(_05570_),
    .Q(\shift_storage.storage [576]));
 sg13g2_dfrbp_1 \shift_storage.storage[577]$_SDFFE_PN0P_  (.CLK(clknet_leaf_20_clk_p2c),
    .RESET_B(net1728),
    .D(_01232_),
    .Q_N(_05569_),
    .Q(\shift_storage.storage [577]));
 sg13g2_dfrbp_1 \shift_storage.storage[578]$_SDFFE_PN0P_  (.CLK(clknet_leaf_15_clk_p2c),
    .RESET_B(net1729),
    .D(_01233_),
    .Q_N(_05568_),
    .Q(\shift_storage.storage [578]));
 sg13g2_dfrbp_1 \shift_storage.storage[579]$_SDFFE_PN0P_  (.CLK(clknet_leaf_15_clk_p2c),
    .RESET_B(net1730),
    .D(_01234_),
    .Q_N(_05567_),
    .Q(\shift_storage.storage [579]));
 sg13g2_dfrbp_1 \shift_storage.storage[57]$_SDFFE_PN0P_  (.CLK(clknet_leaf_20_clk_p2c),
    .RESET_B(net1731),
    .D(_01235_),
    .Q_N(_05566_),
    .Q(\shift_storage.storage [57]));
 sg13g2_dfrbp_1 \shift_storage.storage[580]$_SDFFE_PN0P_  (.CLK(clknet_leaf_15_clk_p2c),
    .RESET_B(net1732),
    .D(_01236_),
    .Q_N(_05565_),
    .Q(\shift_storage.storage [580]));
 sg13g2_dfrbp_1 \shift_storage.storage[581]$_SDFFE_PN0P_  (.CLK(clknet_leaf_15_clk_p2c),
    .RESET_B(net1733),
    .D(_01237_),
    .Q_N(_05564_),
    .Q(\shift_storage.storage [581]));
 sg13g2_dfrbp_1 \shift_storage.storage[582]$_SDFFE_PN0P_  (.CLK(clknet_leaf_14_clk_p2c),
    .RESET_B(net1734),
    .D(_01238_),
    .Q_N(_05563_),
    .Q(\shift_storage.storage [582]));
 sg13g2_dfrbp_1 \shift_storage.storage[583]$_SDFFE_PN0P_  (.CLK(clknet_leaf_14_clk_p2c),
    .RESET_B(net1735),
    .D(_01239_),
    .Q_N(_05562_),
    .Q(\shift_storage.storage [583]));
 sg13g2_dfrbp_1 \shift_storage.storage[584]$_SDFFE_PN0P_  (.CLK(clknet_leaf_14_clk_p2c),
    .RESET_B(net1736),
    .D(_01240_),
    .Q_N(_05561_),
    .Q(\shift_storage.storage [584]));
 sg13g2_dfrbp_1 \shift_storage.storage[585]$_SDFFE_PN0P_  (.CLK(clknet_leaf_21_clk_p2c),
    .RESET_B(net1737),
    .D(_01241_),
    .Q_N(_05560_),
    .Q(\shift_storage.storage [585]));
 sg13g2_dfrbp_1 \shift_storage.storage[586]$_SDFFE_PN0P_  (.CLK(clknet_leaf_21_clk_p2c),
    .RESET_B(net1738),
    .D(_01242_),
    .Q_N(_05559_),
    .Q(\shift_storage.storage [586]));
 sg13g2_dfrbp_1 \shift_storage.storage[587]$_SDFFE_PN0P_  (.CLK(clknet_leaf_33_clk_p2c),
    .RESET_B(net1739),
    .D(_01243_),
    .Q_N(_05558_),
    .Q(\shift_storage.storage [587]));
 sg13g2_dfrbp_1 \shift_storage.storage[588]$_SDFFE_PN0P_  (.CLK(clknet_leaf_33_clk_p2c),
    .RESET_B(net1740),
    .D(_01244_),
    .Q_N(_05557_),
    .Q(\shift_storage.storage [588]));
 sg13g2_dfrbp_1 \shift_storage.storage[589]$_SDFFE_PN0P_  (.CLK(clknet_leaf_33_clk_p2c),
    .RESET_B(net1741),
    .D(_01245_),
    .Q_N(_05556_),
    .Q(\shift_storage.storage [589]));
 sg13g2_dfrbp_1 \shift_storage.storage[58]$_SDFFE_PN0P_  (.CLK(clknet_leaf_14_clk_p2c),
    .RESET_B(net1742),
    .D(_01246_),
    .Q_N(_05555_),
    .Q(\shift_storage.storage [58]));
 sg13g2_dfrbp_1 \shift_storage.storage[590]$_SDFFE_PN0P_  (.CLK(clknet_leaf_33_clk_p2c),
    .RESET_B(net1743),
    .D(_01247_),
    .Q_N(_05554_),
    .Q(\shift_storage.storage [590]));
 sg13g2_dfrbp_1 \shift_storage.storage[591]$_SDFFE_PN0P_  (.CLK(clknet_leaf_34_clk_p2c),
    .RESET_B(net1744),
    .D(_01248_),
    .Q_N(_05553_),
    .Q(\shift_storage.storage [591]));
 sg13g2_dfrbp_1 \shift_storage.storage[592]$_SDFFE_PN0P_  (.CLK(clknet_leaf_13_clk_p2c),
    .RESET_B(net1745),
    .D(_01249_),
    .Q_N(_05552_),
    .Q(\shift_storage.storage [592]));
 sg13g2_dfrbp_1 \shift_storage.storage[593]$_SDFFE_PN0P_  (.CLK(clknet_leaf_34_clk_p2c),
    .RESET_B(net1746),
    .D(_01250_),
    .Q_N(_05551_),
    .Q(\shift_storage.storage [593]));
 sg13g2_dfrbp_1 \shift_storage.storage[594]$_SDFFE_PN0P_  (.CLK(clknet_leaf_14_clk_p2c),
    .RESET_B(net1747),
    .D(_01251_),
    .Q_N(_05550_),
    .Q(\shift_storage.storage [594]));
 sg13g2_dfrbp_1 \shift_storage.storage[595]$_SDFFE_PN0P_  (.CLK(clknet_leaf_14_clk_p2c),
    .RESET_B(net1748),
    .D(_01252_),
    .Q_N(_05549_),
    .Q(\shift_storage.storage [595]));
 sg13g2_dfrbp_1 \shift_storage.storage[596]$_SDFFE_PN0P_  (.CLK(clknet_leaf_13_clk_p2c),
    .RESET_B(net1749),
    .D(_01253_),
    .Q_N(_05548_),
    .Q(\shift_storage.storage [596]));
 sg13g2_dfrbp_1 \shift_storage.storage[597]$_SDFFE_PN0P_  (.CLK(clknet_leaf_13_clk_p2c),
    .RESET_B(net1750),
    .D(_01254_),
    .Q_N(_05547_),
    .Q(\shift_storage.storage [597]));
 sg13g2_dfrbp_1 \shift_storage.storage[598]$_SDFFE_PN0P_  (.CLK(clknet_leaf_13_clk_p2c),
    .RESET_B(net1751),
    .D(_01255_),
    .Q_N(_05546_),
    .Q(\shift_storage.storage [598]));
 sg13g2_dfrbp_1 \shift_storage.storage[599]$_SDFFE_PN0P_  (.CLK(clknet_leaf_12_clk_p2c),
    .RESET_B(net1752),
    .D(_01256_),
    .Q_N(_05545_),
    .Q(\shift_storage.storage [599]));
 sg13g2_dfrbp_1 \shift_storage.storage[59]$_SDFFE_PN0P_  (.CLK(clknet_leaf_15_clk_p2c),
    .RESET_B(net1753),
    .D(_01257_),
    .Q_N(_05544_),
    .Q(\shift_storage.storage [59]));
 sg13g2_dfrbp_1 \shift_storage.storage[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_35_clk_p2c),
    .RESET_B(net1754),
    .D(_01258_),
    .Q_N(_05543_),
    .Q(\shift_storage.storage [5]));
 sg13g2_dfrbp_1 \shift_storage.storage[600]$_SDFFE_PN0P_  (.CLK(clknet_leaf_12_clk_p2c),
    .RESET_B(net1755),
    .D(_01259_),
    .Q_N(_05542_),
    .Q(\shift_storage.storage [600]));
 sg13g2_dfrbp_1 \shift_storage.storage[601]$_SDFFE_PN0P_  (.CLK(clknet_leaf_12_clk_p2c),
    .RESET_B(net1756),
    .D(_01260_),
    .Q_N(_05541_),
    .Q(\shift_storage.storage [601]));
 sg13g2_dfrbp_1 \shift_storage.storage[602]$_SDFFE_PN0P_  (.CLK(clknet_leaf_12_clk_p2c),
    .RESET_B(net1757),
    .D(_01261_),
    .Q_N(_05540_),
    .Q(\shift_storage.storage [602]));
 sg13g2_dfrbp_1 \shift_storage.storage[603]$_SDFFE_PN0P_  (.CLK(clknet_leaf_11_clk_p2c),
    .RESET_B(net1758),
    .D(_01262_),
    .Q_N(_05539_),
    .Q(\shift_storage.storage [603]));
 sg13g2_dfrbp_1 \shift_storage.storage[604]$_SDFFE_PN0P_  (.CLK(clknet_leaf_10_clk_p2c),
    .RESET_B(net1759),
    .D(_01263_),
    .Q_N(_05538_),
    .Q(\shift_storage.storage [604]));
 sg13g2_dfrbp_1 \shift_storage.storage[605]$_SDFFE_PN0P_  (.CLK(clknet_leaf_10_clk_p2c),
    .RESET_B(net1760),
    .D(_01264_),
    .Q_N(_05537_),
    .Q(\shift_storage.storage [605]));
 sg13g2_dfrbp_1 \shift_storage.storage[606]$_SDFFE_PN0P_  (.CLK(clknet_leaf_13_clk_p2c),
    .RESET_B(net1761),
    .D(_01265_),
    .Q_N(_05536_),
    .Q(\shift_storage.storage [606]));
 sg13g2_dfrbp_1 \shift_storage.storage[607]$_SDFFE_PN0P_  (.CLK(clknet_leaf_12_clk_p2c),
    .RESET_B(net1762),
    .D(_01266_),
    .Q_N(_05535_),
    .Q(\shift_storage.storage [607]));
 sg13g2_dfrbp_1 \shift_storage.storage[608]$_SDFFE_PN0P_  (.CLK(clknet_leaf_13_clk_p2c),
    .RESET_B(net1763),
    .D(_01267_),
    .Q_N(_05534_),
    .Q(\shift_storage.storage [608]));
 sg13g2_dfrbp_1 \shift_storage.storage[609]$_SDFFE_PN0P_  (.CLK(clknet_leaf_16_clk_p2c),
    .RESET_B(net1764),
    .D(_01268_),
    .Q_N(_05533_),
    .Q(\shift_storage.storage [609]));
 sg13g2_dfrbp_1 \shift_storage.storage[60]$_SDFFE_PN0P_  (.CLK(clknet_leaf_16_clk_p2c),
    .RESET_B(net1765),
    .D(_01269_),
    .Q_N(_05532_),
    .Q(\shift_storage.storage [60]));
 sg13g2_dfrbp_1 \shift_storage.storage[610]$_SDFFE_PN0P_  (.CLK(clknet_leaf_10_clk_p2c),
    .RESET_B(net1766),
    .D(_01270_),
    .Q_N(_05531_),
    .Q(\shift_storage.storage [610]));
 sg13g2_dfrbp_1 \shift_storage.storage[611]$_SDFFE_PN0P_  (.CLK(clknet_leaf_7_clk_p2c),
    .RESET_B(net1767),
    .D(_01271_),
    .Q_N(_05530_),
    .Q(\shift_storage.storage [611]));
 sg13g2_dfrbp_1 \shift_storage.storage[612]$_SDFFE_PN0P_  (.CLK(clknet_leaf_7_clk_p2c),
    .RESET_B(net1768),
    .D(_01272_),
    .Q_N(_05529_),
    .Q(\shift_storage.storage [612]));
 sg13g2_dfrbp_1 \shift_storage.storage[613]$_SDFFE_PN0P_  (.CLK(clknet_leaf_7_clk_p2c),
    .RESET_B(net1769),
    .D(_01273_),
    .Q_N(_05528_),
    .Q(\shift_storage.storage [613]));
 sg13g2_dfrbp_1 \shift_storage.storage[614]$_SDFFE_PN0P_  (.CLK(clknet_leaf_7_clk_p2c),
    .RESET_B(net1770),
    .D(_01274_),
    .Q_N(_05527_),
    .Q(\shift_storage.storage [614]));
 sg13g2_dfrbp_1 \shift_storage.storage[615]$_SDFFE_PN0P_  (.CLK(clknet_leaf_6_clk_p2c),
    .RESET_B(net1771),
    .D(_01275_),
    .Q_N(_05526_),
    .Q(\shift_storage.storage [615]));
 sg13g2_dfrbp_1 \shift_storage.storage[616]$_SDFFE_PN0P_  (.CLK(clknet_leaf_6_clk_p2c),
    .RESET_B(net1772),
    .D(_01276_),
    .Q_N(_05525_),
    .Q(\shift_storage.storage [616]));
 sg13g2_dfrbp_1 \shift_storage.storage[617]$_SDFFE_PN0P_  (.CLK(clknet_leaf_16_clk_p2c),
    .RESET_B(net1773),
    .D(_01277_),
    .Q_N(_05524_),
    .Q(\shift_storage.storage [617]));
 sg13g2_dfrbp_1 \shift_storage.storage[618]$_SDFFE_PN0P_  (.CLK(clknet_leaf_16_clk_p2c),
    .RESET_B(net1774),
    .D(_01278_),
    .Q_N(_05523_),
    .Q(\shift_storage.storage [618]));
 sg13g2_dfrbp_1 \shift_storage.storage[619]$_SDFFE_PN0P_  (.CLK(clknet_leaf_15_clk_p2c),
    .RESET_B(net1775),
    .D(_01279_),
    .Q_N(_05522_),
    .Q(\shift_storage.storage [619]));
 sg13g2_dfrbp_1 \shift_storage.storage[61]$_SDFFE_PN0P_  (.CLK(clknet_leaf_17_clk_p2c),
    .RESET_B(net1776),
    .D(_01280_),
    .Q_N(_05521_),
    .Q(\shift_storage.storage [61]));
 sg13g2_dfrbp_1 \shift_storage.storage[620]$_SDFFE_PN0P_  (.CLK(clknet_leaf_16_clk_p2c),
    .RESET_B(net1777),
    .D(_01281_),
    .Q_N(_05520_),
    .Q(\shift_storage.storage [620]));
 sg13g2_dfrbp_1 \shift_storage.storage[621]$_SDFFE_PN0P_  (.CLK(clknet_leaf_17_clk_p2c),
    .RESET_B(net1778),
    .D(_01282_),
    .Q_N(_05519_),
    .Q(\shift_storage.storage [621]));
 sg13g2_dfrbp_1 \shift_storage.storage[622]$_SDFFE_PN0P_  (.CLK(clknet_leaf_17_clk_p2c),
    .RESET_B(net1779),
    .D(_01283_),
    .Q_N(_05518_),
    .Q(\shift_storage.storage [622]));
 sg13g2_dfrbp_1 \shift_storage.storage[623]$_SDFFE_PN0P_  (.CLK(clknet_leaf_18_clk_p2c),
    .RESET_B(net1780),
    .D(_01284_),
    .Q_N(_05517_),
    .Q(\shift_storage.storage [623]));
 sg13g2_dfrbp_1 \shift_storage.storage[624]$_SDFFE_PN0P_  (.CLK(clknet_leaf_18_clk_p2c),
    .RESET_B(net1781),
    .D(_01285_),
    .Q_N(_05516_),
    .Q(\shift_storage.storage [624]));
 sg13g2_dfrbp_1 \shift_storage.storage[625]$_SDFFE_PN0P_  (.CLK(clknet_leaf_18_clk_p2c),
    .RESET_B(net1782),
    .D(_01286_),
    .Q_N(_05515_),
    .Q(\shift_storage.storage [625]));
 sg13g2_dfrbp_1 \shift_storage.storage[626]$_SDFFE_PN0P_  (.CLK(clknet_leaf_18_clk_p2c),
    .RESET_B(net1783),
    .D(_01287_),
    .Q_N(_05514_),
    .Q(\shift_storage.storage [626]));
 sg13g2_dfrbp_1 \shift_storage.storage[627]$_SDFFE_PN0P_  (.CLK(clknet_leaf_17_clk_p2c),
    .RESET_B(net1784),
    .D(_01288_),
    .Q_N(_05513_),
    .Q(\shift_storage.storage [627]));
 sg13g2_dfrbp_1 \shift_storage.storage[628]$_SDFFE_PN0P_  (.CLK(clknet_leaf_17_clk_p2c),
    .RESET_B(net1785),
    .D(_01289_),
    .Q_N(_05512_),
    .Q(\shift_storage.storage [628]));
 sg13g2_dfrbp_1 \shift_storage.storage[629]$_SDFFE_PN0P_  (.CLK(clknet_leaf_18_clk_p2c),
    .RESET_B(net1786),
    .D(_01290_),
    .Q_N(_05511_),
    .Q(\shift_storage.storage [629]));
 sg13g2_dfrbp_1 \shift_storage.storage[62]$_SDFFE_PN0P_  (.CLK(clknet_leaf_17_clk_p2c),
    .RESET_B(net1787),
    .D(_01291_),
    .Q_N(_05510_),
    .Q(\shift_storage.storage [62]));
 sg13g2_dfrbp_1 \shift_storage.storage[630]$_SDFFE_PN0P_  (.CLK(clknet_leaf_18_clk_p2c),
    .RESET_B(net1788),
    .D(_01292_),
    .Q_N(_05509_),
    .Q(\shift_storage.storage [630]));
 sg13g2_dfrbp_1 \shift_storage.storage[631]$_SDFFE_PN0P_  (.CLK(clknet_leaf_6_clk_p2c),
    .RESET_B(net1789),
    .D(_01293_),
    .Q_N(_05508_),
    .Q(\shift_storage.storage [631]));
 sg13g2_dfrbp_1 \shift_storage.storage[632]$_SDFFE_PN0P_  (.CLK(clknet_leaf_5_clk_p2c),
    .RESET_B(net1790),
    .D(_01294_),
    .Q_N(_05507_),
    .Q(\shift_storage.storage [632]));
 sg13g2_dfrbp_1 \shift_storage.storage[633]$_SDFFE_PN0P_  (.CLK(clknet_leaf_5_clk_p2c),
    .RESET_B(net1791),
    .D(_01295_),
    .Q_N(_05506_),
    .Q(\shift_storage.storage [633]));
 sg13g2_dfrbp_1 \shift_storage.storage[634]$_SDFFE_PN0P_  (.CLK(clknet_leaf_6_clk_p2c),
    .RESET_B(net1792),
    .D(_01296_),
    .Q_N(_05505_),
    .Q(\shift_storage.storage [634]));
 sg13g2_dfrbp_1 \shift_storage.storage[635]$_SDFFE_PN0P_  (.CLK(clknet_leaf_6_clk_p2c),
    .RESET_B(net1793),
    .D(_01297_),
    .Q_N(_05504_),
    .Q(\shift_storage.storage [635]));
 sg13g2_dfrbp_1 \shift_storage.storage[636]$_SDFFE_PN0P_  (.CLK(clknet_leaf_6_clk_p2c),
    .RESET_B(net1794),
    .D(_01298_),
    .Q_N(_05503_),
    .Q(\shift_storage.storage [636]));
 sg13g2_dfrbp_1 \shift_storage.storage[637]$_SDFFE_PN0P_  (.CLK(clknet_leaf_5_clk_p2c),
    .RESET_B(net1795),
    .D(_01299_),
    .Q_N(_05502_),
    .Q(\shift_storage.storage [637]));
 sg13g2_dfrbp_1 \shift_storage.storage[638]$_SDFFE_PN0P_  (.CLK(clknet_leaf_5_clk_p2c),
    .RESET_B(net1796),
    .D(_01300_),
    .Q_N(_05501_),
    .Q(\shift_storage.storage [638]));
 sg13g2_dfrbp_1 \shift_storage.storage[639]$_SDFFE_PN0P_  (.CLK(clknet_leaf_5_clk_p2c),
    .RESET_B(net1797),
    .D(_01301_),
    .Q_N(_05500_),
    .Q(\shift_storage.storage [639]));
 sg13g2_dfrbp_1 \shift_storage.storage[63]$_SDFFE_PN0P_  (.CLK(clknet_leaf_5_clk_p2c),
    .RESET_B(net1798),
    .D(_01302_),
    .Q_N(_05499_),
    .Q(\shift_storage.storage [63]));
 sg13g2_dfrbp_1 \shift_storage.storage[640]$_SDFFE_PN0P_  (.CLK(clknet_leaf_4_clk_p2c),
    .RESET_B(net1799),
    .D(_01303_),
    .Q_N(_05498_),
    .Q(\shift_storage.storage [640]));
 sg13g2_dfrbp_1 \shift_storage.storage[641]$_SDFFE_PN0P_  (.CLK(clknet_leaf_4_clk_p2c),
    .RESET_B(net1800),
    .D(_01304_),
    .Q_N(_05497_),
    .Q(\shift_storage.storage [641]));
 sg13g2_dfrbp_1 \shift_storage.storage[642]$_SDFFE_PN0P_  (.CLK(clknet_leaf_4_clk_p2c),
    .RESET_B(net1801),
    .D(_01305_),
    .Q_N(_05496_),
    .Q(\shift_storage.storage [642]));
 sg13g2_dfrbp_1 \shift_storage.storage[643]$_SDFFE_PN0P_  (.CLK(clknet_leaf_3_clk_p2c),
    .RESET_B(net1802),
    .D(_01306_),
    .Q_N(_05495_),
    .Q(\shift_storage.storage [643]));
 sg13g2_dfrbp_1 \shift_storage.storage[644]$_SDFFE_PN0P_  (.CLK(clknet_leaf_3_clk_p2c),
    .RESET_B(net1803),
    .D(_01307_),
    .Q_N(_05494_),
    .Q(\shift_storage.storage [644]));
 sg13g2_dfrbp_1 \shift_storage.storage[645]$_SDFFE_PN0P_  (.CLK(clknet_leaf_3_clk_p2c),
    .RESET_B(net1804),
    .D(_01308_),
    .Q_N(_05493_),
    .Q(\shift_storage.storage [645]));
 sg13g2_dfrbp_1 \shift_storage.storage[646]$_SDFFE_PN0P_  (.CLK(clknet_leaf_3_clk_p2c),
    .RESET_B(net1805),
    .D(_01309_),
    .Q_N(_05492_),
    .Q(\shift_storage.storage [646]));
 sg13g2_dfrbp_1 \shift_storage.storage[647]$_SDFFE_PN0P_  (.CLK(clknet_leaf_1_clk_p2c),
    .RESET_B(net1806),
    .D(_01310_),
    .Q_N(_05491_),
    .Q(\shift_storage.storage [647]));
 sg13g2_dfrbp_1 \shift_storage.storage[648]$_SDFFE_PN0P_  (.CLK(clknet_leaf_3_clk_p2c),
    .RESET_B(net1807),
    .D(_01311_),
    .Q_N(_05490_),
    .Q(\shift_storage.storage [648]));
 sg13g2_dfrbp_1 \shift_storage.storage[649]$_SDFFE_PN0P_  (.CLK(clknet_leaf_4_clk_p2c),
    .RESET_B(net1808),
    .D(_01312_),
    .Q_N(_05489_),
    .Q(\shift_storage.storage [649]));
 sg13g2_dfrbp_1 \shift_storage.storage[64]$_SDFFE_PN0P_  (.CLK(clknet_leaf_1_clk_p2c),
    .RESET_B(net1809),
    .D(_01313_),
    .Q_N(_05488_),
    .Q(\shift_storage.storage [64]));
 sg13g2_dfrbp_1 \shift_storage.storage[650]$_SDFFE_PN0P_  (.CLK(clknet_leaf_0_clk_p2c),
    .RESET_B(net1810),
    .D(_01314_),
    .Q_N(_05487_),
    .Q(\shift_storage.storage [650]));
 sg13g2_dfrbp_1 \shift_storage.storage[651]$_SDFFE_PN0P_  (.CLK(clknet_leaf_0_clk_p2c),
    .RESET_B(net1811),
    .D(_01315_),
    .Q_N(_05486_),
    .Q(\shift_storage.storage [651]));
 sg13g2_dfrbp_1 \shift_storage.storage[652]$_SDFFE_PN0P_  (.CLK(clknet_leaf_0_clk_p2c),
    .RESET_B(net1812),
    .D(_01316_),
    .Q_N(_05485_),
    .Q(\shift_storage.storage [652]));
 sg13g2_dfrbp_1 \shift_storage.storage[653]$_SDFFE_PN0P_  (.CLK(clknet_leaf_0_clk_p2c),
    .RESET_B(net1813),
    .D(_01317_),
    .Q_N(_05484_),
    .Q(\shift_storage.storage [653]));
 sg13g2_dfrbp_1 \shift_storage.storage[654]$_SDFFE_PN0P_  (.CLK(clknet_leaf_1_clk_p2c),
    .RESET_B(net1814),
    .D(_01318_),
    .Q_N(_05483_),
    .Q(\shift_storage.storage [654]));
 sg13g2_dfrbp_1 \shift_storage.storage[655]$_SDFFE_PN0P_  (.CLK(clknet_leaf_294_clk_p2c),
    .RESET_B(net1815),
    .D(_01319_),
    .Q_N(_05482_),
    .Q(\shift_storage.storage [655]));
 sg13g2_dfrbp_1 \shift_storage.storage[656]$_SDFFE_PN0P_  (.CLK(clknet_leaf_294_clk_p2c),
    .RESET_B(net1816),
    .D(_01320_),
    .Q_N(_05481_),
    .Q(\shift_storage.storage [656]));
 sg13g2_dfrbp_1 \shift_storage.storage[657]$_SDFFE_PN0P_  (.CLK(clknet_leaf_0_clk_p2c),
    .RESET_B(net1817),
    .D(_01321_),
    .Q_N(_05480_),
    .Q(\shift_storage.storage [657]));
 sg13g2_dfrbp_1 \shift_storage.storage[658]$_SDFFE_PN0P_  (.CLK(clknet_leaf_293_clk_p2c),
    .RESET_B(net1818),
    .D(_01322_),
    .Q_N(_05479_),
    .Q(\shift_storage.storage [658]));
 sg13g2_dfrbp_1 \shift_storage.storage[659]$_SDFFE_PN0P_  (.CLK(clknet_leaf_293_clk_p2c),
    .RESET_B(net1819),
    .D(_01323_),
    .Q_N(_05478_),
    .Q(\shift_storage.storage [659]));
 sg13g2_dfrbp_1 \shift_storage.storage[65]$_SDFFE_PN0P_  (.CLK(clknet_leaf_1_clk_p2c),
    .RESET_B(net1820),
    .D(_01324_),
    .Q_N(_05477_),
    .Q(\shift_storage.storage [65]));
 sg13g2_dfrbp_1 \shift_storage.storage[660]$_SDFFE_PN0P_  (.CLK(clknet_leaf_293_clk_p2c),
    .RESET_B(net1821),
    .D(_01325_),
    .Q_N(_05476_),
    .Q(\shift_storage.storage [660]));
 sg13g2_dfrbp_1 \shift_storage.storage[661]$_SDFFE_PN0P_  (.CLK(clknet_leaf_293_clk_p2c),
    .RESET_B(net1822),
    .D(_01326_),
    .Q_N(_05475_),
    .Q(\shift_storage.storage [661]));
 sg13g2_dfrbp_1 \shift_storage.storage[662]$_SDFFE_PN0P_  (.CLK(clknet_leaf_293_clk_p2c),
    .RESET_B(net1823),
    .D(_01327_),
    .Q_N(_05474_),
    .Q(\shift_storage.storage [662]));
 sg13g2_dfrbp_1 \shift_storage.storage[663]$_SDFFE_PN0P_  (.CLK(clknet_leaf_293_clk_p2c),
    .RESET_B(net1824),
    .D(_01328_),
    .Q_N(_05473_),
    .Q(\shift_storage.storage [663]));
 sg13g2_dfrbp_1 \shift_storage.storage[664]$_SDFFE_PN0P_  (.CLK(clknet_leaf_292_clk_p2c),
    .RESET_B(net1825),
    .D(_01329_),
    .Q_N(_05472_),
    .Q(\shift_storage.storage [664]));
 sg13g2_dfrbp_1 \shift_storage.storage[665]$_SDFFE_PN0P_  (.CLK(clknet_leaf_292_clk_p2c),
    .RESET_B(net1826),
    .D(_01330_),
    .Q_N(_05471_),
    .Q(\shift_storage.storage [665]));
 sg13g2_dfrbp_1 \shift_storage.storage[666]$_SDFFE_PN0P_  (.CLK(clknet_leaf_292_clk_p2c),
    .RESET_B(net1827),
    .D(_01331_),
    .Q_N(_05470_),
    .Q(\shift_storage.storage [666]));
 sg13g2_dfrbp_1 \shift_storage.storage[667]$_SDFFE_PN0P_  (.CLK(clknet_leaf_294_clk_p2c),
    .RESET_B(net1828),
    .D(_01332_),
    .Q_N(_05469_),
    .Q(\shift_storage.storage [667]));
 sg13g2_dfrbp_1 \shift_storage.storage[668]$_SDFFE_PN0P_  (.CLK(clknet_leaf_290_clk_p2c),
    .RESET_B(net1829),
    .D(_01333_),
    .Q_N(_05468_),
    .Q(\shift_storage.storage [668]));
 sg13g2_dfrbp_1 \shift_storage.storage[669]$_SDFFE_PN0P_  (.CLK(clknet_leaf_291_clk_p2c),
    .RESET_B(net1830),
    .D(_01334_),
    .Q_N(_05467_),
    .Q(\shift_storage.storage [669]));
 sg13g2_dfrbp_1 \shift_storage.storage[66]$_SDFFE_PN0P_  (.CLK(clknet_leaf_1_clk_p2c),
    .RESET_B(net1831),
    .D(_01335_),
    .Q_N(_05466_),
    .Q(\shift_storage.storage [66]));
 sg13g2_dfrbp_1 \shift_storage.storage[670]$_SDFFE_PN0P_  (.CLK(clknet_leaf_292_clk_p2c),
    .RESET_B(net1832),
    .D(_01336_),
    .Q_N(_05465_),
    .Q(\shift_storage.storage [670]));
 sg13g2_dfrbp_1 \shift_storage.storage[671]$_SDFFE_PN0P_  (.CLK(clknet_leaf_292_clk_p2c),
    .RESET_B(net1833),
    .D(_01337_),
    .Q_N(_05464_),
    .Q(\shift_storage.storage [671]));
 sg13g2_dfrbp_1 \shift_storage.storage[672]$_SDFFE_PN0P_  (.CLK(clknet_leaf_292_clk_p2c),
    .RESET_B(net1834),
    .D(_01338_),
    .Q_N(_05463_),
    .Q(\shift_storage.storage [672]));
 sg13g2_dfrbp_1 \shift_storage.storage[673]$_SDFFE_PN0P_  (.CLK(clknet_leaf_291_clk_p2c),
    .RESET_B(net1835),
    .D(_01339_),
    .Q_N(_05462_),
    .Q(\shift_storage.storage [673]));
 sg13g2_dfrbp_1 \shift_storage.storage[674]$_SDFFE_PN0P_  (.CLK(clknet_leaf_291_clk_p2c),
    .RESET_B(net1836),
    .D(_01340_),
    .Q_N(_05461_),
    .Q(\shift_storage.storage [674]));
 sg13g2_dfrbp_1 \shift_storage.storage[675]$_SDFFE_PN0P_  (.CLK(clknet_leaf_288_clk_p2c),
    .RESET_B(net1837),
    .D(_01341_),
    .Q_N(_05460_),
    .Q(\shift_storage.storage [675]));
 sg13g2_dfrbp_1 \shift_storage.storage[676]$_SDFFE_PN0P_  (.CLK(clknet_leaf_291_clk_p2c),
    .RESET_B(net1838),
    .D(_01342_),
    .Q_N(_05459_),
    .Q(\shift_storage.storage [676]));
 sg13g2_dfrbp_1 \shift_storage.storage[677]$_SDFFE_PN0P_  (.CLK(clknet_leaf_289_clk_p2c),
    .RESET_B(net1839),
    .D(_01343_),
    .Q_N(_05458_),
    .Q(\shift_storage.storage [677]));
 sg13g2_dfrbp_1 \shift_storage.storage[678]$_SDFFE_PN0P_  (.CLK(clknet_leaf_291_clk_p2c),
    .RESET_B(net1840),
    .D(_01344_),
    .Q_N(_05457_),
    .Q(\shift_storage.storage [678]));
 sg13g2_dfrbp_1 \shift_storage.storage[679]$_SDFFE_PN0P_  (.CLK(clknet_leaf_290_clk_p2c),
    .RESET_B(net1841),
    .D(_01345_),
    .Q_N(_05456_),
    .Q(\shift_storage.storage [679]));
 sg13g2_dfrbp_1 \shift_storage.storage[67]$_SDFFE_PN0P_  (.CLK(clknet_leaf_1_clk_p2c),
    .RESET_B(net1842),
    .D(_01346_),
    .Q_N(_05455_),
    .Q(\shift_storage.storage [67]));
 sg13g2_dfrbp_1 \shift_storage.storage[680]$_SDFFE_PN0P_  (.CLK(clknet_leaf_290_clk_p2c),
    .RESET_B(net1843),
    .D(_01347_),
    .Q_N(_05454_),
    .Q(\shift_storage.storage [680]));
 sg13g2_dfrbp_1 \shift_storage.storage[681]$_SDFFE_PN0P_  (.CLK(clknet_leaf_290_clk_p2c),
    .RESET_B(net1844),
    .D(_01348_),
    .Q_N(_05453_),
    .Q(\shift_storage.storage [681]));
 sg13g2_dfrbp_1 \shift_storage.storage[682]$_SDFFE_PN0P_  (.CLK(clknet_leaf_2_clk_p2c),
    .RESET_B(net1845),
    .D(_01349_),
    .Q_N(_05452_),
    .Q(\shift_storage.storage [682]));
 sg13g2_dfrbp_1 \shift_storage.storage[683]$_SDFFE_PN0P_  (.CLK(clknet_leaf_2_clk_p2c),
    .RESET_B(net1846),
    .D(_01350_),
    .Q_N(_05451_),
    .Q(\shift_storage.storage [683]));
 sg13g2_dfrbp_1 \shift_storage.storage[684]$_SDFFE_PN0P_  (.CLK(clknet_leaf_2_clk_p2c),
    .RESET_B(net1847),
    .D(_01351_),
    .Q_N(_05450_),
    .Q(\shift_storage.storage [684]));
 sg13g2_dfrbp_1 \shift_storage.storage[685]$_SDFFE_PN0P_  (.CLK(clknet_leaf_2_clk_p2c),
    .RESET_B(net1848),
    .D(_01352_),
    .Q_N(_05449_),
    .Q(\shift_storage.storage [685]));
 sg13g2_dfrbp_1 \shift_storage.storage[686]$_SDFFE_PN0P_  (.CLK(clknet_leaf_2_clk_p2c),
    .RESET_B(net1849),
    .D(_01353_),
    .Q_N(_05448_),
    .Q(\shift_storage.storage [686]));
 sg13g2_dfrbp_1 \shift_storage.storage[687]$_SDFFE_PN0P_  (.CLK(clknet_leaf_2_clk_p2c),
    .RESET_B(net1850),
    .D(_01354_),
    .Q_N(_05447_),
    .Q(\shift_storage.storage [687]));
 sg13g2_dfrbp_1 \shift_storage.storage[688]$_SDFFE_PN0P_  (.CLK(clknet_leaf_8_clk_p2c),
    .RESET_B(net1851),
    .D(_01355_),
    .Q_N(_05446_),
    .Q(\shift_storage.storage [688]));
 sg13g2_dfrbp_1 \shift_storage.storage[689]$_SDFFE_PN0P_  (.CLK(clknet_leaf_9_clk_p2c),
    .RESET_B(net1852),
    .D(_01356_),
    .Q_N(_05445_),
    .Q(\shift_storage.storage [689]));
 sg13g2_dfrbp_1 \shift_storage.storage[68]$_SDFFE_PN0P_  (.CLK(clknet_leaf_8_clk_p2c),
    .RESET_B(net1853),
    .D(_01357_),
    .Q_N(_05444_),
    .Q(\shift_storage.storage [68]));
 sg13g2_dfrbp_1 \shift_storage.storage[690]$_SDFFE_PN0P_  (.CLK(clknet_leaf_8_clk_p2c),
    .RESET_B(net1854),
    .D(_01358_),
    .Q_N(_05443_),
    .Q(\shift_storage.storage [690]));
 sg13g2_dfrbp_1 \shift_storage.storage[691]$_SDFFE_PN0P_  (.CLK(clknet_leaf_8_clk_p2c),
    .RESET_B(net1855),
    .D(_01359_),
    .Q_N(_05442_),
    .Q(\shift_storage.storage [691]));
 sg13g2_dfrbp_1 \shift_storage.storage[692]$_SDFFE_PN0P_  (.CLK(clknet_leaf_8_clk_p2c),
    .RESET_B(net1856),
    .D(_01360_),
    .Q_N(_05441_),
    .Q(\shift_storage.storage [692]));
 sg13g2_dfrbp_1 \shift_storage.storage[693]$_SDFFE_PN0P_  (.CLK(clknet_leaf_7_clk_p2c),
    .RESET_B(net1857),
    .D(_01361_),
    .Q_N(_05440_),
    .Q(\shift_storage.storage [693]));
 sg13g2_dfrbp_1 \shift_storage.storage[694]$_SDFFE_PN0P_  (.CLK(clknet_leaf_7_clk_p2c),
    .RESET_B(net1858),
    .D(_01362_),
    .Q_N(_05439_),
    .Q(\shift_storage.storage [694]));
 sg13g2_dfrbp_1 \shift_storage.storage[695]$_SDFFE_PN0P_  (.CLK(clknet_leaf_7_clk_p2c),
    .RESET_B(net1859),
    .D(_01363_),
    .Q_N(_05438_),
    .Q(\shift_storage.storage [695]));
 sg13g2_dfrbp_1 \shift_storage.storage[696]$_SDFFE_PN0P_  (.CLK(clknet_leaf_9_clk_p2c),
    .RESET_B(net1860),
    .D(_01364_),
    .Q_N(_05437_),
    .Q(\shift_storage.storage [696]));
 sg13g2_dfrbp_1 \shift_storage.storage[697]$_SDFFE_PN0P_  (.CLK(clknet_leaf_9_clk_p2c),
    .RESET_B(net1861),
    .D(_01365_),
    .Q_N(_05436_),
    .Q(\shift_storage.storage [697]));
 sg13g2_dfrbp_1 \shift_storage.storage[698]$_SDFFE_PN0P_  (.CLK(clknet_leaf_9_clk_p2c),
    .RESET_B(net1862),
    .D(_01366_),
    .Q_N(_05435_),
    .Q(\shift_storage.storage [698]));
 sg13g2_dfrbp_1 \shift_storage.storage[699]$_SDFFE_PN0P_  (.CLK(clknet_leaf_10_clk_p2c),
    .RESET_B(net1863),
    .D(_01367_),
    .Q_N(_05434_),
    .Q(\shift_storage.storage [699]));
 sg13g2_dfrbp_1 \shift_storage.storage[69]$_SDFFE_PN0P_  (.CLK(clknet_leaf_9_clk_p2c),
    .RESET_B(net1864),
    .D(_01368_),
    .Q_N(_05433_),
    .Q(\shift_storage.storage [69]));
 sg13g2_dfrbp_1 \shift_storage.storage[6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_11_clk_p2c),
    .RESET_B(net1865),
    .D(_01369_),
    .Q_N(_05432_),
    .Q(\shift_storage.storage [6]));
 sg13g2_dfrbp_1 \shift_storage.storage[700]$_SDFFE_PN0P_  (.CLK(clknet_leaf_10_clk_p2c),
    .RESET_B(net1866),
    .D(_01370_),
    .Q_N(_05431_),
    .Q(\shift_storage.storage [700]));
 sg13g2_dfrbp_1 \shift_storage.storage[701]$_SDFFE_PN0P_  (.CLK(clknet_leaf_281_clk_p2c),
    .RESET_B(net1867),
    .D(_01371_),
    .Q_N(_05430_),
    .Q(\shift_storage.storage [701]));
 sg13g2_dfrbp_1 \shift_storage.storage[702]$_SDFFE_PN0P_  (.CLK(clknet_leaf_11_clk_p2c),
    .RESET_B(net1868),
    .D(_01372_),
    .Q_N(_05429_),
    .Q(\shift_storage.storage [702]));
 sg13g2_dfrbp_1 \shift_storage.storage[703]$_SDFFE_PN0P_  (.CLK(clknet_leaf_281_clk_p2c),
    .RESET_B(net1869),
    .D(_01373_),
    .Q_N(_05428_),
    .Q(\shift_storage.storage [703]));
 sg13g2_dfrbp_1 \shift_storage.storage[704]$_SDFFE_PN0P_  (.CLK(clknet_leaf_283_clk_p2c),
    .RESET_B(net1870),
    .D(_01374_),
    .Q_N(_05427_),
    .Q(\shift_storage.storage [704]));
 sg13g2_dfrbp_1 \shift_storage.storage[705]$_SDFFE_PN0P_  (.CLK(clknet_leaf_283_clk_p2c),
    .RESET_B(net1871),
    .D(_01375_),
    .Q_N(_05426_),
    .Q(\shift_storage.storage [705]));
 sg13g2_dfrbp_1 \shift_storage.storage[706]$_SDFFE_PN0P_  (.CLK(clknet_leaf_9_clk_p2c),
    .RESET_B(net1872),
    .D(_01376_),
    .Q_N(_05425_),
    .Q(\shift_storage.storage [706]));
 sg13g2_dfrbp_1 \shift_storage.storage[707]$_SDFFE_PN0P_  (.CLK(clknet_leaf_9_clk_p2c),
    .RESET_B(net1873),
    .D(_01377_),
    .Q_N(_05424_),
    .Q(\shift_storage.storage [707]));
 sg13g2_dfrbp_1 \shift_storage.storage[708]$_SDFFE_PN0P_  (.CLK(clknet_leaf_283_clk_p2c),
    .RESET_B(net1874),
    .D(_01378_),
    .Q_N(_05423_),
    .Q(\shift_storage.storage [708]));
 sg13g2_dfrbp_1 \shift_storage.storage[709]$_SDFFE_PN0P_  (.CLK(clknet_leaf_283_clk_p2c),
    .RESET_B(net1875),
    .D(_01379_),
    .Q_N(_05422_),
    .Q(\shift_storage.storage [709]));
 sg13g2_dfrbp_1 \shift_storage.storage[70]$_SDFFE_PN0P_  (.CLK(clknet_leaf_284_clk_p2c),
    .RESET_B(net1876),
    .D(_01380_),
    .Q_N(_05421_),
    .Q(\shift_storage.storage [70]));
 sg13g2_dfrbp_1 \shift_storage.storage[710]$_SDFFE_PN0P_  (.CLK(clknet_leaf_283_clk_p2c),
    .RESET_B(net1877),
    .D(_01381_),
    .Q_N(_05420_),
    .Q(\shift_storage.storage [710]));
 sg13g2_dfrbp_1 \shift_storage.storage[711]$_SDFFE_PN0P_  (.CLK(clknet_leaf_283_clk_p2c),
    .RESET_B(net1878),
    .D(_01382_),
    .Q_N(_05419_),
    .Q(\shift_storage.storage [711]));
 sg13g2_dfrbp_1 \shift_storage.storage[712]$_SDFFE_PN0P_  (.CLK(clknet_leaf_284_clk_p2c),
    .RESET_B(net1879),
    .D(_01383_),
    .Q_N(_05418_),
    .Q(\shift_storage.storage [712]));
 sg13g2_dfrbp_1 \shift_storage.storage[713]$_SDFFE_PN0P_  (.CLK(clknet_leaf_284_clk_p2c),
    .RESET_B(net1880),
    .D(_01384_),
    .Q_N(_05417_),
    .Q(\shift_storage.storage [713]));
 sg13g2_dfrbp_1 \shift_storage.storage[714]$_SDFFE_PN0P_  (.CLK(clknet_leaf_284_clk_p2c),
    .RESET_B(net1881),
    .D(_01385_),
    .Q_N(_05416_),
    .Q(\shift_storage.storage [714]));
 sg13g2_dfrbp_1 \shift_storage.storage[715]$_SDFFE_PN0P_  (.CLK(clknet_leaf_284_clk_p2c),
    .RESET_B(net1882),
    .D(_01386_),
    .Q_N(_05415_),
    .Q(\shift_storage.storage [715]));
 sg13g2_dfrbp_1 \shift_storage.storage[716]$_SDFFE_PN0P_  (.CLK(clknet_leaf_290_clk_p2c),
    .RESET_B(net1883),
    .D(_01387_),
    .Q_N(_05414_),
    .Q(\shift_storage.storage [716]));
 sg13g2_dfrbp_1 \shift_storage.storage[717]$_SDFFE_PN0P_  (.CLK(clknet_leaf_289_clk_p2c),
    .RESET_B(net1884),
    .D(_01388_),
    .Q_N(_05413_),
    .Q(\shift_storage.storage [717]));
 sg13g2_dfrbp_1 \shift_storage.storage[718]$_SDFFE_PN0P_  (.CLK(clknet_leaf_289_clk_p2c),
    .RESET_B(net1885),
    .D(_01389_),
    .Q_N(_05412_),
    .Q(\shift_storage.storage [718]));
 sg13g2_dfrbp_1 \shift_storage.storage[719]$_SDFFE_PN0P_  (.CLK(clknet_leaf_289_clk_p2c),
    .RESET_B(net1886),
    .D(_01390_),
    .Q_N(_05411_),
    .Q(\shift_storage.storage [719]));
 sg13g2_dfrbp_1 \shift_storage.storage[71]$_SDFFE_PN0P_  (.CLK(clknet_leaf_284_clk_p2c),
    .RESET_B(net1887),
    .D(_01391_),
    .Q_N(_05410_),
    .Q(\shift_storage.storage [71]));
 sg13g2_dfrbp_1 \shift_storage.storage[720]$_SDFFE_PN0P_  (.CLK(clknet_leaf_289_clk_p2c),
    .RESET_B(net1888),
    .D(_01392_),
    .Q_N(_05409_),
    .Q(\shift_storage.storage [720]));
 sg13g2_dfrbp_1 \shift_storage.storage[721]$_SDFFE_PN0P_  (.CLK(clknet_leaf_289_clk_p2c),
    .RESET_B(net1889),
    .D(_01393_),
    .Q_N(_05408_),
    .Q(\shift_storage.storage [721]));
 sg13g2_dfrbp_1 \shift_storage.storage[722]$_SDFFE_PN0P_  (.CLK(clknet_leaf_288_clk_p2c),
    .RESET_B(net1890),
    .D(_01394_),
    .Q_N(_05407_),
    .Q(\shift_storage.storage [722]));
 sg13g2_dfrbp_1 \shift_storage.storage[723]$_SDFFE_PN0P_  (.CLK(clknet_leaf_288_clk_p2c),
    .RESET_B(net1891),
    .D(_01395_),
    .Q_N(_05406_),
    .Q(\shift_storage.storage [723]));
 sg13g2_dfrbp_1 \shift_storage.storage[724]$_SDFFE_PN0P_  (.CLK(clknet_leaf_288_clk_p2c),
    .RESET_B(net1892),
    .D(_01396_),
    .Q_N(_05405_),
    .Q(\shift_storage.storage [724]));
 sg13g2_dfrbp_1 \shift_storage.storage[725]$_SDFFE_PN0P_  (.CLK(clknet_leaf_288_clk_p2c),
    .RESET_B(net1893),
    .D(_01397_),
    .Q_N(_05404_),
    .Q(\shift_storage.storage [725]));
 sg13g2_dfrbp_1 \shift_storage.storage[726]$_SDFFE_PN0P_  (.CLK(clknet_leaf_287_clk_p2c),
    .RESET_B(net1894),
    .D(_01398_),
    .Q_N(_05403_),
    .Q(\shift_storage.storage [726]));
 sg13g2_dfrbp_1 \shift_storage.storage[727]$_SDFFE_PN0P_  (.CLK(clknet_leaf_287_clk_p2c),
    .RESET_B(net1895),
    .D(_01399_),
    .Q_N(_05402_),
    .Q(\shift_storage.storage [727]));
 sg13g2_dfrbp_1 \shift_storage.storage[728]$_SDFFE_PN0P_  (.CLK(clknet_leaf_287_clk_p2c),
    .RESET_B(net1896),
    .D(_01400_),
    .Q_N(_05401_),
    .Q(\shift_storage.storage [728]));
 sg13g2_dfrbp_1 \shift_storage.storage[729]$_SDFFE_PN0P_  (.CLK(clknet_leaf_287_clk_p2c),
    .RESET_B(net1897),
    .D(_01401_),
    .Q_N(_05400_),
    .Q(\shift_storage.storage [729]));
 sg13g2_dfrbp_1 \shift_storage.storage[72]$_SDFFE_PN0P_  (.CLK(clknet_leaf_286_clk_p2c),
    .RESET_B(net1898),
    .D(_01402_),
    .Q_N(_05399_),
    .Q(\shift_storage.storage [72]));
 sg13g2_dfrbp_1 \shift_storage.storage[730]$_SDFFE_PN0P_  (.CLK(clknet_leaf_287_clk_p2c),
    .RESET_B(net1899),
    .D(_01403_),
    .Q_N(_05398_),
    .Q(\shift_storage.storage [730]));
 sg13g2_dfrbp_1 \shift_storage.storage[731]$_SDFFE_PN0P_  (.CLK(clknet_leaf_285_clk_p2c),
    .RESET_B(net1900),
    .D(_01404_),
    .Q_N(_05397_),
    .Q(\shift_storage.storage [731]));
 sg13g2_dfrbp_1 \shift_storage.storage[732]$_SDFFE_PN0P_  (.CLK(clknet_leaf_286_clk_p2c),
    .RESET_B(net1901),
    .D(_01405_),
    .Q_N(_05396_),
    .Q(\shift_storage.storage [732]));
 sg13g2_dfrbp_1 \shift_storage.storage[733]$_SDFFE_PN0P_  (.CLK(clknet_leaf_285_clk_p2c),
    .RESET_B(net1902),
    .D(_01406_),
    .Q_N(_05395_),
    .Q(\shift_storage.storage [733]));
 sg13g2_dfrbp_1 \shift_storage.storage[734]$_SDFFE_PN0P_  (.CLK(clknet_leaf_285_clk_p2c),
    .RESET_B(net1903),
    .D(_01407_),
    .Q_N(_05394_),
    .Q(\shift_storage.storage [734]));
 sg13g2_dfrbp_1 \shift_storage.storage[735]$_SDFFE_PN0P_  (.CLK(clknet_leaf_276_clk_p2c),
    .RESET_B(net1904),
    .D(_01408_),
    .Q_N(_05393_),
    .Q(\shift_storage.storage [735]));
 sg13g2_dfrbp_1 \shift_storage.storage[736]$_SDFFE_PN0P_  (.CLK(clknet_leaf_275_clk_p2c),
    .RESET_B(net1905),
    .D(_01409_),
    .Q_N(_05392_),
    .Q(\shift_storage.storage [736]));
 sg13g2_dfrbp_1 \shift_storage.storage[737]$_SDFFE_PN0P_  (.CLK(clknet_leaf_274_clk_p2c),
    .RESET_B(net1906),
    .D(_01410_),
    .Q_N(_05391_),
    .Q(\shift_storage.storage [737]));
 sg13g2_dfrbp_1 \shift_storage.storage[738]$_SDFFE_PN0P_  (.CLK(clknet_leaf_286_clk_p2c),
    .RESET_B(net1907),
    .D(_01411_),
    .Q_N(_05390_),
    .Q(\shift_storage.storage [738]));
 sg13g2_dfrbp_1 \shift_storage.storage[739]$_SDFFE_PN0P_  (.CLK(clknet_leaf_286_clk_p2c),
    .RESET_B(net1908),
    .D(_01412_),
    .Q_N(_05389_),
    .Q(\shift_storage.storage [739]));
 sg13g2_dfrbp_1 \shift_storage.storage[73]$_SDFFE_PN0P_  (.CLK(clknet_leaf_274_clk_p2c),
    .RESET_B(net1909),
    .D(_01413_),
    .Q_N(_05388_),
    .Q(\shift_storage.storage [73]));
 sg13g2_dfrbp_1 \shift_storage.storage[740]$_SDFFE_PN0P_  (.CLK(clknet_leaf_286_clk_p2c),
    .RESET_B(net1910),
    .D(_01414_),
    .Q_N(_05387_),
    .Q(\shift_storage.storage [740]));
 sg13g2_dfrbp_1 \shift_storage.storage[741]$_SDFFE_PN0P_  (.CLK(clknet_leaf_286_clk_p2c),
    .RESET_B(net1911),
    .D(_01415_),
    .Q_N(_05386_),
    .Q(\shift_storage.storage [741]));
 sg13g2_dfrbp_1 \shift_storage.storage[742]$_SDFFE_PN0P_  (.CLK(clknet_leaf_287_clk_p2c),
    .RESET_B(net1912),
    .D(_01416_),
    .Q_N(_05385_),
    .Q(\shift_storage.storage [742]));
 sg13g2_dfrbp_1 \shift_storage.storage[743]$_SDFFE_PN0P_  (.CLK(clknet_leaf_274_clk_p2c),
    .RESET_B(net1913),
    .D(_01417_),
    .Q_N(_05384_),
    .Q(\shift_storage.storage [743]));
 sg13g2_dfrbp_1 \shift_storage.storage[744]$_SDFFE_PN0P_  (.CLK(clknet_leaf_274_clk_p2c),
    .RESET_B(net1914),
    .D(_01418_),
    .Q_N(_05383_),
    .Q(\shift_storage.storage [744]));
 sg13g2_dfrbp_1 \shift_storage.storage[745]$_SDFFE_PN0P_  (.CLK(clknet_leaf_274_clk_p2c),
    .RESET_B(net1915),
    .D(_01419_),
    .Q_N(_05382_),
    .Q(\shift_storage.storage [745]));
 sg13g2_dfrbp_1 \shift_storage.storage[746]$_SDFFE_PN0P_  (.CLK(clknet_leaf_274_clk_p2c),
    .RESET_B(net1916),
    .D(_01420_),
    .Q_N(_05381_),
    .Q(\shift_storage.storage [746]));
 sg13g2_dfrbp_1 \shift_storage.storage[747]$_SDFFE_PN0P_  (.CLK(clknet_leaf_273_clk_p2c),
    .RESET_B(net1917),
    .D(_01421_),
    .Q_N(_05380_),
    .Q(\shift_storage.storage [747]));
 sg13g2_dfrbp_1 \shift_storage.storage[748]$_SDFFE_PN0P_  (.CLK(clknet_leaf_273_clk_p2c),
    .RESET_B(net1918),
    .D(_01422_),
    .Q_N(_05379_),
    .Q(\shift_storage.storage [748]));
 sg13g2_dfrbp_1 \shift_storage.storage[749]$_SDFFE_PN0P_  (.CLK(clknet_leaf_273_clk_p2c),
    .RESET_B(net1919),
    .D(_01423_),
    .Q_N(_05378_),
    .Q(\shift_storage.storage [749]));
 sg13g2_dfrbp_1 \shift_storage.storage[74]$_SDFFE_PN0P_  (.CLK(clknet_leaf_275_clk_p2c),
    .RESET_B(net1920),
    .D(_01424_),
    .Q_N(_05377_),
    .Q(\shift_storage.storage [74]));
 sg13g2_dfrbp_1 \shift_storage.storage[750]$_SDFFE_PN0P_  (.CLK(clknet_leaf_272_clk_p2c),
    .RESET_B(net1921),
    .D(_01425_),
    .Q_N(_05376_),
    .Q(\shift_storage.storage [750]));
 sg13g2_dfrbp_1 \shift_storage.storage[751]$_SDFFE_PN0P_  (.CLK(clknet_leaf_273_clk_p2c),
    .RESET_B(net1922),
    .D(_01426_),
    .Q_N(_05375_),
    .Q(\shift_storage.storage [751]));
 sg13g2_dfrbp_1 \shift_storage.storage[752]$_SDFFE_PN0P_  (.CLK(clknet_leaf_269_clk_p2c),
    .RESET_B(net1923),
    .D(_01427_),
    .Q_N(_05374_),
    .Q(\shift_storage.storage [752]));
 sg13g2_dfrbp_1 \shift_storage.storage[753]$_SDFFE_PN0P_  (.CLK(clknet_leaf_272_clk_p2c),
    .RESET_B(net1924),
    .D(_01428_),
    .Q_N(_05373_),
    .Q(\shift_storage.storage [753]));
 sg13g2_dfrbp_1 \shift_storage.storage[754]$_SDFFE_PN0P_  (.CLK(clknet_leaf_269_clk_p2c),
    .RESET_B(net1925),
    .D(_01429_),
    .Q_N(_05372_),
    .Q(\shift_storage.storage [754]));
 sg13g2_dfrbp_1 \shift_storage.storage[755]$_SDFFE_PN0P_  (.CLK(clknet_leaf_269_clk_p2c),
    .RESET_B(net1926),
    .D(_01430_),
    .Q_N(_05371_),
    .Q(\shift_storage.storage [755]));
 sg13g2_dfrbp_1 \shift_storage.storage[756]$_SDFFE_PN0P_  (.CLK(clknet_leaf_272_clk_p2c),
    .RESET_B(net1927),
    .D(_01431_),
    .Q_N(_05370_),
    .Q(\shift_storage.storage [756]));
 sg13g2_dfrbp_1 \shift_storage.storage[757]$_SDFFE_PN0P_  (.CLK(clknet_leaf_272_clk_p2c),
    .RESET_B(net1928),
    .D(_01432_),
    .Q_N(_05369_),
    .Q(\shift_storage.storage [757]));
 sg13g2_dfrbp_1 \shift_storage.storage[758]$_SDFFE_PN0P_  (.CLK(clknet_leaf_273_clk_p2c),
    .RESET_B(net1929),
    .D(_01433_),
    .Q_N(_05368_),
    .Q(\shift_storage.storage [758]));
 sg13g2_dfrbp_1 \shift_storage.storage[759]$_SDFFE_PN0P_  (.CLK(clknet_leaf_273_clk_p2c),
    .RESET_B(net1930),
    .D(_01434_),
    .Q_N(_05367_),
    .Q(\shift_storage.storage [759]));
 sg13g2_dfrbp_1 \shift_storage.storage[75]$_SDFFE_PN0P_  (.CLK(clknet_leaf_275_clk_p2c),
    .RESET_B(net1931),
    .D(_01435_),
    .Q_N(_05366_),
    .Q(\shift_storage.storage [75]));
 sg13g2_dfrbp_1 \shift_storage.storage[760]$_SDFFE_PN0P_  (.CLK(clknet_leaf_275_clk_p2c),
    .RESET_B(net1932),
    .D(_01436_),
    .Q_N(_05365_),
    .Q(\shift_storage.storage [760]));
 sg13g2_dfrbp_1 \shift_storage.storage[761]$_SDFFE_PN0P_  (.CLK(clknet_leaf_275_clk_p2c),
    .RESET_B(net1933),
    .D(_01437_),
    .Q_N(_05364_),
    .Q(\shift_storage.storage [761]));
 sg13g2_dfrbp_1 \shift_storage.storage[762]$_SDFFE_PN0P_  (.CLK(clknet_leaf_272_clk_p2c),
    .RESET_B(net1934),
    .D(_01438_),
    .Q_N(_05363_),
    .Q(\shift_storage.storage [762]));
 sg13g2_dfrbp_1 \shift_storage.storage[763]$_SDFFE_PN0P_  (.CLK(clknet_leaf_271_clk_p2c),
    .RESET_B(net1935),
    .D(_01439_),
    .Q_N(_05362_),
    .Q(\shift_storage.storage [763]));
 sg13g2_dfrbp_1 \shift_storage.storage[764]$_SDFFE_PN0P_  (.CLK(clknet_leaf_271_clk_p2c),
    .RESET_B(net1936),
    .D(_01440_),
    .Q_N(_05361_),
    .Q(\shift_storage.storage [764]));
 sg13g2_dfrbp_1 \shift_storage.storage[765]$_SDFFE_PN0P_  (.CLK(clknet_leaf_277_clk_p2c),
    .RESET_B(net1937),
    .D(_01441_),
    .Q_N(_05360_),
    .Q(\shift_storage.storage [765]));
 sg13g2_dfrbp_1 \shift_storage.storage[766]$_SDFFE_PN0P_  (.CLK(clknet_leaf_277_clk_p2c),
    .RESET_B(net1938),
    .D(_01442_),
    .Q_N(_05359_),
    .Q(\shift_storage.storage [766]));
 sg13g2_dfrbp_1 \shift_storage.storage[767]$_SDFFE_PN0P_  (.CLK(clknet_leaf_277_clk_p2c),
    .RESET_B(net1939),
    .D(_01443_),
    .Q_N(_05358_),
    .Q(\shift_storage.storage [767]));
 sg13g2_dfrbp_1 \shift_storage.storage[768]$_SDFFE_PN0P_  (.CLK(clknet_leaf_277_clk_p2c),
    .RESET_B(net1940),
    .D(_01444_),
    .Q_N(_05357_),
    .Q(\shift_storage.storage [768]));
 sg13g2_dfrbp_1 \shift_storage.storage[769]$_SDFFE_PN0P_  (.CLK(clknet_leaf_278_clk_p2c),
    .RESET_B(net1941),
    .D(_01445_),
    .Q_N(_05356_),
    .Q(\shift_storage.storage [769]));
 sg13g2_dfrbp_1 \shift_storage.storage[76]$_SDFFE_PN0P_  (.CLK(clknet_leaf_277_clk_p2c),
    .RESET_B(net1942),
    .D(_01446_),
    .Q_N(_05355_),
    .Q(\shift_storage.storage [76]));
 sg13g2_dfrbp_1 \shift_storage.storage[770]$_SDFFE_PN0P_  (.CLK(clknet_leaf_276_clk_p2c),
    .RESET_B(net1943),
    .D(_01447_),
    .Q_N(_05354_),
    .Q(\shift_storage.storage [770]));
 sg13g2_dfrbp_1 \shift_storage.storage[771]$_SDFFE_PN0P_  (.CLK(clknet_leaf_276_clk_p2c),
    .RESET_B(net1944),
    .D(_01448_),
    .Q_N(_05353_),
    .Q(\shift_storage.storage [771]));
 sg13g2_dfrbp_1 \shift_storage.storage[772]$_SDFFE_PN0P_  (.CLK(clknet_leaf_276_clk_p2c),
    .RESET_B(net1945),
    .D(_01449_),
    .Q_N(_05352_),
    .Q(\shift_storage.storage [772]));
 sg13g2_dfrbp_1 \shift_storage.storage[773]$_SDFFE_PN0P_  (.CLK(clknet_leaf_276_clk_p2c),
    .RESET_B(net1946),
    .D(_01450_),
    .Q_N(_05351_),
    .Q(\shift_storage.storage [773]));
 sg13g2_dfrbp_1 \shift_storage.storage[774]$_SDFFE_PN0P_  (.CLK(clknet_leaf_285_clk_p2c),
    .RESET_B(net1947),
    .D(_01451_),
    .Q_N(_05350_),
    .Q(\shift_storage.storage [774]));
 sg13g2_dfrbp_1 \shift_storage.storage[775]$_SDFFE_PN0P_  (.CLK(clknet_leaf_276_clk_p2c),
    .RESET_B(net1948),
    .D(_01452_),
    .Q_N(_05349_),
    .Q(\shift_storage.storage [775]));
 sg13g2_dfrbp_1 \shift_storage.storage[776]$_SDFFE_PN0P_  (.CLK(clknet_leaf_285_clk_p2c),
    .RESET_B(net1949),
    .D(_01453_),
    .Q_N(_05348_),
    .Q(\shift_storage.storage [776]));
 sg13g2_dfrbp_1 \shift_storage.storage[777]$_SDFFE_PN0P_  (.CLK(clknet_leaf_285_clk_p2c),
    .RESET_B(net1950),
    .D(_01454_),
    .Q_N(_05347_),
    .Q(\shift_storage.storage [777]));
 sg13g2_dfrbp_1 \shift_storage.storage[778]$_SDFFE_PN0P_  (.CLK(clknet_leaf_282_clk_p2c),
    .RESET_B(net1951),
    .D(_01455_),
    .Q_N(_05346_),
    .Q(\shift_storage.storage [778]));
 sg13g2_dfrbp_1 \shift_storage.storage[779]$_SDFFE_PN0P_  (.CLK(clknet_leaf_282_clk_p2c),
    .RESET_B(net1952),
    .D(_01456_),
    .Q_N(_05345_),
    .Q(\shift_storage.storage [779]));
 sg13g2_dfrbp_1 \shift_storage.storage[77]$_SDFFE_PN0P_  (.CLK(clknet_leaf_279_clk_p2c),
    .RESET_B(net1953),
    .D(_01457_),
    .Q_N(_05344_),
    .Q(\shift_storage.storage [77]));
 sg13g2_dfrbp_1 \shift_storage.storage[780]$_SDFFE_PN0P_  (.CLK(clknet_leaf_282_clk_p2c),
    .RESET_B(net1954),
    .D(_01458_),
    .Q_N(_05343_),
    .Q(\shift_storage.storage [780]));
 sg13g2_dfrbp_1 \shift_storage.storage[781]$_SDFFE_PN0P_  (.CLK(clknet_leaf_282_clk_p2c),
    .RESET_B(net1955),
    .D(_01459_),
    .Q_N(_05342_),
    .Q(\shift_storage.storage [781]));
 sg13g2_dfrbp_1 \shift_storage.storage[782]$_SDFFE_PN0P_  (.CLK(clknet_leaf_282_clk_p2c),
    .RESET_B(net1956),
    .D(_01460_),
    .Q_N(_05341_),
    .Q(\shift_storage.storage [782]));
 sg13g2_dfrbp_1 \shift_storage.storage[783]$_SDFFE_PN0P_  (.CLK(clknet_leaf_279_clk_p2c),
    .RESET_B(net1957),
    .D(_01461_),
    .Q_N(_05340_),
    .Q(\shift_storage.storage [783]));
 sg13g2_dfrbp_1 \shift_storage.storage[784]$_SDFFE_PN0P_  (.CLK(clknet_leaf_279_clk_p2c),
    .RESET_B(net1958),
    .D(_01462_),
    .Q_N(_05339_),
    .Q(\shift_storage.storage [784]));
 sg13g2_dfrbp_1 \shift_storage.storage[785]$_SDFFE_PN0P_  (.CLK(clknet_leaf_279_clk_p2c),
    .RESET_B(net1959),
    .D(_01463_),
    .Q_N(_05338_),
    .Q(\shift_storage.storage [785]));
 sg13g2_dfrbp_1 \shift_storage.storage[786]$_SDFFE_PN0P_  (.CLK(clknet_leaf_280_clk_p2c),
    .RESET_B(net1960),
    .D(_01464_),
    .Q_N(_05337_),
    .Q(\shift_storage.storage [786]));
 sg13g2_dfrbp_1 \shift_storage.storage[787]$_SDFFE_PN0P_  (.CLK(clknet_leaf_281_clk_p2c),
    .RESET_B(net1961),
    .D(_01465_),
    .Q_N(_05336_),
    .Q(\shift_storage.storage [787]));
 sg13g2_dfrbp_1 \shift_storage.storage[788]$_SDFFE_PN0P_  (.CLK(clknet_leaf_281_clk_p2c),
    .RESET_B(net1962),
    .D(_01466_),
    .Q_N(_05335_),
    .Q(\shift_storage.storage [788]));
 sg13g2_dfrbp_1 \shift_storage.storage[789]$_SDFFE_PN0P_  (.CLK(clknet_leaf_281_clk_p2c),
    .RESET_B(net1963),
    .D(_01467_),
    .Q_N(_05334_),
    .Q(\shift_storage.storage [789]));
 sg13g2_dfrbp_1 \shift_storage.storage[78]$_SDFFE_PN0P_  (.CLK(clknet_leaf_280_clk_p2c),
    .RESET_B(net1964),
    .D(_01468_),
    .Q_N(_05333_),
    .Q(\shift_storage.storage [78]));
 sg13g2_dfrbp_1 \shift_storage.storage[790]$_SDFFE_PN0P_  (.CLK(clknet_leaf_281_clk_p2c),
    .RESET_B(net1965),
    .D(_01469_),
    .Q_N(_05332_),
    .Q(\shift_storage.storage [790]));
 sg13g2_dfrbp_1 \shift_storage.storage[791]$_SDFFE_PN0P_  (.CLK(clknet_leaf_281_clk_p2c),
    .RESET_B(net1966),
    .D(_01470_),
    .Q_N(_05331_),
    .Q(\shift_storage.storage [791]));
 sg13g2_dfrbp_1 \shift_storage.storage[792]$_SDFFE_PN0P_  (.CLK(clknet_leaf_280_clk_p2c),
    .RESET_B(net1967),
    .D(_01471_),
    .Q_N(_05330_),
    .Q(\shift_storage.storage [792]));
 sg13g2_dfrbp_1 \shift_storage.storage[793]$_SDFFE_PN0P_  (.CLK(clknet_leaf_280_clk_p2c),
    .RESET_B(net1968),
    .D(_01472_),
    .Q_N(_05329_),
    .Q(\shift_storage.storage [793]));
 sg13g2_dfrbp_1 \shift_storage.storage[794]$_SDFFE_PN0P_  (.CLK(clknet_leaf_11_clk_p2c),
    .RESET_B(net1969),
    .D(_01473_),
    .Q_N(_05328_),
    .Q(\shift_storage.storage [794]));
 sg13g2_dfrbp_1 \shift_storage.storage[795]$_SDFFE_PN0P_  (.CLK(clknet_leaf_11_clk_p2c),
    .RESET_B(net1970),
    .D(_01474_),
    .Q_N(_05327_),
    .Q(\shift_storage.storage [795]));
 sg13g2_dfrbp_1 \shift_storage.storage[796]$_SDFFE_PN0P_  (.CLK(clknet_leaf_11_clk_p2c),
    .RESET_B(net1971),
    .D(_01475_),
    .Q_N(_05326_),
    .Q(\shift_storage.storage [796]));
 sg13g2_dfrbp_1 \shift_storage.storage[797]$_SDFFE_PN0P_  (.CLK(clknet_leaf_11_clk_p2c),
    .RESET_B(net1972),
    .D(_01476_),
    .Q_N(_05325_),
    .Q(\shift_storage.storage [797]));
 sg13g2_dfrbp_1 \shift_storage.storage[798]$_SDFFE_PN0P_  (.CLK(clknet_leaf_257_clk_p2c),
    .RESET_B(net1973),
    .D(_01477_),
    .Q_N(_05324_),
    .Q(\shift_storage.storage [798]));
 sg13g2_dfrbp_1 \shift_storage.storage[799]$_SDFFE_PN0P_  (.CLK(clknet_leaf_257_clk_p2c),
    .RESET_B(net1974),
    .D(_01478_),
    .Q_N(_05323_),
    .Q(\shift_storage.storage [799]));
 sg13g2_dfrbp_1 \shift_storage.storage[79]$_SDFFE_PN0P_  (.CLK(clknet_leaf_258_clk_p2c),
    .RESET_B(net1975),
    .D(_01479_),
    .Q_N(_05322_),
    .Q(\shift_storage.storage [79]));
 sg13g2_dfrbp_1 \shift_storage.storage[7]$_SDFFE_PN0P_  (.CLK(clknet_leaf_257_clk_p2c),
    .RESET_B(net1976),
    .D(_01480_),
    .Q_N(_05321_),
    .Q(\shift_storage.storage [7]));
 sg13g2_dfrbp_1 \shift_storage.storage[800]$_SDFFE_PN0P_  (.CLK(clknet_leaf_257_clk_p2c),
    .RESET_B(net1977),
    .D(_01481_),
    .Q_N(_05320_),
    .Q(\shift_storage.storage [800]));
 sg13g2_dfrbp_1 \shift_storage.storage[801]$_SDFFE_PN0P_  (.CLK(clknet_leaf_258_clk_p2c),
    .RESET_B(net1978),
    .D(_01482_),
    .Q_N(_05319_),
    .Q(\shift_storage.storage [801]));
 sg13g2_dfrbp_1 \shift_storage.storage[802]$_SDFFE_PN0P_  (.CLK(clknet_leaf_258_clk_p2c),
    .RESET_B(net1979),
    .D(_01483_),
    .Q_N(_05318_),
    .Q(\shift_storage.storage [802]));
 sg13g2_dfrbp_1 \shift_storage.storage[803]$_SDFFE_PN0P_  (.CLK(clknet_leaf_257_clk_p2c),
    .RESET_B(net1980),
    .D(_01484_),
    .Q_N(_05317_),
    .Q(\shift_storage.storage [803]));
 sg13g2_dfrbp_1 \shift_storage.storage[804]$_SDFFE_PN0P_  (.CLK(clknet_leaf_258_clk_p2c),
    .RESET_B(net1981),
    .D(_01485_),
    .Q_N(_05316_),
    .Q(\shift_storage.storage [804]));
 sg13g2_dfrbp_1 \shift_storage.storage[805]$_SDFFE_PN0P_  (.CLK(clknet_leaf_258_clk_p2c),
    .RESET_B(net1982),
    .D(_01486_),
    .Q_N(_05315_),
    .Q(\shift_storage.storage [805]));
 sg13g2_dfrbp_1 \shift_storage.storage[806]$_SDFFE_PN0P_  (.CLK(clknet_leaf_259_clk_p2c),
    .RESET_B(net1983),
    .D(_01487_),
    .Q_N(_05314_),
    .Q(\shift_storage.storage [806]));
 sg13g2_dfrbp_1 \shift_storage.storage[807]$_SDFFE_PN0P_  (.CLK(clknet_leaf_259_clk_p2c),
    .RESET_B(net1984),
    .D(_01488_),
    .Q_N(_05313_),
    .Q(\shift_storage.storage [807]));
 sg13g2_dfrbp_1 \shift_storage.storage[808]$_SDFFE_PN0P_  (.CLK(clknet_leaf_260_clk_p2c),
    .RESET_B(net1985),
    .D(_01489_),
    .Q_N(_05312_),
    .Q(\shift_storage.storage [808]));
 sg13g2_dfrbp_1 \shift_storage.storage[809]$_SDFFE_PN0P_  (.CLK(clknet_leaf_260_clk_p2c),
    .RESET_B(net1986),
    .D(_01490_),
    .Q_N(_05311_),
    .Q(\shift_storage.storage [809]));
 sg13g2_dfrbp_1 \shift_storage.storage[80]$_SDFFE_PN0P_  (.CLK(clknet_leaf_260_clk_p2c),
    .RESET_B(net1987),
    .D(_01491_),
    .Q_N(_05310_),
    .Q(\shift_storage.storage [80]));
 sg13g2_dfrbp_1 \shift_storage.storage[810]$_SDFFE_PN0P_  (.CLK(clknet_leaf_280_clk_p2c),
    .RESET_B(net1988),
    .D(_01492_),
    .Q_N(_05309_),
    .Q(\shift_storage.storage [810]));
 sg13g2_dfrbp_1 \shift_storage.storage[811]$_SDFFE_PN0P_  (.CLK(clknet_leaf_279_clk_p2c),
    .RESET_B(net1989),
    .D(_01493_),
    .Q_N(_05308_),
    .Q(\shift_storage.storage [811]));
 sg13g2_dfrbp_1 \shift_storage.storage[812]$_SDFFE_PN0P_  (.CLK(clknet_leaf_279_clk_p2c),
    .RESET_B(net1990),
    .D(_01494_),
    .Q_N(_05307_),
    .Q(\shift_storage.storage [812]));
 sg13g2_dfrbp_1 \shift_storage.storage[813]$_SDFFE_PN0P_  (.CLK(clknet_leaf_278_clk_p2c),
    .RESET_B(net1991),
    .D(_01495_),
    .Q_N(_05306_),
    .Q(\shift_storage.storage [813]));
 sg13g2_dfrbp_1 \shift_storage.storage[814]$_SDFFE_PN0P_  (.CLK(clknet_leaf_278_clk_p2c),
    .RESET_B(net1992),
    .D(_01496_),
    .Q_N(_05305_),
    .Q(\shift_storage.storage [814]));
 sg13g2_dfrbp_1 \shift_storage.storage[815]$_SDFFE_PN0P_  (.CLK(clknet_leaf_260_clk_p2c),
    .RESET_B(net1993),
    .D(_01497_),
    .Q_N(_05304_),
    .Q(\shift_storage.storage [815]));
 sg13g2_dfrbp_1 \shift_storage.storage[816]$_SDFFE_PN0P_  (.CLK(clknet_leaf_260_clk_p2c),
    .RESET_B(net1994),
    .D(_01498_),
    .Q_N(_05303_),
    .Q(\shift_storage.storage [816]));
 sg13g2_dfrbp_1 \shift_storage.storage[817]$_SDFFE_PN0P_  (.CLK(clknet_leaf_260_clk_p2c),
    .RESET_B(net1995),
    .D(_01499_),
    .Q_N(_05302_),
    .Q(\shift_storage.storage [817]));
 sg13g2_dfrbp_1 \shift_storage.storage[818]$_SDFFE_PN0P_  (.CLK(clknet_leaf_261_clk_p2c),
    .RESET_B(net1996),
    .D(_01500_),
    .Q_N(_05301_),
    .Q(\shift_storage.storage [818]));
 sg13g2_dfrbp_1 \shift_storage.storage[819]$_SDFFE_PN0P_  (.CLK(clknet_leaf_266_clk_p2c),
    .RESET_B(net1997),
    .D(_01501_),
    .Q_N(_05300_),
    .Q(\shift_storage.storage [819]));
 sg13g2_dfrbp_1 \shift_storage.storage[81]$_SDFFE_PN0P_  (.CLK(clknet_leaf_266_clk_p2c),
    .RESET_B(net1998),
    .D(_01502_),
    .Q_N(_05299_),
    .Q(\shift_storage.storage [81]));
 sg13g2_dfrbp_1 \shift_storage.storage[820]$_SDFFE_PN0P_  (.CLK(clknet_leaf_271_clk_p2c),
    .RESET_B(net1999),
    .D(_01503_),
    .Q_N(_05298_),
    .Q(\shift_storage.storage [820]));
 sg13g2_dfrbp_1 \shift_storage.storage[821]$_SDFFE_PN0P_  (.CLK(clknet_leaf_271_clk_p2c),
    .RESET_B(net2000),
    .D(_01504_),
    .Q_N(_05297_),
    .Q(\shift_storage.storage [821]));
 sg13g2_dfrbp_1 \shift_storage.storage[822]$_SDFFE_PN0P_  (.CLK(clknet_leaf_278_clk_p2c),
    .RESET_B(net2001),
    .D(_01505_),
    .Q_N(_05296_),
    .Q(\shift_storage.storage [822]));
 sg13g2_dfrbp_1 \shift_storage.storage[823]$_SDFFE_PN0P_  (.CLK(clknet_leaf_278_clk_p2c),
    .RESET_B(net2002),
    .D(_01506_),
    .Q_N(_05295_),
    .Q(\shift_storage.storage [823]));
 sg13g2_dfrbp_1 \shift_storage.storage[824]$_SDFFE_PN0P_  (.CLK(clknet_leaf_271_clk_p2c),
    .RESET_B(net2003),
    .D(_01507_),
    .Q_N(_05294_),
    .Q(\shift_storage.storage [824]));
 sg13g2_dfrbp_1 \shift_storage.storage[825]$_SDFFE_PN0P_  (.CLK(clknet_leaf_270_clk_p2c),
    .RESET_B(net2004),
    .D(_01508_),
    .Q_N(_05293_),
    .Q(\shift_storage.storage [825]));
 sg13g2_dfrbp_1 \shift_storage.storage[826]$_SDFFE_PN0P_  (.CLK(clknet_leaf_270_clk_p2c),
    .RESET_B(net2005),
    .D(_01509_),
    .Q_N(_05292_),
    .Q(\shift_storage.storage [826]));
 sg13g2_dfrbp_1 \shift_storage.storage[827]$_SDFFE_PN0P_  (.CLK(clknet_leaf_270_clk_p2c),
    .RESET_B(net2006),
    .D(_01510_),
    .Q_N(_05291_),
    .Q(\shift_storage.storage [827]));
 sg13g2_dfrbp_1 \shift_storage.storage[828]$_SDFFE_PN0P_  (.CLK(clknet_leaf_270_clk_p2c),
    .RESET_B(net2007),
    .D(_01511_),
    .Q_N(_05290_),
    .Q(\shift_storage.storage [828]));
 sg13g2_dfrbp_1 \shift_storage.storage[829]$_SDFFE_PN0P_  (.CLK(clknet_leaf_270_clk_p2c),
    .RESET_B(net2008),
    .D(_01512_),
    .Q_N(_05289_),
    .Q(\shift_storage.storage [829]));
 sg13g2_dfrbp_1 \shift_storage.storage[82]$_SDFFE_PN0P_  (.CLK(clknet_leaf_266_clk_p2c),
    .RESET_B(net2009),
    .D(_01513_),
    .Q_N(_05288_),
    .Q(\shift_storage.storage [82]));
 sg13g2_dfrbp_1 \shift_storage.storage[830]$_SDFFE_PN0P_  (.CLK(clknet_leaf_270_clk_p2c),
    .RESET_B(net2010),
    .D(_01514_),
    .Q_N(_05287_),
    .Q(\shift_storage.storage [830]));
 sg13g2_dfrbp_1 \shift_storage.storage[831]$_SDFFE_PN0P_  (.CLK(clknet_leaf_270_clk_p2c),
    .RESET_B(net2011),
    .D(_01515_),
    .Q_N(_05286_),
    .Q(\shift_storage.storage [831]));
 sg13g2_dfrbp_1 \shift_storage.storage[832]$_SDFFE_PN0P_  (.CLK(clknet_leaf_266_clk_p2c),
    .RESET_B(net2012),
    .D(_01516_),
    .Q_N(_05285_),
    .Q(\shift_storage.storage [832]));
 sg13g2_dfrbp_1 \shift_storage.storage[833]$_SDFFE_PN0P_  (.CLK(clknet_leaf_266_clk_p2c),
    .RESET_B(net2013),
    .D(_01517_),
    .Q_N(_05284_),
    .Q(\shift_storage.storage [833]));
 sg13g2_dfrbp_1 \shift_storage.storage[834]$_SDFFE_PN0P_  (.CLK(clknet_leaf_266_clk_p2c),
    .RESET_B(net2014),
    .D(_01518_),
    .Q_N(_05283_),
    .Q(\shift_storage.storage [834]));
 sg13g2_dfrbp_1 \shift_storage.storage[835]$_SDFFE_PN0P_  (.CLK(clknet_leaf_267_clk_p2c),
    .RESET_B(net2015),
    .D(_01519_),
    .Q_N(_05282_),
    .Q(\shift_storage.storage [835]));
 sg13g2_dfrbp_1 \shift_storage.storage[836]$_SDFFE_PN0P_  (.CLK(clknet_leaf_267_clk_p2c),
    .RESET_B(net2016),
    .D(_01520_),
    .Q_N(_05281_),
    .Q(\shift_storage.storage [836]));
 sg13g2_dfrbp_1 \shift_storage.storage[837]$_SDFFE_PN0P_  (.CLK(clknet_leaf_267_clk_p2c),
    .RESET_B(net2017),
    .D(_01521_),
    .Q_N(_05280_),
    .Q(\shift_storage.storage [837]));
 sg13g2_dfrbp_1 \shift_storage.storage[838]$_SDFFE_PN0P_  (.CLK(clknet_leaf_268_clk_p2c),
    .RESET_B(net2018),
    .D(_01522_),
    .Q_N(_05279_),
    .Q(\shift_storage.storage [838]));
 sg13g2_dfrbp_1 \shift_storage.storage[839]$_SDFFE_PN0P_  (.CLK(clknet_leaf_268_clk_p2c),
    .RESET_B(net2019),
    .D(_01523_),
    .Q_N(_05278_),
    .Q(\shift_storage.storage [839]));
 sg13g2_dfrbp_1 \shift_storage.storage[83]$_SDFFE_PN0P_  (.CLK(clknet_leaf_267_clk_p2c),
    .RESET_B(net2020),
    .D(_01524_),
    .Q_N(_05277_),
    .Q(\shift_storage.storage [83]));
 sg13g2_dfrbp_1 \shift_storage.storage[840]$_SDFFE_PN0P_  (.CLK(clknet_leaf_268_clk_p2c),
    .RESET_B(net2021),
    .D(_01525_),
    .Q_N(_05276_),
    .Q(\shift_storage.storage [840]));
 sg13g2_dfrbp_1 \shift_storage.storage[841]$_SDFFE_PN0P_  (.CLK(clknet_leaf_269_clk_p2c),
    .RESET_B(net2022),
    .D(_01526_),
    .Q_N(_05275_),
    .Q(\shift_storage.storage [841]));
 sg13g2_dfrbp_1 \shift_storage.storage[842]$_SDFFE_PN0P_  (.CLK(clknet_leaf_269_clk_p2c),
    .RESET_B(net2023),
    .D(_01527_),
    .Q_N(_05274_),
    .Q(\shift_storage.storage [842]));
 sg13g2_dfrbp_1 \shift_storage.storage[843]$_SDFFE_PN0P_  (.CLK(clknet_leaf_268_clk_p2c),
    .RESET_B(net2024),
    .D(_01528_),
    .Q_N(_05273_),
    .Q(\shift_storage.storage [843]));
 sg13g2_dfrbp_1 \shift_storage.storage[844]$_SDFFE_PN0P_  (.CLK(clknet_leaf_268_clk_p2c),
    .RESET_B(net2025),
    .D(_01529_),
    .Q_N(_05272_),
    .Q(\shift_storage.storage [844]));
 sg13g2_dfrbp_1 \shift_storage.storage[845]$_SDFFE_PN0P_  (.CLK(clknet_leaf_224_clk_p2c),
    .RESET_B(net2026),
    .D(_01530_),
    .Q_N(_05271_),
    .Q(\shift_storage.storage [845]));
 sg13g2_dfrbp_1 \shift_storage.storage[846]$_SDFFE_PN0P_  (.CLK(clknet_leaf_224_clk_p2c),
    .RESET_B(net2027),
    .D(_01531_),
    .Q_N(_05270_),
    .Q(\shift_storage.storage [846]));
 sg13g2_dfrbp_1 \shift_storage.storage[847]$_SDFFE_PN0P_  (.CLK(clknet_leaf_268_clk_p2c),
    .RESET_B(net2028),
    .D(_01532_),
    .Q_N(_05269_),
    .Q(\shift_storage.storage [847]));
 sg13g2_dfrbp_1 \shift_storage.storage[848]$_SDFFE_PN0P_  (.CLK(clknet_leaf_267_clk_p2c),
    .RESET_B(net2029),
    .D(_01533_),
    .Q_N(_05268_),
    .Q(\shift_storage.storage [848]));
 sg13g2_dfrbp_1 \shift_storage.storage[849]$_SDFFE_PN0P_  (.CLK(clknet_leaf_267_clk_p2c),
    .RESET_B(net2030),
    .D(_01534_),
    .Q_N(_05267_),
    .Q(\shift_storage.storage [849]));
 sg13g2_dfrbp_1 \shift_storage.storage[84]$_SDFFE_PN0P_  (.CLK(clknet_leaf_265_clk_p2c),
    .RESET_B(net2031),
    .D(_01535_),
    .Q_N(_05266_),
    .Q(\shift_storage.storage [84]));
 sg13g2_dfrbp_1 \shift_storage.storage[850]$_SDFFE_PN0P_  (.CLK(clknet_leaf_224_clk_p2c),
    .RESET_B(net2032),
    .D(_01536_),
    .Q_N(_05265_),
    .Q(\shift_storage.storage [850]));
 sg13g2_dfrbp_1 \shift_storage.storage[851]$_SDFFE_PN0P_  (.CLK(clknet_leaf_224_clk_p2c),
    .RESET_B(net2033),
    .D(_01537_),
    .Q_N(_05264_),
    .Q(\shift_storage.storage [851]));
 sg13g2_dfrbp_1 \shift_storage.storage[852]$_SDFFE_PN0P_  (.CLK(clknet_leaf_225_clk_p2c),
    .RESET_B(net2034),
    .D(_01538_),
    .Q_N(_05263_),
    .Q(\shift_storage.storage [852]));
 sg13g2_dfrbp_1 \shift_storage.storage[853]$_SDFFE_PN0P_  (.CLK(clknet_leaf_225_clk_p2c),
    .RESET_B(net2035),
    .D(_01539_),
    .Q_N(_05262_),
    .Q(\shift_storage.storage [853]));
 sg13g2_dfrbp_1 \shift_storage.storage[854]$_SDFFE_PN0P_  (.CLK(clknet_leaf_225_clk_p2c),
    .RESET_B(net2036),
    .D(_01540_),
    .Q_N(_05261_),
    .Q(\shift_storage.storage [854]));
 sg13g2_dfrbp_1 \shift_storage.storage[855]$_SDFFE_PN0P_  (.CLK(clknet_leaf_225_clk_p2c),
    .RESET_B(net2037),
    .D(_01541_),
    .Q_N(_05260_),
    .Q(\shift_storage.storage [855]));
 sg13g2_dfrbp_1 \shift_storage.storage[856]$_SDFFE_PN0P_  (.CLK(clknet_leaf_225_clk_p2c),
    .RESET_B(net2038),
    .D(_01542_),
    .Q_N(_05259_),
    .Q(\shift_storage.storage [856]));
 sg13g2_dfrbp_1 \shift_storage.storage[857]$_SDFFE_PN0P_  (.CLK(clknet_leaf_226_clk_p2c),
    .RESET_B(net2039),
    .D(_01543_),
    .Q_N(_05258_),
    .Q(\shift_storage.storage [857]));
 sg13g2_dfrbp_1 \shift_storage.storage[858]$_SDFFE_PN0P_  (.CLK(clknet_leaf_226_clk_p2c),
    .RESET_B(net2040),
    .D(_01544_),
    .Q_N(_05257_),
    .Q(\shift_storage.storage [858]));
 sg13g2_dfrbp_1 \shift_storage.storage[859]$_SDFFE_PN0P_  (.CLK(clknet_leaf_226_clk_p2c),
    .RESET_B(net2041),
    .D(_01545_),
    .Q_N(_05256_),
    .Q(\shift_storage.storage [859]));
 sg13g2_dfrbp_1 \shift_storage.storage[85]$_SDFFE_PN0P_  (.CLK(clknet_leaf_226_clk_p2c),
    .RESET_B(net2042),
    .D(_01546_),
    .Q_N(_05255_),
    .Q(\shift_storage.storage [85]));
 sg13g2_dfrbp_1 \shift_storage.storage[860]$_SDFFE_PN0P_  (.CLK(clknet_leaf_227_clk_p2c),
    .RESET_B(net2043),
    .D(_01547_),
    .Q_N(_05254_),
    .Q(\shift_storage.storage [860]));
 sg13g2_dfrbp_1 \shift_storage.storage[861]$_SDFFE_PN0P_  (.CLK(clknet_leaf_226_clk_p2c),
    .RESET_B(net2044),
    .D(_01548_),
    .Q_N(_05253_),
    .Q(\shift_storage.storage [861]));
 sg13g2_dfrbp_1 \shift_storage.storage[862]$_SDFFE_PN0P_  (.CLK(clknet_leaf_226_clk_p2c),
    .RESET_B(net2045),
    .D(_01549_),
    .Q_N(_05252_),
    .Q(\shift_storage.storage [862]));
 sg13g2_dfrbp_1 \shift_storage.storage[863]$_SDFFE_PN0P_  (.CLK(clknet_leaf_227_clk_p2c),
    .RESET_B(net2046),
    .D(_01550_),
    .Q_N(_05251_),
    .Q(\shift_storage.storage [863]));
 sg13g2_dfrbp_1 \shift_storage.storage[864]$_SDFFE_PN0P_  (.CLK(clknet_leaf_227_clk_p2c),
    .RESET_B(net2047),
    .D(_01551_),
    .Q_N(_05250_),
    .Q(\shift_storage.storage [864]));
 sg13g2_dfrbp_1 \shift_storage.storage[865]$_SDFFE_PN0P_  (.CLK(clknet_leaf_228_clk_p2c),
    .RESET_B(net2048),
    .D(_01552_),
    .Q_N(_05249_),
    .Q(\shift_storage.storage [865]));
 sg13g2_dfrbp_1 \shift_storage.storage[866]$_SDFFE_PN0P_  (.CLK(clknet_leaf_227_clk_p2c),
    .RESET_B(net2049),
    .D(_01553_),
    .Q_N(_05248_),
    .Q(\shift_storage.storage [866]));
 sg13g2_dfrbp_1 \shift_storage.storage[867]$_SDFFE_PN0P_  (.CLK(clknet_leaf_228_clk_p2c),
    .RESET_B(net2050),
    .D(_01554_),
    .Q_N(_05247_),
    .Q(\shift_storage.storage [867]));
 sg13g2_dfrbp_1 \shift_storage.storage[868]$_SDFFE_PN0P_  (.CLK(clknet_leaf_228_clk_p2c),
    .RESET_B(net2051),
    .D(_01555_),
    .Q_N(_05246_),
    .Q(\shift_storage.storage [868]));
 sg13g2_dfrbp_1 \shift_storage.storage[869]$_SDFFE_PN0P_  (.CLK(clknet_leaf_227_clk_p2c),
    .RESET_B(net2052),
    .D(_01556_),
    .Q_N(_05245_),
    .Q(\shift_storage.storage [869]));
 sg13g2_dfrbp_1 \shift_storage.storage[86]$_SDFFE_PN0P_  (.CLK(clknet_leaf_264_clk_p2c),
    .RESET_B(net2053),
    .D(_01557_),
    .Q_N(_05244_),
    .Q(\shift_storage.storage [86]));
 sg13g2_dfrbp_1 \shift_storage.storage[870]$_SDFFE_PN0P_  (.CLK(clknet_leaf_228_clk_p2c),
    .RESET_B(net2054),
    .D(_01558_),
    .Q_N(_05243_),
    .Q(\shift_storage.storage [870]));
 sg13g2_dfrbp_1 \shift_storage.storage[871]$_SDFFE_PN0P_  (.CLK(clknet_leaf_263_clk_p2c),
    .RESET_B(net2055),
    .D(_01559_),
    .Q_N(_05242_),
    .Q(\shift_storage.storage [871]));
 sg13g2_dfrbp_1 \shift_storage.storage[872]$_SDFFE_PN0P_  (.CLK(clknet_leaf_263_clk_p2c),
    .RESET_B(net2056),
    .D(_01560_),
    .Q_N(_05241_),
    .Q(\shift_storage.storage [872]));
 sg13g2_dfrbp_1 \shift_storage.storage[873]$_SDFFE_PN0P_  (.CLK(clknet_leaf_263_clk_p2c),
    .RESET_B(net2057),
    .D(_01561_),
    .Q_N(_05240_),
    .Q(\shift_storage.storage [873]));
 sg13g2_dfrbp_1 \shift_storage.storage[874]$_SDFFE_PN0P_  (.CLK(clknet_leaf_264_clk_p2c),
    .RESET_B(net2058),
    .D(_01562_),
    .Q_N(_05239_),
    .Q(\shift_storage.storage [874]));
 sg13g2_dfrbp_1 \shift_storage.storage[875]$_SDFFE_PN0P_  (.CLK(clknet_leaf_264_clk_p2c),
    .RESET_B(net2059),
    .D(_01563_),
    .Q_N(_05238_),
    .Q(\shift_storage.storage [875]));
 sg13g2_dfrbp_1 \shift_storage.storage[876]$_SDFFE_PN0P_  (.CLK(clknet_leaf_264_clk_p2c),
    .RESET_B(net2060),
    .D(_01564_),
    .Q_N(_05237_),
    .Q(\shift_storage.storage [876]));
 sg13g2_dfrbp_1 \shift_storage.storage[877]$_SDFFE_PN0P_  (.CLK(clknet_leaf_264_clk_p2c),
    .RESET_B(net2061),
    .D(_01565_),
    .Q_N(_05236_),
    .Q(\shift_storage.storage [877]));
 sg13g2_dfrbp_1 \shift_storage.storage[878]$_SDFFE_PN0P_  (.CLK(clknet_leaf_265_clk_p2c),
    .RESET_B(net2062),
    .D(_01566_),
    .Q_N(_05235_),
    .Q(\shift_storage.storage [878]));
 sg13g2_dfrbp_1 \shift_storage.storage[879]$_SDFFE_PN0P_  (.CLK(clknet_leaf_265_clk_p2c),
    .RESET_B(net2063),
    .D(_01567_),
    .Q_N(_05234_),
    .Q(\shift_storage.storage [879]));
 sg13g2_dfrbp_1 \shift_storage.storage[87]$_SDFFE_PN0P_  (.CLK(clknet_leaf_264_clk_p2c),
    .RESET_B(net2064),
    .D(_01568_),
    .Q_N(_05233_),
    .Q(\shift_storage.storage [87]));
 sg13g2_dfrbp_1 \shift_storage.storage[880]$_SDFFE_PN0P_  (.CLK(clknet_leaf_265_clk_p2c),
    .RESET_B(net2065),
    .D(_01569_),
    .Q_N(_05232_),
    .Q(\shift_storage.storage [880]));
 sg13g2_dfrbp_1 \shift_storage.storage[881]$_SDFFE_PN0P_  (.CLK(clknet_leaf_265_clk_p2c),
    .RESET_B(net2066),
    .D(_01570_),
    .Q_N(_05231_),
    .Q(\shift_storage.storage [881]));
 sg13g2_dfrbp_1 \shift_storage.storage[882]$_SDFFE_PN0P_  (.CLK(clknet_leaf_265_clk_p2c),
    .RESET_B(net2067),
    .D(_01571_),
    .Q_N(_05230_),
    .Q(\shift_storage.storage [882]));
 sg13g2_dfrbp_1 \shift_storage.storage[883]$_SDFFE_PN0P_  (.CLK(clknet_leaf_265_clk_p2c),
    .RESET_B(net2068),
    .D(_01572_),
    .Q_N(_05229_),
    .Q(\shift_storage.storage [883]));
 sg13g2_dfrbp_1 \shift_storage.storage[884]$_SDFFE_PN0P_  (.CLK(clknet_leaf_261_clk_p2c),
    .RESET_B(net2069),
    .D(_01573_),
    .Q_N(_05228_),
    .Q(\shift_storage.storage [884]));
 sg13g2_dfrbp_1 \shift_storage.storage[885]$_SDFFE_PN0P_  (.CLK(clknet_leaf_261_clk_p2c),
    .RESET_B(net2070),
    .D(_01574_),
    .Q_N(_05227_),
    .Q(\shift_storage.storage [885]));
 sg13g2_dfrbp_1 \shift_storage.storage[886]$_SDFFE_PN0P_  (.CLK(clknet_leaf_261_clk_p2c),
    .RESET_B(net2071),
    .D(_01575_),
    .Q_N(_05226_),
    .Q(\shift_storage.storage [886]));
 sg13g2_dfrbp_1 \shift_storage.storage[887]$_SDFFE_PN0P_  (.CLK(clknet_leaf_261_clk_p2c),
    .RESET_B(net2072),
    .D(_01576_),
    .Q_N(_05225_),
    .Q(\shift_storage.storage [887]));
 sg13g2_dfrbp_1 \shift_storage.storage[888]$_SDFFE_PN0P_  (.CLK(clknet_leaf_261_clk_p2c),
    .RESET_B(net2073),
    .D(_01577_),
    .Q_N(_05224_),
    .Q(\shift_storage.storage [888]));
 sg13g2_dfrbp_1 \shift_storage.storage[889]$_SDFFE_PN0P_  (.CLK(clknet_leaf_263_clk_p2c),
    .RESET_B(net2074),
    .D(_01578_),
    .Q_N(_05223_),
    .Q(\shift_storage.storage [889]));
 sg13g2_dfrbp_1 \shift_storage.storage[88]$_SDFFE_PN0P_  (.CLK(clknet_leaf_252_clk_p2c),
    .RESET_B(net2075),
    .D(_01579_),
    .Q_N(_05222_),
    .Q(\shift_storage.storage [88]));
 sg13g2_dfrbp_1 \shift_storage.storage[890]$_SDFFE_PN0P_  (.CLK(clknet_leaf_262_clk_p2c),
    .RESET_B(net2076),
    .D(_01580_),
    .Q_N(_05221_),
    .Q(\shift_storage.storage [890]));
 sg13g2_dfrbp_1 \shift_storage.storage[891]$_SDFFE_PN0P_  (.CLK(clknet_leaf_263_clk_p2c),
    .RESET_B(net2077),
    .D(_01581_),
    .Q_N(_05220_),
    .Q(\shift_storage.storage [891]));
 sg13g2_dfrbp_1 \shift_storage.storage[892]$_SDFFE_PN0P_  (.CLK(clknet_leaf_252_clk_p2c),
    .RESET_B(net2078),
    .D(_01582_),
    .Q_N(_05219_),
    .Q(\shift_storage.storage [892]));
 sg13g2_dfrbp_1 \shift_storage.storage[893]$_SDFFE_PN0P_  (.CLK(clknet_leaf_262_clk_p2c),
    .RESET_B(net2079),
    .D(_01583_),
    .Q_N(_05218_),
    .Q(\shift_storage.storage [893]));
 sg13g2_dfrbp_1 \shift_storage.storage[894]$_SDFFE_PN0P_  (.CLK(clknet_leaf_262_clk_p2c),
    .RESET_B(net2080),
    .D(_01584_),
    .Q_N(_05217_),
    .Q(\shift_storage.storage [894]));
 sg13g2_dfrbp_1 \shift_storage.storage[895]$_SDFFE_PN0P_  (.CLK(clknet_leaf_262_clk_p2c),
    .RESET_B(net2081),
    .D(_01585_),
    .Q_N(_05216_),
    .Q(\shift_storage.storage [895]));
 sg13g2_dfrbp_1 \shift_storage.storage[896]$_SDFFE_PN0P_  (.CLK(clknet_leaf_262_clk_p2c),
    .RESET_B(net2082),
    .D(_01586_),
    .Q_N(_05215_),
    .Q(\shift_storage.storage [896]));
 sg13g2_dfrbp_1 \shift_storage.storage[897]$_SDFFE_PN0P_  (.CLK(clknet_leaf_259_clk_p2c),
    .RESET_B(net2083),
    .D(_01587_),
    .Q_N(_05214_),
    .Q(\shift_storage.storage [897]));
 sg13g2_dfrbp_1 \shift_storage.storage[898]$_SDFFE_PN0P_  (.CLK(clknet_leaf_262_clk_p2c),
    .RESET_B(net2084),
    .D(_01588_),
    .Q_N(_05213_),
    .Q(\shift_storage.storage [898]));
 sg13g2_dfrbp_1 \shift_storage.storage[899]$_SDFFE_PN0P_  (.CLK(clknet_leaf_259_clk_p2c),
    .RESET_B(net2085),
    .D(_01589_),
    .Q_N(_05212_),
    .Q(\shift_storage.storage [899]));
 sg13g2_dfrbp_1 \shift_storage.storage[89]$_SDFFE_PN0P_  (.CLK(clknet_leaf_252_clk_p2c),
    .RESET_B(net2086),
    .D(_01590_),
    .Q_N(_05211_),
    .Q(\shift_storage.storage [89]));
 sg13g2_dfrbp_1 \shift_storage.storage[8]$_SDFFE_PN0P_  (.CLK(clknet_leaf_252_clk_p2c),
    .RESET_B(net2087),
    .D(_01591_),
    .Q_N(_05210_),
    .Q(\shift_storage.storage [8]));
 sg13g2_dfrbp_1 \shift_storage.storage[900]$_SDFFE_PN0P_  (.CLK(clknet_leaf_252_clk_p2c),
    .RESET_B(net2088),
    .D(_01592_),
    .Q_N(_05209_),
    .Q(\shift_storage.storage [900]));
 sg13g2_dfrbp_1 \shift_storage.storage[901]$_SDFFE_PN0P_  (.CLK(clknet_leaf_255_clk_p2c),
    .RESET_B(net2089),
    .D(_01593_),
    .Q_N(_05208_),
    .Q(\shift_storage.storage [901]));
 sg13g2_dfrbp_1 \shift_storage.storage[902]$_SDFFE_PN0P_  (.CLK(clknet_leaf_259_clk_p2c),
    .RESET_B(net2090),
    .D(_01594_),
    .Q_N(_05207_),
    .Q(\shift_storage.storage [902]));
 sg13g2_dfrbp_1 \shift_storage.storage[903]$_SDFFE_PN0P_  (.CLK(clknet_leaf_256_clk_p2c),
    .RESET_B(net2091),
    .D(_01595_),
    .Q_N(_05206_),
    .Q(\shift_storage.storage [903]));
 sg13g2_dfrbp_1 \shift_storage.storage[904]$_SDFFE_PN0P_  (.CLK(clknet_leaf_256_clk_p2c),
    .RESET_B(net2092),
    .D(_01596_),
    .Q_N(_05205_),
    .Q(\shift_storage.storage [904]));
 sg13g2_dfrbp_1 \shift_storage.storage[905]$_SDFFE_PN0P_  (.CLK(clknet_leaf_255_clk_p2c),
    .RESET_B(net2093),
    .D(_01597_),
    .Q_N(_05204_),
    .Q(\shift_storage.storage [905]));
 sg13g2_dfrbp_1 \shift_storage.storage[906]$_SDFFE_PN0P_  (.CLK(clknet_leaf_253_clk_p2c),
    .RESET_B(net2094),
    .D(_01598_),
    .Q_N(_05203_),
    .Q(\shift_storage.storage [906]));
 sg13g2_dfrbp_1 \shift_storage.storage[907]$_SDFFE_PN0P_  (.CLK(clknet_leaf_255_clk_p2c),
    .RESET_B(net2095),
    .D(_01599_),
    .Q_N(_05202_),
    .Q(\shift_storage.storage [907]));
 sg13g2_dfrbp_1 \shift_storage.storage[908]$_SDFFE_PN0P_  (.CLK(clknet_leaf_253_clk_p2c),
    .RESET_B(net2096),
    .D(_01600_),
    .Q_N(_05201_),
    .Q(\shift_storage.storage [908]));
 sg13g2_dfrbp_1 \shift_storage.storage[909]$_SDFFE_PN0P_  (.CLK(clknet_leaf_253_clk_p2c),
    .RESET_B(net2097),
    .D(_01601_),
    .Q_N(_05200_),
    .Q(\shift_storage.storage [909]));
 sg13g2_dfrbp_1 \shift_storage.storage[90]$_SDFFE_PN0P_  (.CLK(clknet_leaf_255_clk_p2c),
    .RESET_B(net2098),
    .D(_01602_),
    .Q_N(_05199_),
    .Q(\shift_storage.storage [90]));
 sg13g2_dfrbp_1 \shift_storage.storage[910]$_SDFFE_PN0P_  (.CLK(clknet_leaf_254_clk_p2c),
    .RESET_B(net2099),
    .D(_01603_),
    .Q_N(_05198_),
    .Q(\shift_storage.storage [910]));
 sg13g2_dfrbp_1 \shift_storage.storage[911]$_SDFFE_PN0P_  (.CLK(clknet_leaf_254_clk_p2c),
    .RESET_B(net2100),
    .D(_01604_),
    .Q_N(_05197_),
    .Q(\shift_storage.storage [911]));
 sg13g2_dfrbp_1 \shift_storage.storage[912]$_SDFFE_PN0P_  (.CLK(clknet_leaf_254_clk_p2c),
    .RESET_B(net2101),
    .D(_01605_),
    .Q_N(_05196_),
    .Q(\shift_storage.storage [912]));
 sg13g2_dfrbp_1 \shift_storage.storage[913]$_SDFFE_PN0P_  (.CLK(clknet_leaf_254_clk_p2c),
    .RESET_B(net2102),
    .D(_01606_),
    .Q_N(_05195_),
    .Q(\shift_storage.storage [913]));
 sg13g2_dfrbp_1 \shift_storage.storage[914]$_SDFFE_PN0P_  (.CLK(clknet_leaf_254_clk_p2c),
    .RESET_B(net2103),
    .D(_01607_),
    .Q_N(_05194_),
    .Q(\shift_storage.storage [914]));
 sg13g2_dfrbp_1 \shift_storage.storage[915]$_SDFFE_PN0P_  (.CLK(clknet_leaf_254_clk_p2c),
    .RESET_B(net2104),
    .D(_01608_),
    .Q_N(_05193_),
    .Q(\shift_storage.storage [915]));
 sg13g2_dfrbp_1 \shift_storage.storage[916]$_SDFFE_PN0P_  (.CLK(clknet_leaf_38_clk_p2c),
    .RESET_B(net2105),
    .D(_01609_),
    .Q_N(_05192_),
    .Q(\shift_storage.storage [916]));
 sg13g2_dfrbp_1 \shift_storage.storage[917]$_SDFFE_PN0P_  (.CLK(clknet_leaf_38_clk_p2c),
    .RESET_B(net2106),
    .D(_01610_),
    .Q_N(_05191_),
    .Q(\shift_storage.storage [917]));
 sg13g2_dfrbp_1 \shift_storage.storage[918]$_SDFFE_PN0P_  (.CLK(clknet_leaf_37_clk_p2c),
    .RESET_B(net2107),
    .D(_01611_),
    .Q_N(_05190_),
    .Q(\shift_storage.storage [918]));
 sg13g2_dfrbp_1 \shift_storage.storage[919]$_SDFFE_PN0P_  (.CLK(clknet_leaf_255_clk_p2c),
    .RESET_B(net2108),
    .D(_01612_),
    .Q_N(_05189_),
    .Q(\shift_storage.storage [919]));
 sg13g2_dfrbp_1 \shift_storage.storage[91]$_SDFFE_PN0P_  (.CLK(clknet_leaf_37_clk_p2c),
    .RESET_B(net2109),
    .D(_01613_),
    .Q_N(_05188_),
    .Q(\shift_storage.storage [91]));
 sg13g2_dfrbp_1 \shift_storage.storage[920]$_SDFFE_PN0P_  (.CLK(clknet_leaf_256_clk_p2c),
    .RESET_B(net2110),
    .D(_01614_),
    .Q_N(_05187_),
    .Q(\shift_storage.storage [920]));
 sg13g2_dfrbp_1 \shift_storage.storage[921]$_SDFFE_PN0P_  (.CLK(clknet_leaf_256_clk_p2c),
    .RESET_B(net2111),
    .D(_01615_),
    .Q_N(_05186_),
    .Q(\shift_storage.storage [921]));
 sg13g2_dfrbp_1 \shift_storage.storage[922]$_SDFFE_PN0P_  (.CLK(clknet_leaf_256_clk_p2c),
    .RESET_B(net2112),
    .D(_01616_),
    .Q_N(_05185_),
    .Q(\shift_storage.storage [922]));
 sg13g2_dfrbp_1 \shift_storage.storage[923]$_SDFFE_PN0P_  (.CLK(clknet_leaf_257_clk_p2c),
    .RESET_B(net2113),
    .D(_01617_),
    .Q_N(_05184_),
    .Q(\shift_storage.storage [923]));
 sg13g2_dfrbp_1 \shift_storage.storage[924]$_SDFFE_PN0P_  (.CLK(clknet_leaf_256_clk_p2c),
    .RESET_B(net2114),
    .D(_01618_),
    .Q_N(_05183_),
    .Q(\shift_storage.storage [924]));
 sg13g2_dfrbp_1 \shift_storage.storage[925]$_SDFFE_PN0P_  (.CLK(clknet_leaf_36_clk_p2c),
    .RESET_B(net2115),
    .D(_01619_),
    .Q_N(_05182_),
    .Q(\shift_storage.storage [925]));
 sg13g2_dfrbp_1 \shift_storage.storage[926]$_SDFFE_PN0P_  (.CLK(clknet_leaf_36_clk_p2c),
    .RESET_B(net2116),
    .D(_01620_),
    .Q_N(_05181_),
    .Q(\shift_storage.storage [926]));
 sg13g2_dfrbp_1 \shift_storage.storage[927]$_SDFFE_PN0P_  (.CLK(clknet_leaf_36_clk_p2c),
    .RESET_B(net2117),
    .D(_01621_),
    .Q_N(_05180_),
    .Q(\shift_storage.storage [927]));
 sg13g2_dfrbp_1 \shift_storage.storage[928]$_SDFFE_PN0P_  (.CLK(clknet_leaf_36_clk_p2c),
    .RESET_B(net2118),
    .D(_01622_),
    .Q_N(_05179_),
    .Q(\shift_storage.storage [928]));
 sg13g2_dfrbp_1 \shift_storage.storage[929]$_SDFFE_PN0P_  (.CLK(clknet_leaf_36_clk_p2c),
    .RESET_B(net2119),
    .D(_01623_),
    .Q_N(_05178_),
    .Q(\shift_storage.storage [929]));
 sg13g2_dfrbp_1 \shift_storage.storage[92]$_SDFFE_PN0P_  (.CLK(clknet_leaf_37_clk_p2c),
    .RESET_B(net2120),
    .D(_01624_),
    .Q_N(_05177_),
    .Q(\shift_storage.storage [92]));
 sg13g2_dfrbp_1 \shift_storage.storage[930]$_SDFFE_PN0P_  (.CLK(clknet_leaf_36_clk_p2c),
    .RESET_B(net2121),
    .D(_01625_),
    .Q_N(_05176_),
    .Q(\shift_storage.storage [930]));
 sg13g2_dfrbp_1 \shift_storage.storage[931]$_SDFFE_PN0P_  (.CLK(clknet_leaf_12_clk_p2c),
    .RESET_B(net2122),
    .D(_01626_),
    .Q_N(_05175_),
    .Q(\shift_storage.storage [931]));
 sg13g2_dfrbp_1 \shift_storage.storage[932]$_SDFFE_PN0P_  (.CLK(clknet_leaf_35_clk_p2c),
    .RESET_B(net2123),
    .D(_01627_),
    .Q_N(_05174_),
    .Q(\shift_storage.storage [932]));
 sg13g2_dfrbp_1 \shift_storage.storage[933]$_SDFFE_PN0P_  (.CLK(clknet_leaf_35_clk_p2c),
    .RESET_B(net2124),
    .D(_01628_),
    .Q_N(_05173_),
    .Q(\shift_storage.storage [933]));
 sg13g2_dfrbp_1 \shift_storage.storage[934]$_SDFFE_PN0P_  (.CLK(clknet_leaf_35_clk_p2c),
    .RESET_B(net2125),
    .D(_01629_),
    .Q_N(_05172_),
    .Q(\shift_storage.storage [934]));
 sg13g2_dfrbp_1 \shift_storage.storage[935]$_SDFFE_PN0P_  (.CLK(clknet_leaf_35_clk_p2c),
    .RESET_B(net2126),
    .D(_01630_),
    .Q_N(_05171_),
    .Q(\shift_storage.storage [935]));
 sg13g2_dfrbp_1 \shift_storage.storage[936]$_SDFFE_PN0P_  (.CLK(clknet_leaf_37_clk_p2c),
    .RESET_B(net2127),
    .D(_01631_),
    .Q_N(_05170_),
    .Q(\shift_storage.storage [936]));
 sg13g2_dfrbp_1 \shift_storage.storage[937]$_SDFFE_PN0P_  (.CLK(clknet_leaf_35_clk_p2c),
    .RESET_B(net2128),
    .D(_01632_),
    .Q_N(_05169_),
    .Q(\shift_storage.storage [937]));
 sg13g2_dfrbp_1 \shift_storage.storage[938]$_SDFFE_PN0P_  (.CLK(clknet_leaf_34_clk_p2c),
    .RESET_B(net2129),
    .D(_01633_),
    .Q_N(_05168_),
    .Q(\shift_storage.storage [938]));
 sg13g2_dfrbp_1 \shift_storage.storage[939]$_SDFFE_PN0P_  (.CLK(clknet_leaf_34_clk_p2c),
    .RESET_B(net2130),
    .D(_01634_),
    .Q_N(_05167_),
    .Q(\shift_storage.storage [939]));
 sg13g2_dfrbp_1 \shift_storage.storage[93]$_SDFFE_PN0P_  (.CLK(clknet_leaf_32_clk_p2c),
    .RESET_B(net2131),
    .D(_01635_),
    .Q_N(_05166_),
    .Q(\shift_storage.storage [93]));
 sg13g2_dfrbp_1 \shift_storage.storage[940]$_SDFFE_PN0P_  (.CLK(clknet_leaf_34_clk_p2c),
    .RESET_B(net2132),
    .D(_01636_),
    .Q_N(_05165_),
    .Q(\shift_storage.storage [940]));
 sg13g2_dfrbp_1 \shift_storage.storage[941]$_SDFFE_PN0P_  (.CLK(clknet_leaf_34_clk_p2c),
    .RESET_B(net2133),
    .D(_01637_),
    .Q_N(_05164_),
    .Q(\shift_storage.storage [941]));
 sg13g2_dfrbp_1 \shift_storage.storage[942]$_SDFFE_PN0P_  (.CLK(clknet_leaf_32_clk_p2c),
    .RESET_B(net2134),
    .D(_01638_),
    .Q_N(_05163_),
    .Q(\shift_storage.storage [942]));
 sg13g2_dfrbp_1 \shift_storage.storage[943]$_SDFFE_PN0P_  (.CLK(clknet_leaf_33_clk_p2c),
    .RESET_B(net2135),
    .D(_01639_),
    .Q_N(_05162_),
    .Q(\shift_storage.storage [943]));
 sg13g2_dfrbp_1 \shift_storage.storage[944]$_SDFFE_PN0P_  (.CLK(clknet_leaf_32_clk_p2c),
    .RESET_B(net2136),
    .D(_01640_),
    .Q_N(_05161_),
    .Q(\shift_storage.storage [944]));
 sg13g2_dfrbp_1 \shift_storage.storage[945]$_SDFFE_PN0P_  (.CLK(clknet_leaf_32_clk_p2c),
    .RESET_B(net2137),
    .D(_01641_),
    .Q_N(_05160_),
    .Q(\shift_storage.storage [945]));
 sg13g2_dfrbp_1 \shift_storage.storage[946]$_SDFFE_PN0P_  (.CLK(clknet_leaf_31_clk_p2c),
    .RESET_B(net2138),
    .D(_01642_),
    .Q_N(_05159_),
    .Q(\shift_storage.storage [946]));
 sg13g2_dfrbp_1 \shift_storage.storage[947]$_SDFFE_PN0P_  (.CLK(clknet_leaf_31_clk_p2c),
    .RESET_B(net2139),
    .D(_01643_),
    .Q_N(_05158_),
    .Q(\shift_storage.storage [947]));
 sg13g2_dfrbp_1 \shift_storage.storage[948]$_SDFFE_PN0P_  (.CLK(clknet_leaf_30_clk_p2c),
    .RESET_B(net2140),
    .D(_01644_),
    .Q_N(_05157_),
    .Q(\shift_storage.storage [948]));
 sg13g2_dfrbp_1 \shift_storage.storage[949]$_SDFFE_PN0P_  (.CLK(clknet_leaf_32_clk_p2c),
    .RESET_B(net2141),
    .D(_01645_),
    .Q_N(_05156_),
    .Q(\shift_storage.storage [949]));
 sg13g2_dfrbp_1 \shift_storage.storage[94]$_SDFFE_PN0P_  (.CLK(clknet_leaf_31_clk_p2c),
    .RESET_B(net2142),
    .D(_01646_),
    .Q_N(_05155_),
    .Q(\shift_storage.storage [94]));
 sg13g2_dfrbp_1 \shift_storage.storage[950]$_SDFFE_PN0P_  (.CLK(clknet_leaf_31_clk_p2c),
    .RESET_B(net2143),
    .D(_01647_),
    .Q_N(_05154_),
    .Q(\shift_storage.storage [950]));
 sg13g2_dfrbp_1 \shift_storage.storage[951]$_SDFFE_PN0P_  (.CLK(clknet_leaf_31_clk_p2c),
    .RESET_B(net2144),
    .D(_01648_),
    .Q_N(_05153_),
    .Q(\shift_storage.storage [951]));
 sg13g2_dfrbp_1 \shift_storage.storage[952]$_SDFFE_PN0P_  (.CLK(clknet_leaf_30_clk_p2c),
    .RESET_B(net2145),
    .D(_01649_),
    .Q_N(_05152_),
    .Q(\shift_storage.storage [952]));
 sg13g2_dfrbp_1 \shift_storage.storage[953]$_SDFFE_PN0P_  (.CLK(clknet_leaf_29_clk_p2c),
    .RESET_B(net2146),
    .D(_01650_),
    .Q_N(_05151_),
    .Q(\shift_storage.storage [953]));
 sg13g2_dfrbp_1 \shift_storage.storage[954]$_SDFFE_PN0P_  (.CLK(clknet_leaf_29_clk_p2c),
    .RESET_B(net2147),
    .D(_01651_),
    .Q_N(_05150_),
    .Q(\shift_storage.storage [954]));
 sg13g2_dfrbp_1 \shift_storage.storage[955]$_SDFFE_PN0P_  (.CLK(clknet_leaf_30_clk_p2c),
    .RESET_B(net2148),
    .D(_01652_),
    .Q_N(_05149_),
    .Q(\shift_storage.storage [955]));
 sg13g2_dfrbp_1 \shift_storage.storage[956]$_SDFFE_PN0P_  (.CLK(clknet_leaf_30_clk_p2c),
    .RESET_B(net2149),
    .D(_01653_),
    .Q_N(_05148_),
    .Q(\shift_storage.storage [956]));
 sg13g2_dfrbp_1 \shift_storage.storage[957]$_SDFFE_PN0P_  (.CLK(clknet_leaf_30_clk_p2c),
    .RESET_B(net2150),
    .D(_01654_),
    .Q_N(_05147_),
    .Q(\shift_storage.storage [957]));
 sg13g2_dfrbp_1 \shift_storage.storage[958]$_SDFFE_PN0P_  (.CLK(clknet_leaf_30_clk_p2c),
    .RESET_B(net2151),
    .D(_01655_),
    .Q_N(_05146_),
    .Q(\shift_storage.storage [958]));
 sg13g2_dfrbp_1 \shift_storage.storage[959]$_SDFFE_PN0P_  (.CLK(clknet_leaf_65_clk_p2c),
    .RESET_B(net2152),
    .D(_01656_),
    .Q_N(_05145_),
    .Q(\shift_storage.storage [959]));
 sg13g2_dfrbp_1 \shift_storage.storage[95]$_SDFFE_PN0P_  (.CLK(clknet_leaf_40_clk_p2c),
    .RESET_B(net2153),
    .D(_01657_),
    .Q_N(_05144_),
    .Q(\shift_storage.storage [95]));
 sg13g2_dfrbp_1 \shift_storage.storage[960]$_SDFFE_PN0P_  (.CLK(clknet_leaf_65_clk_p2c),
    .RESET_B(net2154),
    .D(_01658_),
    .Q_N(_05143_),
    .Q(\shift_storage.storage [960]));
 sg13g2_dfrbp_1 \shift_storage.storage[961]$_SDFFE_PN0P_  (.CLK(clknet_leaf_52_clk_p2c),
    .RESET_B(net2155),
    .D(_01659_),
    .Q_N(_05142_),
    .Q(\shift_storage.storage [961]));
 sg13g2_dfrbp_1 \shift_storage.storage[962]$_SDFFE_PN0P_  (.CLK(clknet_leaf_53_clk_p2c),
    .RESET_B(net2156),
    .D(_01660_),
    .Q_N(_05141_),
    .Q(\shift_storage.storage [962]));
 sg13g2_dfrbp_1 \shift_storage.storage[963]$_SDFFE_PN0P_  (.CLK(clknet_leaf_53_clk_p2c),
    .RESET_B(net2157),
    .D(_01661_),
    .Q_N(_05140_),
    .Q(\shift_storage.storage [963]));
 sg13g2_dfrbp_1 \shift_storage.storage[964]$_SDFFE_PN0P_  (.CLK(clknet_leaf_41_clk_p2c),
    .RESET_B(net2158),
    .D(_01662_),
    .Q_N(_05139_),
    .Q(\shift_storage.storage [964]));
 sg13g2_dfrbp_1 \shift_storage.storage[965]$_SDFFE_PN0P_  (.CLK(clknet_leaf_41_clk_p2c),
    .RESET_B(net2159),
    .D(_01663_),
    .Q_N(_05138_),
    .Q(\shift_storage.storage [965]));
 sg13g2_dfrbp_1 \shift_storage.storage[966]$_SDFFE_PN0P_  (.CLK(clknet_leaf_41_clk_p2c),
    .RESET_B(net2160),
    .D(_01664_),
    .Q_N(_05137_),
    .Q(\shift_storage.storage [966]));
 sg13g2_dfrbp_1 \shift_storage.storage[967]$_SDFFE_PN0P_  (.CLK(clknet_leaf_41_clk_p2c),
    .RESET_B(net2161),
    .D(_01665_),
    .Q_N(_05136_),
    .Q(\shift_storage.storage [967]));
 sg13g2_dfrbp_1 \shift_storage.storage[968]$_SDFFE_PN0P_  (.CLK(clknet_leaf_41_clk_p2c),
    .RESET_B(net2162),
    .D(_01666_),
    .Q_N(_05135_),
    .Q(\shift_storage.storage [968]));
 sg13g2_dfrbp_1 \shift_storage.storage[969]$_SDFFE_PN0P_  (.CLK(clknet_leaf_40_clk_p2c),
    .RESET_B(net2163),
    .D(_01667_),
    .Q_N(_05134_),
    .Q(\shift_storage.storage [969]));
 sg13g2_dfrbp_1 \shift_storage.storage[96]$_SDFFE_PN0P_  (.CLK(clknet_leaf_40_clk_p2c),
    .RESET_B(net2164),
    .D(_01668_),
    .Q_N(_05133_),
    .Q(\shift_storage.storage [96]));
 sg13g2_dfrbp_1 \shift_storage.storage[970]$_SDFFE_PN0P_  (.CLK(clknet_leaf_39_clk_p2c),
    .RESET_B(net2165),
    .D(_01669_),
    .Q_N(_05132_),
    .Q(\shift_storage.storage [970]));
 sg13g2_dfrbp_1 \shift_storage.storage[971]$_SDFFE_PN0P_  (.CLK(clknet_leaf_39_clk_p2c),
    .RESET_B(net2166),
    .D(_01670_),
    .Q_N(_05131_),
    .Q(\shift_storage.storage [971]));
 sg13g2_dfrbp_1 \shift_storage.storage[972]$_SDFFE_PN0P_  (.CLK(clknet_leaf_40_clk_p2c),
    .RESET_B(net2167),
    .D(_01671_),
    .Q_N(_05130_),
    .Q(\shift_storage.storage [972]));
 sg13g2_dfrbp_1 \shift_storage.storage[973]$_SDFFE_PN0P_  (.CLK(clknet_leaf_40_clk_p2c),
    .RESET_B(net2168),
    .D(_01672_),
    .Q_N(_05129_),
    .Q(\shift_storage.storage [973]));
 sg13g2_dfrbp_1 \shift_storage.storage[974]$_SDFFE_PN0P_  (.CLK(clknet_leaf_40_clk_p2c),
    .RESET_B(net2169),
    .D(_01673_),
    .Q_N(_05128_),
    .Q(\shift_storage.storage [974]));
 sg13g2_dfrbp_1 \shift_storage.storage[975]$_SDFFE_PN0P_  (.CLK(clknet_leaf_37_clk_p2c),
    .RESET_B(net2170),
    .D(_01674_),
    .Q_N(_05127_),
    .Q(\shift_storage.storage [975]));
 sg13g2_dfrbp_1 \shift_storage.storage[976]$_SDFFE_PN0P_  (.CLK(clknet_leaf_37_clk_p2c),
    .RESET_B(net2171),
    .D(_01675_),
    .Q_N(_05126_),
    .Q(\shift_storage.storage [976]));
 sg13g2_dfrbp_1 \shift_storage.storage[977]$_SDFFE_PN0P_  (.CLK(clknet_leaf_37_clk_p2c),
    .RESET_B(net2172),
    .D(_01676_),
    .Q_N(_05125_),
    .Q(\shift_storage.storage [977]));
 sg13g2_dfrbp_1 \shift_storage.storage[978]$_SDFFE_PN0P_  (.CLK(clknet_leaf_38_clk_p2c),
    .RESET_B(net2173),
    .D(_01677_),
    .Q_N(_05124_),
    .Q(\shift_storage.storage [978]));
 sg13g2_dfrbp_1 \shift_storage.storage[979]$_SDFFE_PN0P_  (.CLK(clknet_leaf_38_clk_p2c),
    .RESET_B(net2174),
    .D(_01678_),
    .Q_N(_05123_),
    .Q(\shift_storage.storage [979]));
 sg13g2_dfrbp_1 \shift_storage.storage[97]$_SDFFE_PN0P_  (.CLK(clknet_leaf_42_clk_p2c),
    .RESET_B(net2175),
    .D(_01679_),
    .Q_N(_05122_),
    .Q(\shift_storage.storage [97]));
 sg13g2_dfrbp_1 \shift_storage.storage[980]$_SDFFE_PN0P_  (.CLK(clknet_leaf_38_clk_p2c),
    .RESET_B(net2176),
    .D(_01680_),
    .Q_N(_05121_),
    .Q(\shift_storage.storage [980]));
 sg13g2_dfrbp_1 \shift_storage.storage[981]$_SDFFE_PN0P_  (.CLK(clknet_leaf_39_clk_p2c),
    .RESET_B(net2177),
    .D(_01681_),
    .Q_N(_05120_),
    .Q(\shift_storage.storage [981]));
 sg13g2_dfrbp_1 \shift_storage.storage[982]$_SDFFE_PN0P_  (.CLK(clknet_leaf_39_clk_p2c),
    .RESET_B(net2178),
    .D(_01682_),
    .Q_N(_05119_),
    .Q(\shift_storage.storage [982]));
 sg13g2_dfrbp_1 \shift_storage.storage[983]$_SDFFE_PN0P_  (.CLK(clknet_leaf_44_clk_p2c),
    .RESET_B(net2179),
    .D(_01683_),
    .Q_N(_05118_),
    .Q(\shift_storage.storage [983]));
 sg13g2_dfrbp_1 \shift_storage.storage[984]$_SDFFE_PN0P_  (.CLK(clknet_leaf_44_clk_p2c),
    .RESET_B(net2180),
    .D(_01684_),
    .Q_N(_05117_),
    .Q(\shift_storage.storage [984]));
 sg13g2_dfrbp_1 \shift_storage.storage[985]$_SDFFE_PN0P_  (.CLK(clknet_leaf_44_clk_p2c),
    .RESET_B(net2181),
    .D(_01685_),
    .Q_N(_05116_),
    .Q(\shift_storage.storage [985]));
 sg13g2_dfrbp_1 \shift_storage.storage[986]$_SDFFE_PN0P_  (.CLK(clknet_leaf_39_clk_p2c),
    .RESET_B(net2182),
    .D(_01686_),
    .Q_N(_05115_),
    .Q(\shift_storage.storage [986]));
 sg13g2_dfrbp_1 \shift_storage.storage[987]$_SDFFE_PN0P_  (.CLK(clknet_leaf_44_clk_p2c),
    .RESET_B(net2183),
    .D(_01687_),
    .Q_N(_05114_),
    .Q(\shift_storage.storage [987]));
 sg13g2_dfrbp_1 \shift_storage.storage[988]$_SDFFE_PN0P_  (.CLK(clknet_leaf_43_clk_p2c),
    .RESET_B(net2184),
    .D(_01688_),
    .Q_N(_05113_),
    .Q(\shift_storage.storage [988]));
 sg13g2_dfrbp_1 \shift_storage.storage[989]$_SDFFE_PN0P_  (.CLK(clknet_leaf_42_clk_p2c),
    .RESET_B(net2185),
    .D(_01689_),
    .Q_N(_05112_),
    .Q(\shift_storage.storage [989]));
 sg13g2_dfrbp_1 \shift_storage.storage[98]$_SDFFE_PN0P_  (.CLK(clknet_leaf_43_clk_p2c),
    .RESET_B(net2186),
    .D(_01690_),
    .Q_N(_05111_),
    .Q(\shift_storage.storage [98]));
 sg13g2_dfrbp_1 \shift_storage.storage[990]$_SDFFE_PN0P_  (.CLK(clknet_leaf_42_clk_p2c),
    .RESET_B(net2187),
    .D(_01691_),
    .Q_N(_05110_),
    .Q(\shift_storage.storage [990]));
 sg13g2_dfrbp_1 \shift_storage.storage[991]$_SDFFE_PN0P_  (.CLK(clknet_leaf_43_clk_p2c),
    .RESET_B(net2188),
    .D(_01692_),
    .Q_N(_05109_),
    .Q(\shift_storage.storage [991]));
 sg13g2_dfrbp_1 \shift_storage.storage[992]$_SDFFE_PN0P_  (.CLK(clknet_leaf_44_clk_p2c),
    .RESET_B(net2189),
    .D(_01693_),
    .Q_N(_05108_),
    .Q(\shift_storage.storage [992]));
 sg13g2_dfrbp_1 \shift_storage.storage[993]$_SDFFE_PN0P_  (.CLK(clknet_leaf_44_clk_p2c),
    .RESET_B(net2190),
    .D(_01694_),
    .Q_N(_05107_),
    .Q(\shift_storage.storage [993]));
 sg13g2_dfrbp_1 \shift_storage.storage[994]$_SDFFE_PN0P_  (.CLK(clknet_leaf_45_clk_p2c),
    .RESET_B(net2191),
    .D(_01695_),
    .Q_N(_05106_),
    .Q(\shift_storage.storage [994]));
 sg13g2_dfrbp_1 \shift_storage.storage[995]$_SDFFE_PN0P_  (.CLK(clknet_leaf_45_clk_p2c),
    .RESET_B(net2192),
    .D(_01696_),
    .Q_N(_05105_),
    .Q(\shift_storage.storage [995]));
 sg13g2_dfrbp_1 \shift_storage.storage[996]$_SDFFE_PN0P_  (.CLK(clknet_leaf_45_clk_p2c),
    .RESET_B(net2193),
    .D(_01697_),
    .Q_N(_05104_),
    .Q(\shift_storage.storage [996]));
 sg13g2_dfrbp_1 \shift_storage.storage[997]$_SDFFE_PN0P_  (.CLK(clknet_leaf_45_clk_p2c),
    .RESET_B(net2194),
    .D(_01698_),
    .Q_N(_05103_),
    .Q(\shift_storage.storage [997]));
 sg13g2_dfrbp_1 \shift_storage.storage[998]$_SDFFE_PN0P_  (.CLK(clknet_leaf_45_clk_p2c),
    .RESET_B(net2195),
    .D(_01699_),
    .Q_N(_05102_),
    .Q(\shift_storage.storage [998]));
 sg13g2_dfrbp_1 \shift_storage.storage[999]$_SDFFE_PN0P_  (.CLK(clknet_leaf_46_clk_p2c),
    .RESET_B(net2196),
    .D(_01700_),
    .Q_N(_05101_),
    .Q(\shift_storage.storage [999]));
 sg13g2_dfrbp_1 \shift_storage.storage[99]$_SDFFE_PN0P_  (.CLK(clknet_leaf_43_clk_p2c),
    .RESET_B(net2197),
    .D(_01701_),
    .Q_N(_05100_),
    .Q(\shift_storage.storage [99]));
 sg13g2_dfrbp_1 \shift_storage.storage[9]$_SDFFE_PN0P_  (.CLK(clknet_leaf_45_clk_p2c),
    .RESET_B(net2198),
    .D(_01702_),
    .Q_N(_05099_),
    .Q(\shift_storage.storage [9]));
 sg13g2_IOPadVdd VDD ();
 sg13g2_IOPadIOVdd IOVDD ();
 sg13g2_IOPadVss VSS ();
 sg13g2_IOPadIOVss IOVSS ();
 sg13g2_Corner IO_CORNER_NORTH_WEST_INST ();
 sg13g2_Corner IO_CORNER_NORTH_EAST_INST ();
 sg13g2_Corner IO_CORNER_SOUTH_WEST_INST ();
 sg13g2_Corner IO_CORNER_SOUTH_EAST_INST ();
 sg13g2_Filler200 IO_FILL_IO_NORTH_0_0 ();
 sg13g2_Filler200 IO_FILL_IO_NORTH_0_1 ();
 sg13g2_Filler200 IO_FILL_IO_NORTH_0_2 ();
 sg13g2_Filler200 IO_FILL_IO_NORTH_0_3 ();
 sg13g2_Filler200 IO_FILL_IO_NORTH_0_4 ();
 sg13g2_Filler200 IO_FILL_IO_NORTH_0_5 ();
 sg13g2_Filler200 IO_FILL_IO_NORTH_0_6 ();
 sg13g2_Filler200 IO_FILL_IO_NORTH_0_7 ();
 sg13g2_Filler200 IO_FILL_IO_NORTH_0_8 ();
 sg13g2_Filler200 IO_FILL_IO_NORTH_0_9 ();
 sg13g2_Filler200 IO_FILL_IO_NORTH_1_0 ();
 sg13g2_Filler200 IO_FILL_IO_NORTH_1_1 ();
 sg13g2_Filler200 IO_FILL_IO_NORTH_1_2 ();
 sg13g2_Filler200 IO_FILL_IO_NORTH_1_3 ();
 sg13g2_Filler200 IO_FILL_IO_NORTH_1_4 ();
 sg13g2_Filler200 IO_FILL_IO_NORTH_1_5 ();
 sg13g2_Filler200 IO_FILL_IO_NORTH_1_6 ();
 sg13g2_Filler200 IO_FILL_IO_NORTH_1_7 ();
 sg13g2_Filler200 IO_FILL_IO_NORTH_1_8 ();
 sg13g2_Filler200 IO_FILL_IO_NORTH_1_9 ();
 sg13g2_Filler200 IO_FILL_IO_NORTH_2_0 ();
 sg13g2_Filler200 IO_FILL_IO_NORTH_2_1 ();
 sg13g2_Filler200 IO_FILL_IO_NORTH_2_2 ();
 sg13g2_Filler200 IO_FILL_IO_NORTH_2_3 ();
 sg13g2_Filler200 IO_FILL_IO_NORTH_2_4 ();
 sg13g2_Filler200 IO_FILL_IO_NORTH_2_5 ();
 sg13g2_Filler200 IO_FILL_IO_NORTH_2_6 ();
 sg13g2_Filler200 IO_FILL_IO_NORTH_2_7 ();
 sg13g2_Filler200 IO_FILL_IO_NORTH_2_8 ();
 sg13g2_Filler200 IO_FILL_IO_NORTH_2_9 ();
 sg13g2_Filler200 IO_FILL_IO_NORTH_3_0 ();
 sg13g2_Filler200 IO_FILL_IO_NORTH_3_1 ();
 sg13g2_Filler200 IO_FILL_IO_NORTH_3_2 ();
 sg13g2_Filler200 IO_FILL_IO_NORTH_3_3 ();
 sg13g2_Filler200 IO_FILL_IO_NORTH_3_4 ();
 sg13g2_Filler200 IO_FILL_IO_NORTH_3_5 ();
 sg13g2_Filler200 IO_FILL_IO_NORTH_3_6 ();
 sg13g2_Filler200 IO_FILL_IO_NORTH_3_7 ();
 sg13g2_Filler200 IO_FILL_IO_NORTH_3_8 ();
 sg13g2_Filler200 IO_FILL_IO_NORTH_3_9 ();
 sg13g2_Filler200 IO_FILL_IO_NORTH_4_0 ();
 sg13g2_Filler200 IO_FILL_IO_NORTH_4_1 ();
 sg13g2_Filler200 IO_FILL_IO_NORTH_4_2 ();
 sg13g2_Filler200 IO_FILL_IO_NORTH_4_3 ();
 sg13g2_Filler200 IO_FILL_IO_NORTH_4_4 ();
 sg13g2_Filler200 IO_FILL_IO_NORTH_4_5 ();
 sg13g2_Filler200 IO_FILL_IO_NORTH_4_6 ();
 sg13g2_Filler200 IO_FILL_IO_NORTH_4_7 ();
 sg13g2_Filler200 IO_FILL_IO_NORTH_4_8 ();
 sg13g2_Filler200 IO_FILL_IO_NORTH_4_9 ();
 sg13g2_Filler200 IO_FILL_IO_NORTH_5_0 ();
 sg13g2_Filler200 IO_FILL_IO_NORTH_5_1 ();
 sg13g2_Filler200 IO_FILL_IO_NORTH_5_2 ();
 sg13g2_Filler200 IO_FILL_IO_NORTH_5_3 ();
 sg13g2_Filler200 IO_FILL_IO_NORTH_5_4 ();
 sg13g2_Filler200 IO_FILL_IO_NORTH_5_5 ();
 sg13g2_Filler200 IO_FILL_IO_NORTH_5_6 ();
 sg13g2_Filler200 IO_FILL_IO_NORTH_5_7 ();
 sg13g2_Filler200 IO_FILL_IO_NORTH_5_8 ();
 sg13g2_Filler200 IO_FILL_IO_NORTH_5_9 ();
 sg13g2_Filler200 IO_FILL_IO_NORTH_6_0 ();
 sg13g2_Filler200 IO_FILL_IO_NORTH_6_1 ();
 sg13g2_Filler200 IO_FILL_IO_NORTH_6_2 ();
 sg13g2_Filler200 IO_FILL_IO_NORTH_6_3 ();
 sg13g2_Filler200 IO_FILL_IO_NORTH_6_4 ();
 sg13g2_Filler200 IO_FILL_IO_NORTH_6_5 ();
 sg13g2_Filler200 IO_FILL_IO_NORTH_6_6 ();
 sg13g2_Filler200 IO_FILL_IO_NORTH_6_7 ();
 sg13g2_Filler200 IO_FILL_IO_NORTH_6_8 ();
 sg13g2_Filler200 IO_FILL_IO_NORTH_6_9 ();
 sg13g2_Filler200 IO_FILL_IO_NORTH_7_0 ();
 sg13g2_Filler200 IO_FILL_IO_NORTH_7_1 ();
 sg13g2_Filler200 IO_FILL_IO_NORTH_7_2 ();
 sg13g2_Filler200 IO_FILL_IO_NORTH_7_3 ();
 sg13g2_Filler200 IO_FILL_IO_NORTH_7_4 ();
 sg13g2_Filler200 IO_FILL_IO_NORTH_7_5 ();
 sg13g2_Filler200 IO_FILL_IO_NORTH_7_6 ();
 sg13g2_Filler200 IO_FILL_IO_NORTH_7_7 ();
 sg13g2_Filler200 IO_FILL_IO_NORTH_7_8 ();
 sg13g2_Filler200 IO_FILL_IO_NORTH_7_9 ();
 sg13g2_Filler200 IO_FILL_IO_NORTH_8_0 ();
 sg13g2_Filler200 IO_FILL_IO_NORTH_8_1 ();
 sg13g2_Filler200 IO_FILL_IO_NORTH_8_2 ();
 sg13g2_Filler200 IO_FILL_IO_NORTH_8_3 ();
 sg13g2_Filler200 IO_FILL_IO_NORTH_8_4 ();
 sg13g2_Filler200 IO_FILL_IO_NORTH_8_5 ();
 sg13g2_Filler200 IO_FILL_IO_NORTH_8_6 ();
 sg13g2_Filler200 IO_FILL_IO_NORTH_8_7 ();
 sg13g2_Filler200 IO_FILL_IO_NORTH_8_8 ();
 sg13g2_Filler200 IO_FILL_IO_NORTH_8_9 ();
 sg13g2_Filler200 IO_FILL_IO_SOUTH_0_0 ();
 sg13g2_Filler200 IO_FILL_IO_SOUTH_0_1 ();
 sg13g2_Filler200 IO_FILL_IO_SOUTH_0_2 ();
 sg13g2_Filler200 IO_FILL_IO_SOUTH_0_3 ();
 sg13g2_Filler200 IO_FILL_IO_SOUTH_0_4 ();
 sg13g2_Filler200 IO_FILL_IO_SOUTH_0_5 ();
 sg13g2_Filler200 IO_FILL_IO_SOUTH_0_6 ();
 sg13g2_Filler200 IO_FILL_IO_SOUTH_0_7 ();
 sg13g2_Filler200 IO_FILL_IO_SOUTH_0_8 ();
 sg13g2_Filler200 IO_FILL_IO_SOUTH_0_9 ();
 sg13g2_Filler200 IO_FILL_IO_SOUTH_1_0 ();
 sg13g2_Filler200 IO_FILL_IO_SOUTH_1_1 ();
 sg13g2_Filler200 IO_FILL_IO_SOUTH_1_2 ();
 sg13g2_Filler200 IO_FILL_IO_SOUTH_1_3 ();
 sg13g2_Filler200 IO_FILL_IO_SOUTH_1_4 ();
 sg13g2_Filler200 IO_FILL_IO_SOUTH_1_5 ();
 sg13g2_Filler200 IO_FILL_IO_SOUTH_1_6 ();
 sg13g2_Filler200 IO_FILL_IO_SOUTH_1_7 ();
 sg13g2_Filler200 IO_FILL_IO_SOUTH_1_8 ();
 sg13g2_Filler200 IO_FILL_IO_SOUTH_1_9 ();
 sg13g2_Filler200 IO_FILL_IO_SOUTH_2_0 ();
 sg13g2_Filler200 IO_FILL_IO_SOUTH_2_1 ();
 sg13g2_Filler200 IO_FILL_IO_SOUTH_2_2 ();
 sg13g2_Filler200 IO_FILL_IO_SOUTH_2_3 ();
 sg13g2_Filler200 IO_FILL_IO_SOUTH_2_4 ();
 sg13g2_Filler200 IO_FILL_IO_SOUTH_2_5 ();
 sg13g2_Filler200 IO_FILL_IO_SOUTH_2_6 ();
 sg13g2_Filler200 IO_FILL_IO_SOUTH_2_7 ();
 sg13g2_Filler200 IO_FILL_IO_SOUTH_2_8 ();
 sg13g2_Filler200 IO_FILL_IO_SOUTH_2_9 ();
 sg13g2_Filler200 IO_FILL_IO_SOUTH_3_0 ();
 sg13g2_Filler200 IO_FILL_IO_SOUTH_3_1 ();
 sg13g2_Filler200 IO_FILL_IO_SOUTH_3_2 ();
 sg13g2_Filler200 IO_FILL_IO_SOUTH_3_3 ();
 sg13g2_Filler200 IO_FILL_IO_SOUTH_3_4 ();
 sg13g2_Filler200 IO_FILL_IO_SOUTH_3_5 ();
 sg13g2_Filler200 IO_FILL_IO_SOUTH_3_6 ();
 sg13g2_Filler200 IO_FILL_IO_SOUTH_3_7 ();
 sg13g2_Filler200 IO_FILL_IO_SOUTH_3_8 ();
 sg13g2_Filler200 IO_FILL_IO_SOUTH_3_9 ();
 sg13g2_Filler200 IO_FILL_IO_SOUTH_4_0 ();
 sg13g2_Filler200 IO_FILL_IO_SOUTH_4_1 ();
 sg13g2_Filler200 IO_FILL_IO_SOUTH_4_2 ();
 sg13g2_Filler200 IO_FILL_IO_SOUTH_4_3 ();
 sg13g2_Filler200 IO_FILL_IO_SOUTH_4_4 ();
 sg13g2_Filler200 IO_FILL_IO_SOUTH_4_5 ();
 sg13g2_Filler200 IO_FILL_IO_SOUTH_4_6 ();
 sg13g2_Filler200 IO_FILL_IO_SOUTH_4_7 ();
 sg13g2_Filler200 IO_FILL_IO_SOUTH_4_8 ();
 sg13g2_Filler200 IO_FILL_IO_SOUTH_4_9 ();
 sg13g2_Filler200 IO_FILL_IO_SOUTH_5_0 ();
 sg13g2_Filler200 IO_FILL_IO_SOUTH_5_1 ();
 sg13g2_Filler200 IO_FILL_IO_SOUTH_5_2 ();
 sg13g2_Filler200 IO_FILL_IO_SOUTH_5_3 ();
 sg13g2_Filler200 IO_FILL_IO_SOUTH_5_4 ();
 sg13g2_Filler200 IO_FILL_IO_SOUTH_5_5 ();
 sg13g2_Filler200 IO_FILL_IO_SOUTH_5_6 ();
 sg13g2_Filler200 IO_FILL_IO_SOUTH_5_7 ();
 sg13g2_Filler200 IO_FILL_IO_SOUTH_5_8 ();
 sg13g2_Filler200 IO_FILL_IO_SOUTH_5_9 ();
 sg13g2_Filler200 IO_FILL_IO_SOUTH_6_0 ();
 sg13g2_Filler200 IO_FILL_IO_SOUTH_6_1 ();
 sg13g2_Filler200 IO_FILL_IO_SOUTH_6_2 ();
 sg13g2_Filler200 IO_FILL_IO_SOUTH_6_3 ();
 sg13g2_Filler200 IO_FILL_IO_SOUTH_6_4 ();
 sg13g2_Filler200 IO_FILL_IO_SOUTH_6_5 ();
 sg13g2_Filler200 IO_FILL_IO_SOUTH_6_6 ();
 sg13g2_Filler200 IO_FILL_IO_SOUTH_6_7 ();
 sg13g2_Filler200 IO_FILL_IO_SOUTH_6_8 ();
 sg13g2_Filler200 IO_FILL_IO_SOUTH_6_9 ();
 sg13g2_Filler200 IO_FILL_IO_SOUTH_7_0 ();
 sg13g2_Filler200 IO_FILL_IO_SOUTH_7_1 ();
 sg13g2_Filler200 IO_FILL_IO_SOUTH_7_2 ();
 sg13g2_Filler200 IO_FILL_IO_SOUTH_7_3 ();
 sg13g2_Filler200 IO_FILL_IO_SOUTH_7_4 ();
 sg13g2_Filler200 IO_FILL_IO_SOUTH_7_5 ();
 sg13g2_Filler200 IO_FILL_IO_SOUTH_7_6 ();
 sg13g2_Filler200 IO_FILL_IO_SOUTH_7_7 ();
 sg13g2_Filler200 IO_FILL_IO_SOUTH_7_8 ();
 sg13g2_Filler200 IO_FILL_IO_SOUTH_7_9 ();
 sg13g2_Filler200 IO_FILL_IO_SOUTH_8_0 ();
 sg13g2_Filler200 IO_FILL_IO_SOUTH_8_1 ();
 sg13g2_Filler200 IO_FILL_IO_SOUTH_8_2 ();
 sg13g2_Filler200 IO_FILL_IO_SOUTH_8_3 ();
 sg13g2_Filler200 IO_FILL_IO_SOUTH_8_4 ();
 sg13g2_Filler200 IO_FILL_IO_SOUTH_8_5 ();
 sg13g2_Filler200 IO_FILL_IO_SOUTH_8_6 ();
 sg13g2_Filler200 IO_FILL_IO_SOUTH_8_7 ();
 sg13g2_Filler200 IO_FILL_IO_SOUTH_8_8 ();
 sg13g2_Filler200 IO_FILL_IO_SOUTH_8_9 ();
 sg13g2_Filler200 IO_FILL_IO_WEST_0_0 ();
 sg13g2_Filler200 IO_FILL_IO_WEST_0_1 ();
 sg13g2_Filler200 IO_FILL_IO_WEST_0_2 ();
 sg13g2_Filler200 IO_FILL_IO_WEST_0_3 ();
 sg13g2_Filler200 IO_FILL_IO_WEST_0_4 ();
 sg13g2_Filler200 IO_FILL_IO_WEST_0_5 ();
 sg13g2_Filler200 IO_FILL_IO_WEST_0_6 ();
 sg13g2_Filler200 IO_FILL_IO_WEST_0_7 ();
 sg13g2_Filler200 IO_FILL_IO_WEST_0_8 ();
 sg13g2_Filler200 IO_FILL_IO_WEST_0_9 ();
 sg13g2_Filler200 IO_FILL_IO_WEST_1_0 ();
 sg13g2_Filler200 IO_FILL_IO_WEST_1_1 ();
 sg13g2_Filler200 IO_FILL_IO_WEST_1_2 ();
 sg13g2_Filler200 IO_FILL_IO_WEST_1_3 ();
 sg13g2_Filler200 IO_FILL_IO_WEST_1_4 ();
 sg13g2_Filler200 IO_FILL_IO_WEST_1_5 ();
 sg13g2_Filler200 IO_FILL_IO_WEST_1_6 ();
 sg13g2_Filler200 IO_FILL_IO_WEST_1_7 ();
 sg13g2_Filler200 IO_FILL_IO_WEST_1_8 ();
 sg13g2_Filler200 IO_FILL_IO_WEST_1_9 ();
 sg13g2_Filler200 IO_FILL_IO_WEST_2_0 ();
 sg13g2_Filler200 IO_FILL_IO_WEST_2_1 ();
 sg13g2_Filler200 IO_FILL_IO_WEST_2_2 ();
 sg13g2_Filler200 IO_FILL_IO_WEST_2_3 ();
 sg13g2_Filler200 IO_FILL_IO_WEST_2_4 ();
 sg13g2_Filler200 IO_FILL_IO_WEST_2_5 ();
 sg13g2_Filler200 IO_FILL_IO_WEST_2_6 ();
 sg13g2_Filler200 IO_FILL_IO_WEST_2_7 ();
 sg13g2_Filler200 IO_FILL_IO_WEST_2_8 ();
 sg13g2_Filler200 IO_FILL_IO_WEST_2_9 ();
 sg13g2_Filler200 IO_FILL_IO_WEST_3_0 ();
 sg13g2_Filler200 IO_FILL_IO_WEST_3_1 ();
 sg13g2_Filler200 IO_FILL_IO_WEST_3_2 ();
 sg13g2_Filler200 IO_FILL_IO_WEST_3_3 ();
 sg13g2_Filler200 IO_FILL_IO_WEST_3_4 ();
 sg13g2_Filler200 IO_FILL_IO_WEST_3_5 ();
 sg13g2_Filler200 IO_FILL_IO_WEST_3_6 ();
 sg13g2_Filler200 IO_FILL_IO_WEST_3_7 ();
 sg13g2_Filler200 IO_FILL_IO_WEST_3_8 ();
 sg13g2_Filler200 IO_FILL_IO_WEST_3_9 ();
 sg13g2_Filler200 IO_FILL_IO_WEST_4_0 ();
 sg13g2_Filler200 IO_FILL_IO_WEST_4_1 ();
 sg13g2_Filler200 IO_FILL_IO_WEST_4_2 ();
 sg13g2_Filler200 IO_FILL_IO_WEST_4_3 ();
 sg13g2_Filler200 IO_FILL_IO_WEST_4_4 ();
 sg13g2_Filler200 IO_FILL_IO_WEST_4_5 ();
 sg13g2_Filler200 IO_FILL_IO_WEST_4_6 ();
 sg13g2_Filler200 IO_FILL_IO_WEST_4_7 ();
 sg13g2_Filler200 IO_FILL_IO_WEST_4_8 ();
 sg13g2_Filler200 IO_FILL_IO_WEST_4_9 ();
 sg13g2_Filler200 IO_FILL_IO_WEST_5_0 ();
 sg13g2_Filler200 IO_FILL_IO_WEST_5_1 ();
 sg13g2_Filler200 IO_FILL_IO_WEST_5_2 ();
 sg13g2_Filler200 IO_FILL_IO_WEST_5_3 ();
 sg13g2_Filler200 IO_FILL_IO_WEST_5_4 ();
 sg13g2_Filler200 IO_FILL_IO_WEST_5_5 ();
 sg13g2_Filler200 IO_FILL_IO_WEST_5_6 ();
 sg13g2_Filler200 IO_FILL_IO_WEST_5_7 ();
 sg13g2_Filler200 IO_FILL_IO_WEST_5_8 ();
 sg13g2_Filler200 IO_FILL_IO_WEST_5_9 ();
 sg13g2_Filler200 IO_FILL_IO_WEST_6_0 ();
 sg13g2_Filler200 IO_FILL_IO_WEST_6_1 ();
 sg13g2_Filler200 IO_FILL_IO_WEST_6_2 ();
 sg13g2_Filler200 IO_FILL_IO_WEST_6_3 ();
 sg13g2_Filler200 IO_FILL_IO_WEST_6_4 ();
 sg13g2_Filler200 IO_FILL_IO_WEST_6_5 ();
 sg13g2_Filler200 IO_FILL_IO_WEST_6_6 ();
 sg13g2_Filler200 IO_FILL_IO_WEST_6_7 ();
 sg13g2_Filler200 IO_FILL_IO_WEST_6_8 ();
 sg13g2_Filler200 IO_FILL_IO_WEST_6_9 ();
 sg13g2_Filler200 IO_FILL_IO_WEST_7_0 ();
 sg13g2_Filler200 IO_FILL_IO_WEST_7_1 ();
 sg13g2_Filler200 IO_FILL_IO_WEST_7_2 ();
 sg13g2_Filler200 IO_FILL_IO_WEST_7_3 ();
 sg13g2_Filler200 IO_FILL_IO_WEST_7_4 ();
 sg13g2_Filler200 IO_FILL_IO_WEST_7_5 ();
 sg13g2_Filler200 IO_FILL_IO_WEST_7_6 ();
 sg13g2_Filler200 IO_FILL_IO_WEST_7_7 ();
 sg13g2_Filler200 IO_FILL_IO_WEST_7_8 ();
 sg13g2_Filler200 IO_FILL_IO_WEST_7_9 ();
 sg13g2_Filler200 IO_FILL_IO_WEST_8_0 ();
 sg13g2_Filler200 IO_FILL_IO_WEST_8_1 ();
 sg13g2_Filler200 IO_FILL_IO_WEST_8_2 ();
 sg13g2_Filler200 IO_FILL_IO_WEST_8_3 ();
 sg13g2_Filler200 IO_FILL_IO_WEST_8_4 ();
 sg13g2_Filler200 IO_FILL_IO_WEST_8_5 ();
 sg13g2_Filler200 IO_FILL_IO_WEST_8_6 ();
 sg13g2_Filler200 IO_FILL_IO_WEST_8_7 ();
 sg13g2_Filler200 IO_FILL_IO_WEST_8_8 ();
 sg13g2_Filler200 IO_FILL_IO_WEST_8_9 ();
 sg13g2_Filler200 IO_FILL_IO_EAST_0_0 ();
 sg13g2_Filler200 IO_FILL_IO_EAST_0_1 ();
 sg13g2_Filler200 IO_FILL_IO_EAST_0_2 ();
 sg13g2_Filler200 IO_FILL_IO_EAST_0_3 ();
 sg13g2_Filler200 IO_FILL_IO_EAST_0_4 ();
 sg13g2_Filler200 IO_FILL_IO_EAST_0_5 ();
 sg13g2_Filler200 IO_FILL_IO_EAST_0_6 ();
 sg13g2_Filler200 IO_FILL_IO_EAST_0_7 ();
 sg13g2_Filler200 IO_FILL_IO_EAST_0_8 ();
 sg13g2_Filler200 IO_FILL_IO_EAST_0_9 ();
 sg13g2_Filler200 IO_FILL_IO_EAST_1_0 ();
 sg13g2_Filler200 IO_FILL_IO_EAST_1_1 ();
 sg13g2_Filler200 IO_FILL_IO_EAST_1_2 ();
 sg13g2_Filler200 IO_FILL_IO_EAST_1_3 ();
 sg13g2_Filler200 IO_FILL_IO_EAST_1_4 ();
 sg13g2_Filler200 IO_FILL_IO_EAST_1_5 ();
 sg13g2_Filler200 IO_FILL_IO_EAST_1_6 ();
 sg13g2_Filler200 IO_FILL_IO_EAST_1_7 ();
 sg13g2_Filler200 IO_FILL_IO_EAST_1_8 ();
 sg13g2_Filler200 IO_FILL_IO_EAST_1_9 ();
 sg13g2_Filler200 IO_FILL_IO_EAST_2_0 ();
 sg13g2_Filler200 IO_FILL_IO_EAST_2_1 ();
 sg13g2_Filler200 IO_FILL_IO_EAST_2_2 ();
 sg13g2_Filler200 IO_FILL_IO_EAST_2_3 ();
 sg13g2_Filler200 IO_FILL_IO_EAST_2_4 ();
 sg13g2_Filler200 IO_FILL_IO_EAST_2_5 ();
 sg13g2_Filler200 IO_FILL_IO_EAST_2_6 ();
 sg13g2_Filler200 IO_FILL_IO_EAST_2_7 ();
 sg13g2_Filler200 IO_FILL_IO_EAST_2_8 ();
 sg13g2_Filler200 IO_FILL_IO_EAST_2_9 ();
 sg13g2_Filler200 IO_FILL_IO_EAST_3_0 ();
 sg13g2_Filler200 IO_FILL_IO_EAST_3_1 ();
 sg13g2_Filler200 IO_FILL_IO_EAST_3_2 ();
 sg13g2_Filler200 IO_FILL_IO_EAST_3_3 ();
 sg13g2_Filler200 IO_FILL_IO_EAST_3_4 ();
 sg13g2_Filler200 IO_FILL_IO_EAST_3_5 ();
 sg13g2_Filler200 IO_FILL_IO_EAST_3_6 ();
 sg13g2_Filler200 IO_FILL_IO_EAST_3_7 ();
 sg13g2_Filler200 IO_FILL_IO_EAST_3_8 ();
 sg13g2_Filler200 IO_FILL_IO_EAST_3_9 ();
 sg13g2_Filler200 IO_FILL_IO_EAST_4_0 ();
 sg13g2_Filler200 IO_FILL_IO_EAST_4_1 ();
 sg13g2_Filler200 IO_FILL_IO_EAST_4_2 ();
 sg13g2_Filler200 IO_FILL_IO_EAST_4_3 ();
 sg13g2_Filler200 IO_FILL_IO_EAST_4_4 ();
 sg13g2_Filler200 IO_FILL_IO_EAST_4_5 ();
 sg13g2_Filler200 IO_FILL_IO_EAST_4_6 ();
 sg13g2_Filler200 IO_FILL_IO_EAST_4_7 ();
 sg13g2_Filler200 IO_FILL_IO_EAST_4_8 ();
 sg13g2_Filler200 IO_FILL_IO_EAST_4_9 ();
 sg13g2_Filler200 IO_FILL_IO_EAST_5_0 ();
 sg13g2_Filler200 IO_FILL_IO_EAST_5_1 ();
 sg13g2_Filler200 IO_FILL_IO_EAST_5_2 ();
 sg13g2_Filler200 IO_FILL_IO_EAST_5_3 ();
 sg13g2_Filler200 IO_FILL_IO_EAST_5_4 ();
 sg13g2_Filler200 IO_FILL_IO_EAST_5_5 ();
 sg13g2_Filler200 IO_FILL_IO_EAST_5_6 ();
 sg13g2_Filler200 IO_FILL_IO_EAST_5_7 ();
 sg13g2_Filler200 IO_FILL_IO_EAST_5_8 ();
 sg13g2_Filler200 IO_FILL_IO_EAST_5_9 ();
 sg13g2_Filler200 IO_FILL_IO_EAST_6_0 ();
 sg13g2_Filler200 IO_FILL_IO_EAST_6_1 ();
 sg13g2_Filler200 IO_FILL_IO_EAST_6_2 ();
 sg13g2_Filler200 IO_FILL_IO_EAST_6_3 ();
 sg13g2_Filler200 IO_FILL_IO_EAST_6_4 ();
 sg13g2_Filler200 IO_FILL_IO_EAST_6_5 ();
 sg13g2_Filler200 IO_FILL_IO_EAST_6_6 ();
 sg13g2_Filler200 IO_FILL_IO_EAST_6_7 ();
 sg13g2_Filler200 IO_FILL_IO_EAST_6_8 ();
 sg13g2_Filler200 IO_FILL_IO_EAST_6_9 ();
 sg13g2_Filler200 IO_FILL_IO_EAST_7_0 ();
 sg13g2_Filler200 IO_FILL_IO_EAST_7_1 ();
 sg13g2_Filler200 IO_FILL_IO_EAST_7_2 ();
 sg13g2_Filler200 IO_FILL_IO_EAST_7_3 ();
 sg13g2_Filler200 IO_FILL_IO_EAST_7_4 ();
 sg13g2_Filler200 IO_FILL_IO_EAST_7_5 ();
 sg13g2_Filler200 IO_FILL_IO_EAST_7_6 ();
 sg13g2_Filler200 IO_FILL_IO_EAST_7_7 ();
 sg13g2_Filler200 IO_FILL_IO_EAST_7_8 ();
 sg13g2_Filler200 IO_FILL_IO_EAST_7_9 ();
 sg13g2_Filler200 IO_FILL_IO_EAST_8_0 ();
 sg13g2_Filler200 IO_FILL_IO_EAST_8_1 ();
 sg13g2_Filler200 IO_FILL_IO_EAST_8_2 ();
 sg13g2_Filler200 IO_FILL_IO_EAST_8_3 ();
 sg13g2_Filler200 IO_FILL_IO_EAST_8_4 ();
 sg13g2_Filler200 IO_FILL_IO_EAST_8_5 ();
 sg13g2_Filler200 IO_FILL_IO_EAST_8_6 ();
 sg13g2_Filler200 IO_FILL_IO_EAST_8_7 ();
 sg13g2_Filler200 IO_FILL_IO_EAST_8_8 ();
 sg13g2_Filler200 IO_FILL_IO_EAST_8_9 ();
 bondpad_70x70 IO_BOND_port_aux_enable_cell (.pad(aux_enable_pad));
 bondpad_70x70 IO_BOND_port_clk_cell (.pad(clk_pad));
 bondpad_70x70 IO_BOND_port_data_in1_cell (.pad(data_in_pad[0]));
 bondpad_70x70 IO_BOND_port_data_in2_cell (.pad(data_in_pad[1]));
 bondpad_70x70 IO_BOND_port_data_in3_cell (.pad(data_in_pad[2]));
 bondpad_70x70 IO_BOND_port_data_in4_cell (.pad(data_in_pad[3]));
 bondpad_70x70 IO_BOND_port_data_in5_cell (.pad(data_in_pad[4]));
 bondpad_70x70 IO_BOND_port_data_in6_cell (.pad(data_in_pad[5]));
 bondpad_70x70 IO_BOND_port_data_in7_cell (.pad(data_in_pad[6]));
 bondpad_70x70 IO_BOND_port_data_in8_cell (.pad(data_in_pad[7]));
 bondpad_70x70 IO_BOND_port_data_out1_cell (.pad(data_out_pad[0]));
 bondpad_70x70 IO_BOND_port_data_out2_cell (.pad(data_out_pad[1]));
 bondpad_70x70 IO_BOND_port_data_out3_cell (.pad(data_out_pad[2]));
 bondpad_70x70 IO_BOND_port_data_out4_cell (.pad(data_out_pad[3]));
 bondpad_70x70 IO_BOND_port_data_out5_cell (.pad(data_out_pad[4]));
 bondpad_70x70 IO_BOND_port_data_out6_cell (.pad(data_out_pad[5]));
 bondpad_70x70 IO_BOND_port_data_out7_cell (.pad(data_out_pad[6]));
 bondpad_70x70 IO_BOND_port_data_out8_cell (.pad(data_out_pad[7]));
 bondpad_70x70 IO_BOND_port_lfsr_out_cell (.pad(lfsr_out_pad));
 bondpad_70x70 IO_BOND_port_out_select1_cell (.pad(out_select_pad[0]));
 bondpad_70x70 IO_BOND_port_out_select2_cell (.pad(out_select_pad[1]));
 bondpad_70x70 IO_BOND_port_reg_addr1_cell (.pad(reg_addr_pad[0]));
 bondpad_70x70 IO_BOND_port_reg_addr2_cell (.pad(reg_addr_pad[1]));
 bondpad_70x70 IO_BOND_port_reg_addr3_cell (.pad(reg_addr_pad[2]));
 bondpad_70x70 IO_BOND_port_rst_cell (.pad(rst_pad));
 bondpad_70x70 IO_BOND_port_shreg_in_cell (.pad(shreg_in_pad));
 bondpad_70x70 IO_BOND_port_shreg_out_cell (.pad(shreg_out_pad));
 bondpad_70x70 IO_BOND_port_wr_enable_cell (.pad(wr_enable_pad));
 bondpad_70x70 IO_BOND_VSS (.pad(\IO_CORNER_NORTH_WEST_INST.vss_RING ));
 bondpad_70x70 IO_BOND_VDD (.pad(\IO_CORNER_NORTH_WEST_INST.vdd_RING ));
 bondpad_70x70 IO_BOND_IOVDD (.pad(\IO_CORNER_NORTH_WEST_INST.iovdd_RING ));
 bondpad_70x70 IO_BOND_IOVSS (.pad(\IO_CORNER_NORTH_WEST_INST.iovss_RING ));
 sg13g2_buf_2 fanout1 (.A(_02815_),
    .X(net1));
 sg13g2_buf_2 fanout2 (.A(_02546_),
    .X(net2));
 sg13g2_buf_8 wire3 (.A(net3),
    .X(data_out_c2p[7]));
 sg13g2_buf_2 fanout4 (.A(_02545_),
    .X(net4));
 sg13g2_buf_2 fanout5 (.A(_02829_),
    .X(net5));
 sg13g2_buf_2 fanout6 (.A(_02820_),
    .X(net6));
 sg13g2_buf_2 fanout7 (.A(_02016_),
    .X(net7));
 sg13g2_buf_8 wire8 (.A(net8),
    .X(data_out_c2p[6]));
 sg13g2_buf_2 fanout9 (.A(_02825_),
    .X(net9));
 sg13g2_buf_2 fanout10 (.A(_02718_),
    .X(net10));
 sg13g2_buf_8 wire11 (.A(net11),
    .X(data_out_c2p[5]));
 sg13g2_buf_8 wire12 (.A(net12),
    .X(data_out_c2p[4]));
 sg13g2_buf_8 wire13 (.A(net13),
    .X(data_out_c2p[3]));
 sg13g2_buf_2 fanout14 (.A(_02048_),
    .X(net14));
 sg13g2_buf_2 fanout15 (.A(_02671_),
    .X(net15));
 sg13g2_buf_2 fanout16 (.A(_02370_),
    .X(net16));
 sg13g2_buf_2 fanout17 (.A(_02289_),
    .X(net17));
 sg13g2_buf_2 fanout18 (.A(_02754_),
    .X(net18));
 sg13g2_buf_2 fanout19 (.A(_02628_),
    .X(net19));
 sg13g2_buf_2 fanout20 (.A(_02464_),
    .X(net20));
 sg13g2_buf_2 fanout21 (.A(_02394_),
    .X(net21));
 sg13g2_buf_2 fanout22 (.A(_02226_),
    .X(net22));
 sg13g2_buf_2 fanout23 (.A(_02166_),
    .X(net23));
 sg13g2_buf_2 fanout24 (.A(_01896_),
    .X(net24));
 sg13g2_buf_2 fanout25 (.A(_01852_),
    .X(net25));
 sg13g2_buf_2 fanout26 (.A(_02201_),
    .X(net26));
 sg13g2_buf_8 wire27 (.A(net27),
    .X(data_out_c2p[2]));
 sg13g2_buf_2 fanout28 (.A(_01805_),
    .X(net28));
 sg13g2_buf_8 wire29 (.A(net29),
    .X(data_out_c2p[1]));
 sg13g2_buf_2 fanout30 (.A(_03065_),
    .X(net30));
 sg13g2_buf_2 fanout31 (.A(_03064_),
    .X(net31));
 sg13g2_buf_2 fanout32 (.A(_03062_),
    .X(net32));
 sg13g2_buf_1 fanout33 (.A(_04267_),
    .X(net33));
 sg13g2_buf_2 fanout34 (.A(_04255_),
    .X(net34));
 sg13g2_buf_1 fanout35 (.A(_04243_),
    .X(net35));
 sg13g2_buf_1 fanout36 (.A(_04231_),
    .X(net36));
 sg13g2_buf_1 fanout37 (.A(_04219_),
    .X(net37));
 sg13g2_buf_1 fanout38 (.A(_04207_),
    .X(net38));
 sg13g2_buf_1 fanout39 (.A(_04195_),
    .X(net39));
 sg13g2_buf_1 fanout40 (.A(_04183_),
    .X(net40));
 sg13g2_buf_1 fanout41 (.A(_04171_),
    .X(net41));
 sg13g2_buf_1 fanout42 (.A(_04159_),
    .X(net42));
 sg13g2_buf_1 fanout43 (.A(_04145_),
    .X(net43));
 sg13g2_buf_4 fanout44 (.X(net44),
    .A(_04138_));
 sg13g2_buf_1 fanout45 (.A(_04133_),
    .X(net45));
 sg13g2_buf_4 fanout46 (.X(net46),
    .A(_04126_));
 sg13g2_buf_2 fanout47 (.A(_04121_),
    .X(net47));
 sg13g2_buf_4 fanout48 (.X(net48),
    .A(_04114_));
 sg13g2_buf_1 fanout49 (.A(_04109_),
    .X(net49));
 sg13g2_buf_4 fanout50 (.X(net50),
    .A(_04102_));
 sg13g2_buf_1 fanout51 (.A(_04097_),
    .X(net51));
 sg13g2_buf_4 fanout52 (.X(net52),
    .A(_04090_));
 sg13g2_buf_1 fanout53 (.A(_04085_),
    .X(net53));
 sg13g2_buf_4 fanout54 (.X(net54),
    .A(_04078_));
 sg13g2_buf_1 fanout55 (.A(_04073_),
    .X(net55));
 sg13g2_buf_4 fanout56 (.X(net56),
    .A(_04066_));
 sg13g2_buf_1 fanout57 (.A(_04061_),
    .X(net57));
 sg13g2_buf_4 fanout58 (.X(net58),
    .A(_04054_));
 sg13g2_buf_2 fanout59 (.A(_04049_),
    .X(net59));
 sg13g2_buf_4 fanout60 (.X(net60),
    .A(_04042_));
 sg13g2_buf_1 fanout61 (.A(_04037_),
    .X(net61));
 sg13g2_buf_4 fanout62 (.X(net62),
    .A(_04029_));
 sg13g2_buf_1 fanout63 (.A(_04023_),
    .X(net63));
 sg13g2_buf_4 fanout64 (.X(net64),
    .A(_04016_));
 sg13g2_buf_1 fanout65 (.A(_04011_),
    .X(net65));
 sg13g2_buf_4 fanout66 (.X(net66),
    .A(_04004_));
 sg13g2_buf_1 fanout67 (.A(_03999_),
    .X(net67));
 sg13g2_buf_4 fanout68 (.X(net68),
    .A(_03992_));
 sg13g2_buf_1 fanout69 (.A(_03987_),
    .X(net69));
 sg13g2_buf_4 fanout70 (.X(net70),
    .A(_03980_));
 sg13g2_buf_1 fanout71 (.A(_03975_),
    .X(net71));
 sg13g2_buf_4 fanout72 (.X(net72),
    .A(_03968_));
 sg13g2_buf_1 fanout73 (.A(_03963_),
    .X(net73));
 sg13g2_buf_4 fanout74 (.X(net74),
    .A(_03956_));
 sg13g2_buf_1 fanout75 (.A(_03951_),
    .X(net75));
 sg13g2_buf_4 fanout76 (.X(net76),
    .A(_03944_));
 sg13g2_buf_2 fanout77 (.A(_03939_),
    .X(net77));
 sg13g2_buf_4 fanout78 (.X(net78),
    .A(_03932_));
 sg13g2_buf_1 fanout79 (.A(_03927_),
    .X(net79));
 sg13g2_buf_4 fanout80 (.X(net80),
    .A(_03920_));
 sg13g2_buf_1 fanout81 (.A(_03915_),
    .X(net81));
 sg13g2_buf_4 fanout82 (.X(net82),
    .A(_03907_));
 sg13g2_buf_2 fanout83 (.A(_03901_),
    .X(net83));
 sg13g2_buf_4 fanout84 (.X(net84),
    .A(_03894_));
 sg13g2_buf_2 fanout85 (.A(_03889_),
    .X(net85));
 sg13g2_buf_4 fanout86 (.X(net86),
    .A(_03882_));
 sg13g2_buf_1 fanout87 (.A(_03877_),
    .X(net87));
 sg13g2_buf_4 fanout88 (.X(net88),
    .A(_03870_));
 sg13g2_buf_1 fanout89 (.A(_03865_),
    .X(net89));
 sg13g2_buf_4 fanout90 (.X(net90),
    .A(_03858_));
 sg13g2_buf_1 fanout91 (.A(_03853_),
    .X(net91));
 sg13g2_buf_4 fanout92 (.X(net92),
    .A(_03846_));
 sg13g2_buf_1 fanout93 (.A(_03841_),
    .X(net93));
 sg13g2_buf_4 fanout94 (.X(net94),
    .A(_03834_));
 sg13g2_buf_1 fanout95 (.A(_03829_),
    .X(net95));
 sg13g2_buf_4 fanout96 (.X(net96),
    .A(_03822_));
 sg13g2_buf_1 fanout97 (.A(_03817_),
    .X(net97));
 sg13g2_buf_4 fanout98 (.X(net98),
    .A(_03810_));
 sg13g2_buf_1 fanout99 (.A(_03805_),
    .X(net99));
 sg13g2_buf_4 fanout100 (.X(net100),
    .A(_03798_));
 sg13g2_buf_1 fanout101 (.A(_03793_),
    .X(net101));
 sg13g2_buf_4 fanout102 (.X(net102),
    .A(_03785_));
 sg13g2_buf_1 fanout103 (.A(_03779_),
    .X(net103));
 sg13g2_buf_4 fanout104 (.X(net104),
    .A(_03772_));
 sg13g2_buf_2 fanout105 (.A(_03767_),
    .X(net105));
 sg13g2_buf_4 fanout106 (.X(net106),
    .A(_03760_));
 sg13g2_buf_1 fanout107 (.A(_03755_),
    .X(net107));
 sg13g2_buf_4 fanout108 (.X(net108),
    .A(_03748_));
 sg13g2_buf_1 fanout109 (.A(_03743_),
    .X(net109));
 sg13g2_buf_4 fanout110 (.X(net110),
    .A(_03736_));
 sg13g2_buf_1 fanout111 (.A(_03731_),
    .X(net111));
 sg13g2_buf_4 fanout112 (.X(net112),
    .A(_03724_));
 sg13g2_buf_1 fanout113 (.A(_03719_),
    .X(net113));
 sg13g2_buf_4 fanout114 (.X(net114),
    .A(_03712_));
 sg13g2_buf_1 fanout115 (.A(_03707_),
    .X(net115));
 sg13g2_buf_4 fanout116 (.X(net116),
    .A(_03700_));
 sg13g2_buf_1 fanout117 (.A(_03695_),
    .X(net117));
 sg13g2_buf_4 fanout118 (.X(net118),
    .A(_03688_));
 sg13g2_buf_1 fanout119 (.A(_03683_),
    .X(net119));
 sg13g2_buf_4 fanout120 (.X(net120),
    .A(_03676_));
 sg13g2_buf_1 fanout121 (.A(_03671_),
    .X(net121));
 sg13g2_buf_4 fanout122 (.X(net122),
    .A(_03663_));
 sg13g2_buf_1 fanout123 (.A(_03657_),
    .X(net123));
 sg13g2_buf_4 fanout124 (.X(net124),
    .A(_03650_));
 sg13g2_buf_2 fanout125 (.A(_03645_),
    .X(net125));
 sg13g2_buf_4 fanout126 (.X(net126),
    .A(_03638_));
 sg13g2_buf_1 fanout127 (.A(_03633_),
    .X(net127));
 sg13g2_buf_4 fanout128 (.X(net128),
    .A(_03626_));
 sg13g2_buf_1 fanout129 (.A(_03621_),
    .X(net129));
 sg13g2_buf_4 fanout130 (.X(net130),
    .A(_03614_));
 sg13g2_buf_1 fanout131 (.A(_03609_),
    .X(net131));
 sg13g2_buf_4 fanout132 (.X(net132),
    .A(_03602_));
 sg13g2_buf_1 fanout133 (.A(_03597_),
    .X(net133));
 sg13g2_buf_4 fanout134 (.X(net134),
    .A(_03590_));
 sg13g2_buf_1 fanout135 (.A(_03585_),
    .X(net135));
 sg13g2_buf_4 fanout136 (.X(net136),
    .A(_03578_));
 sg13g2_buf_1 fanout137 (.A(_03573_),
    .X(net137));
 sg13g2_buf_4 fanout138 (.X(net138),
    .A(_03566_));
 sg13g2_buf_1 fanout139 (.A(_03561_),
    .X(net139));
 sg13g2_buf_4 fanout140 (.X(net140),
    .A(_03554_));
 sg13g2_buf_1 fanout141 (.A(_03549_),
    .X(net141));
 sg13g2_buf_4 fanout142 (.X(net142),
    .A(_03541_));
 sg13g2_buf_1 fanout143 (.A(_03535_),
    .X(net143));
 sg13g2_buf_4 fanout144 (.X(net144),
    .A(_03528_));
 sg13g2_buf_2 fanout145 (.A(_03523_),
    .X(net145));
 sg13g2_buf_4 fanout146 (.X(net146),
    .A(_03516_));
 sg13g2_buf_1 fanout147 (.A(_03511_),
    .X(net147));
 sg13g2_buf_4 fanout148 (.X(net148),
    .A(_03504_));
 sg13g2_buf_1 fanout149 (.A(_03499_),
    .X(net149));
 sg13g2_buf_4 fanout150 (.X(net150),
    .A(_03492_));
 sg13g2_buf_1 fanout151 (.A(_03487_),
    .X(net151));
 sg13g2_buf_4 fanout152 (.X(net152),
    .A(_03480_));
 sg13g2_buf_1 fanout153 (.A(_03475_),
    .X(net153));
 sg13g2_buf_4 fanout154 (.X(net154),
    .A(_03468_));
 sg13g2_buf_2 fanout155 (.A(_03463_),
    .X(net155));
 sg13g2_buf_4 fanout156 (.X(net156),
    .A(_03456_));
 sg13g2_buf_1 fanout157 (.A(_03451_),
    .X(net157));
 sg13g2_buf_4 fanout158 (.X(net158),
    .A(_03444_));
 sg13g2_buf_2 fanout159 (.A(_03439_),
    .X(net159));
 sg13g2_buf_4 fanout160 (.X(net160),
    .A(_03432_));
 sg13g2_buf_1 fanout161 (.A(_03427_),
    .X(net161));
 sg13g2_buf_4 fanout162 (.X(net162),
    .A(_03419_));
 sg13g2_buf_1 fanout163 (.A(_03413_),
    .X(net163));
 sg13g2_buf_4 fanout164 (.X(net164),
    .A(_03406_));
 sg13g2_buf_2 fanout165 (.A(_03401_),
    .X(net165));
 sg13g2_buf_4 fanout166 (.X(net166),
    .A(_03394_));
 sg13g2_buf_2 fanout167 (.A(_03389_),
    .X(net167));
 sg13g2_buf_4 fanout168 (.X(net168),
    .A(_03382_));
 sg13g2_buf_1 fanout169 (.A(_03377_),
    .X(net169));
 sg13g2_buf_4 fanout170 (.X(net170),
    .A(_03370_));
 sg13g2_buf_1 fanout171 (.A(_03365_),
    .X(net171));
 sg13g2_buf_4 fanout172 (.X(net172),
    .A(_03358_));
 sg13g2_buf_1 fanout173 (.A(_03353_),
    .X(net173));
 sg13g2_buf_4 fanout174 (.X(net174),
    .A(_03346_));
 sg13g2_buf_1 fanout175 (.A(_03341_),
    .X(net175));
 sg13g2_buf_4 fanout176 (.X(net176),
    .A(_03334_));
 sg13g2_buf_2 fanout177 (.A(_03329_),
    .X(net177));
 sg13g2_buf_4 fanout178 (.X(net178),
    .A(_03322_));
 sg13g2_buf_1 fanout179 (.A(_03317_),
    .X(net179));
 sg13g2_buf_4 fanout180 (.X(net180),
    .A(_03310_));
 sg13g2_buf_2 fanout181 (.A(_03305_),
    .X(net181));
 sg13g2_buf_4 fanout182 (.X(net182),
    .A(_03297_));
 sg13g2_buf_1 fanout183 (.A(_03291_),
    .X(net183));
 sg13g2_buf_4 fanout184 (.X(net184),
    .A(_03284_));
 sg13g2_buf_1 fanout185 (.A(_03279_),
    .X(net185));
 sg13g2_buf_4 fanout186 (.X(net186),
    .A(_03272_));
 sg13g2_buf_1 fanout187 (.A(_03267_),
    .X(net187));
 sg13g2_buf_4 fanout188 (.X(net188),
    .A(_03260_));
 sg13g2_buf_1 fanout189 (.A(_03255_),
    .X(net189));
 sg13g2_buf_4 fanout190 (.X(net190),
    .A(_03248_));
 sg13g2_buf_1 fanout191 (.A(_03243_),
    .X(net191));
 sg13g2_buf_4 fanout192 (.X(net192),
    .A(_03236_));
 sg13g2_buf_1 fanout193 (.A(_03231_),
    .X(net193));
 sg13g2_buf_4 fanout194 (.X(net194),
    .A(_03224_));
 sg13g2_buf_1 fanout195 (.A(_03219_),
    .X(net195));
 sg13g2_buf_4 fanout196 (.X(net196),
    .A(_03212_));
 sg13g2_buf_2 fanout197 (.A(_03207_),
    .X(net197));
 sg13g2_buf_4 fanout198 (.X(net198),
    .A(_03200_));
 sg13g2_buf_1 fanout199 (.A(_03195_),
    .X(net199));
 sg13g2_buf_4 fanout200 (.X(net200),
    .A(_03188_));
 sg13g2_buf_1 fanout201 (.A(_03183_),
    .X(net201));
 sg13g2_buf_4 fanout202 (.X(net202),
    .A(_03175_));
 sg13g2_buf_2 fanout203 (.A(_03169_),
    .X(net203));
 sg13g2_buf_4 fanout204 (.X(net204),
    .A(_03162_));
 sg13g2_buf_2 fanout205 (.A(_03157_),
    .X(net205));
 sg13g2_buf_4 fanout206 (.X(net206),
    .A(_03150_));
 sg13g2_buf_1 fanout207 (.A(_03145_),
    .X(net207));
 sg13g2_buf_4 fanout208 (.X(net208),
    .A(_03138_));
 sg13g2_buf_1 fanout209 (.A(_03133_),
    .X(net209));
 sg13g2_buf_4 fanout210 (.X(net210),
    .A(_03126_));
 sg13g2_buf_2 fanout211 (.A(_03121_),
    .X(net211));
 sg13g2_buf_4 fanout212 (.X(net212),
    .A(_03114_));
 sg13g2_buf_1 fanout213 (.A(_03109_),
    .X(net213));
 sg13g2_buf_4 fanout214 (.X(net214),
    .A(_03102_));
 sg13g2_buf_1 fanout215 (.A(_03097_),
    .X(net215));
 sg13g2_buf_4 fanout216 (.X(net216),
    .A(_03090_));
 sg13g2_buf_1 fanout217 (.A(_03085_),
    .X(net217));
 sg13g2_buf_4 fanout218 (.X(net218),
    .A(_03078_));
 sg13g2_buf_1 fanout219 (.A(_03073_),
    .X(net219));
 sg13g2_buf_4 fanout220 (.X(net220),
    .A(_03066_));
 sg13g2_buf_2 fanout221 (.A(_03052_),
    .X(net221));
 sg13g2_buf_2 fanout222 (.A(_01902_),
    .X(net222));
 sg13g2_buf_4 fanout223 (.X(net223),
    .A(_05004_));
 sg13g2_buf_1 fanout224 (.A(_04999_),
    .X(net224));
 sg13g2_buf_4 fanout225 (.X(net225),
    .A(_04992_));
 sg13g2_buf_2 fanout226 (.A(_04987_),
    .X(net226));
 sg13g2_buf_4 fanout227 (.X(net227),
    .A(_04980_));
 sg13g2_buf_1 fanout228 (.A(_04975_),
    .X(net228));
 sg13g2_buf_4 fanout229 (.X(net229),
    .A(_04968_));
 sg13g2_buf_1 fanout230 (.A(_04963_),
    .X(net230));
 sg13g2_buf_4 fanout231 (.X(net231),
    .A(_04956_));
 sg13g2_buf_1 fanout232 (.A(_04951_),
    .X(net232));
 sg13g2_buf_4 fanout233 (.X(net233),
    .A(_04944_));
 sg13g2_buf_1 fanout234 (.A(_04939_),
    .X(net234));
 sg13g2_buf_4 fanout235 (.X(net235),
    .A(_04932_));
 sg13g2_buf_1 fanout236 (.A(_04927_),
    .X(net236));
 sg13g2_buf_4 fanout237 (.X(net237),
    .A(_04920_));
 sg13g2_buf_1 fanout238 (.A(_04915_),
    .X(net238));
 sg13g2_buf_4 fanout239 (.X(net239),
    .A(_04908_));
 sg13g2_buf_1 fanout240 (.A(_04903_),
    .X(net240));
 sg13g2_buf_4 fanout241 (.X(net241),
    .A(_04896_));
 sg13g2_buf_1 fanout242 (.A(_04891_),
    .X(net242));
 sg13g2_buf_4 fanout243 (.X(net243),
    .A(_04883_));
 sg13g2_buf_1 fanout244 (.A(_04877_),
    .X(net244));
 sg13g2_buf_4 fanout245 (.X(net245),
    .A(_04870_));
 sg13g2_buf_2 fanout246 (.A(_04865_),
    .X(net246));
 sg13g2_buf_4 fanout247 (.X(net247),
    .A(_04858_));
 sg13g2_buf_1 fanout248 (.A(_04853_),
    .X(net248));
 sg13g2_buf_4 fanout249 (.X(net249),
    .A(_04846_));
 sg13g2_buf_1 fanout250 (.A(_04841_),
    .X(net250));
 sg13g2_buf_4 fanout251 (.X(net251),
    .A(_04834_));
 sg13g2_buf_1 fanout252 (.A(_04829_),
    .X(net252));
 sg13g2_buf_4 fanout253 (.X(net253),
    .A(_04822_));
 sg13g2_buf_1 fanout254 (.A(_04817_),
    .X(net254));
 sg13g2_buf_4 fanout255 (.X(net255),
    .A(_04810_));
 sg13g2_buf_1 fanout256 (.A(_04805_),
    .X(net256));
 sg13g2_buf_4 fanout257 (.X(net257),
    .A(_04798_));
 sg13g2_buf_1 fanout258 (.A(_04793_),
    .X(net258));
 sg13g2_buf_4 fanout259 (.X(net259),
    .A(_04786_));
 sg13g2_buf_1 fanout260 (.A(_04781_),
    .X(net260));
 sg13g2_buf_4 fanout261 (.X(net261),
    .A(_04774_));
 sg13g2_buf_1 fanout262 (.A(_04769_),
    .X(net262));
 sg13g2_buf_4 fanout263 (.X(net263),
    .A(_04761_));
 sg13g2_buf_1 fanout264 (.A(_04755_),
    .X(net264));
 sg13g2_buf_4 fanout265 (.X(net265),
    .A(_04748_));
 sg13g2_buf_1 fanout266 (.A(_04743_),
    .X(net266));
 sg13g2_buf_4 fanout267 (.X(net267),
    .A(_04736_));
 sg13g2_buf_1 fanout268 (.A(_04731_),
    .X(net268));
 sg13g2_buf_4 fanout269 (.X(net269),
    .A(_04724_));
 sg13g2_buf_1 fanout270 (.A(_04719_),
    .X(net270));
 sg13g2_buf_4 fanout271 (.X(net271),
    .A(_04712_));
 sg13g2_buf_1 fanout272 (.A(_04707_),
    .X(net272));
 sg13g2_buf_4 fanout273 (.X(net273),
    .A(_04700_));
 sg13g2_buf_1 fanout274 (.A(_04695_),
    .X(net274));
 sg13g2_buf_4 fanout275 (.X(net275),
    .A(_04688_));
 sg13g2_buf_1 fanout276 (.A(_04683_),
    .X(net276));
 sg13g2_buf_4 fanout277 (.X(net277),
    .A(_04676_));
 sg13g2_buf_1 fanout278 (.A(_04671_),
    .X(net278));
 sg13g2_buf_4 fanout279 (.X(net279),
    .A(_04664_));
 sg13g2_buf_1 fanout280 (.A(_04659_),
    .X(net280));
 sg13g2_buf_4 fanout281 (.X(net281),
    .A(_04652_));
 sg13g2_buf_1 fanout282 (.A(_04647_),
    .X(net282));
 sg13g2_buf_4 fanout283 (.X(net283),
    .A(_04639_));
 sg13g2_buf_1 fanout284 (.A(_04633_),
    .X(net284));
 sg13g2_buf_4 fanout285 (.X(net285),
    .A(_04626_));
 sg13g2_buf_1 fanout286 (.A(_04621_),
    .X(net286));
 sg13g2_buf_4 fanout287 (.X(net287),
    .A(_04614_));
 sg13g2_buf_1 fanout288 (.A(_04609_),
    .X(net288));
 sg13g2_buf_4 fanout289 (.X(net289),
    .A(_04602_));
 sg13g2_buf_1 fanout290 (.A(_04597_),
    .X(net290));
 sg13g2_buf_4 fanout291 (.X(net291),
    .A(_04590_));
 sg13g2_buf_1 fanout292 (.A(_04585_),
    .X(net292));
 sg13g2_buf_4 fanout293 (.X(net293),
    .A(_04578_));
 sg13g2_buf_1 fanout294 (.A(_04573_),
    .X(net294));
 sg13g2_buf_4 fanout295 (.X(net295),
    .A(_04566_));
 sg13g2_buf_1 fanout296 (.A(_04561_),
    .X(net296));
 sg13g2_buf_4 fanout297 (.X(net297),
    .A(_04554_));
 sg13g2_buf_1 fanout298 (.A(_04549_),
    .X(net298));
 sg13g2_buf_4 fanout299 (.X(net299),
    .A(_04542_));
 sg13g2_buf_1 fanout300 (.A(_04537_),
    .X(net300));
 sg13g2_buf_4 fanout301 (.X(net301),
    .A(_04530_));
 sg13g2_buf_1 fanout302 (.A(_04525_),
    .X(net302));
 sg13g2_buf_4 fanout303 (.X(net303),
    .A(_04517_));
 sg13g2_buf_1 fanout304 (.A(_04511_),
    .X(net304));
 sg13g2_buf_4 fanout305 (.X(net305),
    .A(_04504_));
 sg13g2_buf_1 fanout306 (.A(_04499_),
    .X(net306));
 sg13g2_buf_4 fanout307 (.X(net307),
    .A(_04492_));
 sg13g2_buf_1 fanout308 (.A(_04487_),
    .X(net308));
 sg13g2_buf_4 fanout309 (.X(net309),
    .A(_04480_));
 sg13g2_buf_1 fanout310 (.A(_04475_),
    .X(net310));
 sg13g2_buf_4 fanout311 (.X(net311),
    .A(_04468_));
 sg13g2_buf_1 fanout312 (.A(_04463_),
    .X(net312));
 sg13g2_buf_4 fanout313 (.X(net313),
    .A(_04456_));
 sg13g2_buf_1 fanout314 (.A(_04451_),
    .X(net314));
 sg13g2_buf_4 fanout315 (.X(net315),
    .A(_04444_));
 sg13g2_buf_1 fanout316 (.A(_04439_),
    .X(net316));
 sg13g2_buf_4 fanout317 (.X(net317),
    .A(_04432_));
 sg13g2_buf_2 fanout318 (.A(_04427_),
    .X(net318));
 sg13g2_buf_4 fanout319 (.X(net319),
    .A(_04420_));
 sg13g2_buf_1 fanout320 (.A(_04415_),
    .X(net320));
 sg13g2_buf_4 fanout321 (.X(net321),
    .A(_04408_));
 sg13g2_buf_1 fanout322 (.A(_04403_),
    .X(net322));
 sg13g2_buf_4 fanout323 (.X(net323),
    .A(_04395_));
 sg13g2_buf_2 fanout324 (.A(_04389_),
    .X(net324));
 sg13g2_buf_4 fanout325 (.X(net325),
    .A(_04382_));
 sg13g2_buf_1 fanout326 (.A(_04377_),
    .X(net326));
 sg13g2_buf_4 fanout327 (.X(net327),
    .A(_04370_));
 sg13g2_buf_1 fanout328 (.A(_04365_),
    .X(net328));
 sg13g2_buf_4 fanout329 (.X(net329),
    .A(_04358_));
 sg13g2_buf_1 fanout330 (.A(_04353_),
    .X(net330));
 sg13g2_buf_4 fanout331 (.X(net331),
    .A(_04346_));
 sg13g2_buf_1 fanout332 (.A(_04341_),
    .X(net332));
 sg13g2_buf_4 fanout333 (.X(net333),
    .A(_04334_));
 sg13g2_buf_1 fanout334 (.A(_04329_),
    .X(net334));
 sg13g2_buf_4 fanout335 (.X(net335),
    .A(_04322_));
 sg13g2_buf_1 fanout336 (.A(_04317_),
    .X(net336));
 sg13g2_buf_4 fanout337 (.X(net337),
    .A(_04310_));
 sg13g2_buf_1 fanout338 (.A(_04305_),
    .X(net338));
 sg13g2_buf_4 fanout339 (.X(net339),
    .A(_04298_));
 sg13g2_buf_2 fanout340 (.A(_04293_),
    .X(net340));
 sg13g2_buf_4 fanout341 (.X(net341),
    .A(_04286_));
 sg13g2_buf_1 fanout342 (.A(_04281_),
    .X(net342));
 sg13g2_buf_4 fanout343 (.X(net343),
    .A(_04273_));
 sg13g2_buf_4 fanout344 (.X(net344),
    .A(_04260_));
 sg13g2_buf_4 fanout345 (.X(net345),
    .A(_04248_));
 sg13g2_buf_4 fanout346 (.X(net346),
    .A(_04236_));
 sg13g2_buf_4 fanout347 (.X(net347),
    .A(_04224_));
 sg13g2_buf_4 fanout348 (.X(net348),
    .A(_04212_));
 sg13g2_buf_4 fanout349 (.X(net349),
    .A(_04200_));
 sg13g2_buf_4 fanout350 (.X(net350),
    .A(_04188_));
 sg13g2_buf_4 fanout351 (.X(net351),
    .A(_04176_));
 sg13g2_buf_4 fanout352 (.X(net352),
    .A(_04164_));
 sg13g2_buf_2 fanout353 (.A(_04158_),
    .X(net353));
 sg13g2_buf_4 fanout354 (.X(net354),
    .A(_04151_));
 sg13g2_buf_1 fanout355 (.A(_04036_),
    .X(net355));
 sg13g2_buf_1 fanout356 (.A(_04028_),
    .X(net356));
 sg13g2_buf_1 fanout357 (.A(_03914_),
    .X(net357));
 sg13g2_buf_2 fanout358 (.A(_03906_),
    .X(net358));
 sg13g2_buf_2 fanout359 (.A(_03792_),
    .X(net359));
 sg13g2_buf_2 fanout360 (.A(_03784_),
    .X(net360));
 sg13g2_buf_1 fanout361 (.A(_03670_),
    .X(net361));
 sg13g2_buf_1 fanout362 (.A(_03662_),
    .X(net362));
 sg13g2_buf_1 fanout363 (.A(_03548_),
    .X(net363));
 sg13g2_buf_2 fanout364 (.A(_03540_),
    .X(net364));
 sg13g2_buf_2 fanout365 (.A(_03426_),
    .X(net365));
 sg13g2_buf_2 fanout366 (.A(_03418_),
    .X(net366));
 sg13g2_buf_2 fanout367 (.A(_03304_),
    .X(net367));
 sg13g2_buf_2 fanout368 (.A(_03296_),
    .X(net368));
 sg13g2_buf_2 fanout369 (.A(_03182_),
    .X(net369));
 sg13g2_buf_1 fanout370 (.A(_03174_),
    .X(net370));
 sg13g2_buf_1 fanout371 (.A(_03060_),
    .X(net371));
 sg13g2_buf_1 fanout372 (.A(_03051_),
    .X(net372));
 sg13g2_buf_2 fanout373 (.A(_03038_),
    .X(net373));
 sg13g2_buf_2 fanout374 (.A(_03034_),
    .X(net374));
 sg13g2_buf_2 fanout375 (.A(_03018_),
    .X(net375));
 sg13g2_buf_2 fanout376 (.A(_03011_),
    .X(net376));
 sg13g2_buf_2 fanout377 (.A(_03000_),
    .X(net377));
 sg13g2_buf_2 fanout378 (.A(_02990_),
    .X(net378));
 sg13g2_buf_2 fanout379 (.A(_02979_),
    .X(net379));
 sg13g2_buf_1 fanout380 (.A(_02966_),
    .X(net380));
 sg13g2_buf_2 fanout381 (.A(_02957_),
    .X(net381));
 sg13g2_buf_2 fanout382 (.A(_02943_),
    .X(net382));
 sg13g2_buf_2 fanout383 (.A(_02936_),
    .X(net383));
 sg13g2_buf_2 fanout384 (.A(_02919_),
    .X(net384));
 sg13g2_buf_2 fanout385 (.A(_02916_),
    .X(net385));
 sg13g2_buf_2 fanout386 (.A(_02911_),
    .X(net386));
 sg13g2_buf_2 fanout387 (.A(_02306_),
    .X(net387));
 sg13g2_buf_2 fanout388 (.A(_02223_),
    .X(net388));
 sg13g2_buf_2 fanout389 (.A(_02035_),
    .X(net389));
 sg13g2_buf_2 fanout390 (.A(_02020_),
    .X(net390));
 sg13g2_buf_2 fanout391 (.A(_01944_),
    .X(net391));
 sg13g2_buf_2 fanout392 (.A(_01929_),
    .X(net392));
 sg13g2_buf_2 fanout393 (.A(_01848_),
    .X(net393));
 sg13g2_buf_2 fanout394 (.A(_01847_),
    .X(net394));
 sg13g2_buf_2 fanout395 (.A(_01833_),
    .X(net395));
 sg13g2_buf_2 fanout396 (.A(_01719_),
    .X(net396));
 sg13g2_buf_1 fanout397 (.A(_04890_),
    .X(net397));
 sg13g2_buf_1 fanout398 (.A(_04882_),
    .X(net398));
 sg13g2_buf_1 fanout399 (.A(_04768_),
    .X(net399));
 sg13g2_buf_1 fanout400 (.A(_04760_),
    .X(net400));
 sg13g2_buf_1 fanout401 (.A(_04646_),
    .X(net401));
 sg13g2_buf_1 fanout402 (.A(_04638_),
    .X(net402));
 sg13g2_buf_1 fanout403 (.A(_04524_),
    .X(net403));
 sg13g2_buf_1 fanout404 (.A(_04516_),
    .X(net404));
 sg13g2_buf_2 fanout405 (.A(_04402_),
    .X(net405));
 sg13g2_buf_1 fanout406 (.A(_04394_),
    .X(net406));
 sg13g2_buf_1 fanout407 (.A(_04280_),
    .X(net407));
 sg13g2_buf_2 fanout408 (.A(_04272_),
    .X(net408));
 sg13g2_buf_1 fanout409 (.A(_04150_),
    .X(net409));
 sg13g2_buf_2 fanout410 (.A(_03059_),
    .X(net410));
 sg13g2_buf_2 fanout411 (.A(_03050_),
    .X(net411));
 sg13g2_buf_2 fanout412 (.A(_02910_),
    .X(net412));
 sg13g2_buf_2 fanout413 (.A(_02422_),
    .X(net413));
 sg13g2_buf_2 fanout414 (.A(_02177_),
    .X(net414));
 sg13g2_buf_2 fanout415 (.A(_02168_),
    .X(net415));
 sg13g2_buf_2 fanout416 (.A(_02150_),
    .X(net416));
 sg13g2_buf_2 fanout417 (.A(_02141_),
    .X(net417));
 sg13g2_buf_2 fanout418 (.A(_02137_),
    .X(net418));
 sg13g2_buf_2 fanout419 (.A(_02133_),
    .X(net419));
 sg13g2_buf_2 fanout420 (.A(_02104_),
    .X(net420));
 sg13g2_buf_2 fanout421 (.A(_02072_),
    .X(net421));
 sg13g2_buf_2 fanout422 (.A(_02061_),
    .X(net422));
 sg13g2_buf_2 fanout423 (.A(_02059_),
    .X(net423));
 sg13g2_buf_2 fanout424 (.A(_02051_),
    .X(net424));
 sg13g2_buf_2 fanout425 (.A(_02050_),
    .X(net425));
 sg13g2_buf_2 fanout426 (.A(_02038_),
    .X(net426));
 sg13g2_buf_2 fanout427 (.A(_02034_),
    .X(net427));
 sg13g2_buf_2 fanout428 (.A(_02026_),
    .X(net428));
 sg13g2_buf_2 fanout429 (.A(_02023_),
    .X(net429));
 sg13g2_buf_2 fanout430 (.A(_02021_),
    .X(net430));
 sg13g2_buf_2 fanout431 (.A(_02019_),
    .X(net431));
 sg13g2_buf_2 fanout432 (.A(_02018_),
    .X(net432));
 sg13g2_buf_2 fanout433 (.A(_01984_),
    .X(net433));
 sg13g2_buf_2 fanout434 (.A(_01981_),
    .X(net434));
 sg13g2_buf_2 fanout435 (.A(_01978_),
    .X(net435));
 sg13g2_buf_2 fanout436 (.A(_01972_),
    .X(net436));
 sg13g2_buf_2 fanout437 (.A(_01968_),
    .X(net437));
 sg13g2_buf_2 fanout438 (.A(_01967_),
    .X(net438));
 sg13g2_buf_2 fanout439 (.A(_01962_),
    .X(net439));
 sg13g2_buf_2 fanout440 (.A(_01946_),
    .X(net440));
 sg13g2_buf_2 fanout441 (.A(_01912_),
    .X(net441));
 sg13g2_buf_2 fanout442 (.A(_01910_),
    .X(net442));
 sg13g2_buf_2 fanout443 (.A(_01904_),
    .X(net443));
 sg13g2_buf_2 fanout444 (.A(_01900_),
    .X(net444));
 sg13g2_buf_2 fanout445 (.A(_01897_),
    .X(net445));
 sg13g2_buf_2 fanout446 (.A(_01867_),
    .X(net446));
 sg13g2_buf_2 fanout447 (.A(_01863_),
    .X(net447));
 sg13g2_buf_2 fanout448 (.A(_01859_),
    .X(net448));
 sg13g2_buf_2 fanout449 (.A(_01857_),
    .X(net449));
 sg13g2_buf_2 fanout450 (.A(_01855_),
    .X(net450));
 sg13g2_buf_2 fanout451 (.A(_01853_),
    .X(net451));
 sg13g2_buf_2 fanout452 (.A(_01843_),
    .X(net452));
 sg13g2_buf_2 fanout453 (.A(_01834_),
    .X(net453));
 sg13g2_buf_2 fanout454 (.A(_01825_),
    .X(net454));
 sg13g2_buf_2 fanout455 (.A(_01823_),
    .X(net455));
 sg13g2_buf_2 fanout456 (.A(_01822_),
    .X(net456));
 sg13g2_buf_2 fanout457 (.A(_01818_),
    .X(net457));
 sg13g2_buf_2 fanout458 (.A(_01817_),
    .X(net458));
 sg13g2_buf_2 fanout459 (.A(_01815_),
    .X(net459));
 sg13g2_buf_2 fanout460 (.A(_01801_),
    .X(net460));
 sg13g2_buf_2 fanout461 (.A(_01752_),
    .X(net461));
 sg13g2_buf_2 fanout462 (.A(_01751_),
    .X(net462));
 sg13g2_buf_2 fanout463 (.A(_01738_),
    .X(net463));
 sg13g2_buf_2 fanout464 (.A(_01732_),
    .X(net464));
 sg13g2_buf_2 fanout465 (.A(_01731_),
    .X(net465));
 sg13g2_buf_2 fanout466 (.A(_01730_),
    .X(net466));
 sg13g2_buf_2 fanout467 (.A(_01725_),
    .X(net467));
 sg13g2_buf_2 fanout468 (.A(_01721_),
    .X(net468));
 sg13g2_buf_2 fanout469 (.A(_01707_),
    .X(net469));
 sg13g2_buf_2 fanout470 (.A(_01706_),
    .X(net470));
 sg13g2_buf_2 fanout471 (.A(_01703_),
    .X(net471));
 sg13g2_buf_2 fanout472 (.A(\median_processor.input_storage [7]),
    .X(net472));
 sg13g2_buf_2 fanout473 (.A(\median_processor.input_storage [63]),
    .X(net473));
 sg13g2_buf_2 fanout474 (.A(\median_processor.input_storage [49]),
    .X(net474));
 sg13g2_buf_2 fanout475 (.A(\median_processor.input_storage [41]),
    .X(net475));
 sg13g2_buf_2 fanout476 (.A(\median_processor.input_storage [37]),
    .X(net476));
 sg13g2_buf_2 fanout477 (.A(\median_processor.input_storage [32]),
    .X(net477));
 sg13g2_buf_2 fanout478 (.A(\median_processor.input_storage [2]),
    .X(net478));
 sg13g2_buf_2 fanout479 (.A(\median_processor.input_storage [25]),
    .X(net479));
 sg13g2_buf_2 fanout480 (.A(\median_processor.input_storage [21]),
    .X(net480));
 sg13g2_buf_2 fanout481 (.A(\median_processor.input_storage [15]),
    .X(net481));
 sg13g2_buf_2 fanout482 (.A(\median_processor.input_storage [13]),
    .X(net482));
 sg13g2_buf_2 fanout483 (.A(\median_processor.input_storage [12]),
    .X(net483));
 sg13g2_buf_2 fanout484 (.A(\median_processor.input_storage [0]),
    .X(net484));
 sg13g2_buf_2 fanout485 (.A(_05020_),
    .X(net485));
 sg13g2_buf_2 fanout486 (.A(_05017_),
    .X(net486));
 sg13g2_buf_2 fanout487 (.A(_05015_),
    .X(net487));
 sg13g2_buf_2 fanout488 (.A(_02939_),
    .X(net488));
 sg13g2_buf_2 fanout489 (.A(_02932_),
    .X(net489));
 sg13g2_buf_2 fanout490 (.A(_02927_),
    .X(net490));
 sg13g2_buf_2 fanout491 (.A(_02925_),
    .X(net491));
 sg13g2_buf_2 fanout492 (.A(_02923_),
    .X(net492));
 sg13g2_buf_2 fanout493 (.A(_02912_),
    .X(net493));
 sg13g2_buf_2 fanout494 (.A(_02909_),
    .X(net494));
 sg13g2_buf_2 fanout495 (.A(data_in_p2c_7),
    .X(net495));
 sg13g2_tiehi \median_processor.input_storage[0]$_SDFFE_PN0P__496  (.L_HI(net496));
 sg13g2_tiehi \median_processor.input_storage[10]$_SDFFE_PN0P__497  (.L_HI(net497));
 sg13g2_tiehi \median_processor.input_storage[11]$_SDFFE_PN0P__498  (.L_HI(net498));
 sg13g2_tiehi \median_processor.input_storage[12]$_SDFFE_PN0P__499  (.L_HI(net499));
 sg13g2_tiehi \median_processor.input_storage[13]$_SDFFE_PN0P__500  (.L_HI(net500));
 sg13g2_tiehi \median_processor.input_storage[14]$_SDFFE_PN0P__501  (.L_HI(net501));
 sg13g2_tiehi \median_processor.input_storage[15]$_SDFFE_PN0P__502  (.L_HI(net502));
 sg13g2_tiehi \median_processor.input_storage[16]$_SDFFE_PN0P__503  (.L_HI(net503));
 sg13g2_tiehi \median_processor.input_storage[17]$_SDFFE_PN0P__504  (.L_HI(net504));
 sg13g2_tiehi \median_processor.input_storage[18]$_SDFFE_PN0P__505  (.L_HI(net505));
 sg13g2_tiehi \median_processor.input_storage[19]$_SDFFE_PN0P__506  (.L_HI(net506));
 sg13g2_tiehi \median_processor.input_storage[1]$_SDFFE_PN0P__507  (.L_HI(net507));
 sg13g2_tiehi \median_processor.input_storage[20]$_SDFFE_PN0P__508  (.L_HI(net508));
 sg13g2_tiehi \median_processor.input_storage[21]$_SDFFE_PN0P__509  (.L_HI(net509));
 sg13g2_tiehi \median_processor.input_storage[22]$_SDFFE_PN0P__510  (.L_HI(net510));
 sg13g2_tiehi \median_processor.input_storage[23]$_SDFFE_PN0P__511  (.L_HI(net511));
 sg13g2_tiehi \median_processor.input_storage[24]$_SDFFE_PN0P__512  (.L_HI(net512));
 sg13g2_tiehi \median_processor.input_storage[25]$_SDFFE_PN0P__513  (.L_HI(net513));
 sg13g2_tiehi \median_processor.input_storage[26]$_SDFFE_PN0P__514  (.L_HI(net514));
 sg13g2_tiehi \median_processor.input_storage[27]$_SDFFE_PN0P__515  (.L_HI(net515));
 sg13g2_tiehi \median_processor.input_storage[28]$_SDFFE_PN0P__516  (.L_HI(net516));
 sg13g2_tiehi \median_processor.input_storage[29]$_SDFFE_PN0P__517  (.L_HI(net517));
 sg13g2_tiehi \median_processor.input_storage[2]$_SDFFE_PN0P__518  (.L_HI(net518));
 sg13g2_tiehi \median_processor.input_storage[30]$_SDFFE_PN0P__519  (.L_HI(net519));
 sg13g2_tiehi \median_processor.input_storage[31]$_SDFFE_PN0P__520  (.L_HI(net520));
 sg13g2_tiehi \median_processor.input_storage[32]$_SDFFE_PN0P__521  (.L_HI(net521));
 sg13g2_tiehi \median_processor.input_storage[33]$_SDFFE_PN0P__522  (.L_HI(net522));
 sg13g2_tiehi \median_processor.input_storage[34]$_SDFFE_PN0P__523  (.L_HI(net523));
 sg13g2_tiehi \median_processor.input_storage[35]$_SDFFE_PN0P__524  (.L_HI(net524));
 sg13g2_tiehi \median_processor.input_storage[36]$_SDFFE_PN0P__525  (.L_HI(net525));
 sg13g2_tiehi \median_processor.input_storage[37]$_SDFFE_PN0P__526  (.L_HI(net526));
 sg13g2_tiehi \median_processor.input_storage[38]$_SDFFE_PN0P__527  (.L_HI(net527));
 sg13g2_tiehi \median_processor.input_storage[39]$_SDFFE_PN0P__528  (.L_HI(net528));
 sg13g2_tiehi \median_processor.input_storage[3]$_SDFFE_PN0P__529  (.L_HI(net529));
 sg13g2_tiehi \median_processor.input_storage[40]$_SDFFE_PN0P__530  (.L_HI(net530));
 sg13g2_tiehi \median_processor.input_storage[41]$_SDFFE_PN0P__531  (.L_HI(net531));
 sg13g2_tiehi \median_processor.input_storage[42]$_SDFFE_PN0P__532  (.L_HI(net532));
 sg13g2_tiehi \median_processor.input_storage[43]$_SDFFE_PN0P__533  (.L_HI(net533));
 sg13g2_tiehi \median_processor.input_storage[44]$_SDFFE_PN0P__534  (.L_HI(net534));
 sg13g2_tiehi \median_processor.input_storage[45]$_SDFFE_PN0P__535  (.L_HI(net535));
 sg13g2_tiehi \median_processor.input_storage[46]$_SDFFE_PN0P__536  (.L_HI(net536));
 sg13g2_tiehi \median_processor.input_storage[47]$_SDFFE_PN0P__537  (.L_HI(net537));
 sg13g2_tiehi \median_processor.input_storage[48]$_SDFFE_PN0P__538  (.L_HI(net538));
 sg13g2_tiehi \median_processor.input_storage[49]$_SDFFE_PN0P__539  (.L_HI(net539));
 sg13g2_tiehi \median_processor.input_storage[4]$_SDFFE_PN0P__540  (.L_HI(net540));
 sg13g2_tiehi \median_processor.input_storage[50]$_SDFFE_PN0P__541  (.L_HI(net541));
 sg13g2_tiehi \median_processor.input_storage[51]$_SDFFE_PN0P__542  (.L_HI(net542));
 sg13g2_tiehi \median_processor.input_storage[52]$_SDFFE_PN0P__543  (.L_HI(net543));
 sg13g2_tiehi \median_processor.input_storage[53]$_SDFFE_PN0P__544  (.L_HI(net544));
 sg13g2_tiehi \median_processor.input_storage[54]$_SDFFE_PN0P__545  (.L_HI(net545));
 sg13g2_tiehi \median_processor.input_storage[55]$_SDFFE_PN0P__546  (.L_HI(net546));
 sg13g2_tiehi \median_processor.input_storage[56]$_SDFFE_PN0P__547  (.L_HI(net547));
 sg13g2_tiehi \median_processor.input_storage[57]$_SDFFE_PN0P__548  (.L_HI(net548));
 sg13g2_tiehi \median_processor.input_storage[58]$_SDFFE_PN0P__549  (.L_HI(net549));
 sg13g2_tiehi \median_processor.input_storage[59]$_SDFFE_PN0P__550  (.L_HI(net550));
 sg13g2_tiehi \median_processor.input_storage[5]$_SDFFE_PN0P__551  (.L_HI(net551));
 sg13g2_tiehi \median_processor.input_storage[60]$_SDFFE_PN0P__552  (.L_HI(net552));
 sg13g2_tiehi \median_processor.input_storage[61]$_SDFFE_PN0P__553  (.L_HI(net553));
 sg13g2_tiehi \median_processor.input_storage[62]$_SDFFE_PN0P__554  (.L_HI(net554));
 sg13g2_tiehi \median_processor.input_storage[63]$_SDFFE_PN0P__555  (.L_HI(net555));
 sg13g2_tiehi \median_processor.input_storage[6]$_SDFFE_PN0P__556  (.L_HI(net556));
 sg13g2_tiehi \median_processor.input_storage[7]$_SDFFE_PN0P__557  (.L_HI(net557));
 sg13g2_tiehi \median_processor.input_storage[8]$_SDFFE_PN0P__558  (.L_HI(net558));
 sg13g2_tiehi \median_processor.input_storage[9]$_SDFFE_PN0P__559  (.L_HI(net559));
 sg13g2_tiehi \median_processor.median_processor.median_out[0]$_DFFE_PP__560  (.L_HI(net560));
 sg13g2_tiehi \median_processor.median_processor.median_out[1]$_DFFE_PP__561  (.L_HI(net561));
 sg13g2_tiehi \median_processor.median_processor.median_out[2]$_DFFE_PP__562  (.L_HI(net562));
 sg13g2_tiehi \median_processor.median_processor.median_out[3]$_DFFE_PP__563  (.L_HI(net563));
 sg13g2_tiehi \median_processor.median_processor.median_out[4]$_DFFE_PP__564  (.L_HI(net564));
 sg13g2_tiehi \median_processor.median_processor.median_out[5]$_DFFE_PP__565  (.L_HI(net565));
 sg13g2_tiehi \median_processor.median_processor.median_out[6]$_DFFE_PP__566  (.L_HI(net566));
 sg13g2_tiehi \median_processor.median_processor.median_out[7]$_DFFE_PP__567  (.L_HI(net567));
 sg13g2_tiehi \rando_generator.lfsr_reg[0]$_SDFF_PN0__568  (.L_HI(net568));
 sg13g2_tiehi \rando_generator.lfsr_reg[10]$_SDFF_PN0__569  (.L_HI(net569));
 sg13g2_tiehi \rando_generator.lfsr_reg[11]$_SDFF_PN0__570  (.L_HI(net570));
 sg13g2_tiehi \rando_generator.lfsr_reg[12]$_SDFF_PN0__571  (.L_HI(net571));
 sg13g2_tiehi \rando_generator.lfsr_reg[13]$_SDFF_PN0__572  (.L_HI(net572));
 sg13g2_tiehi \rando_generator.lfsr_reg[14]$_SDFF_PN0__573  (.L_HI(net573));
 sg13g2_tiehi \rando_generator.lfsr_reg[15]$_SDFF_PN0__574  (.L_HI(net574));
 sg13g2_tiehi \rando_generator.lfsr_reg[16]$_SDFF_PN0__575  (.L_HI(net575));
 sg13g2_tiehi \rando_generator.lfsr_reg[17]$_SDFF_PN0__576  (.L_HI(net576));
 sg13g2_tiehi \rando_generator.lfsr_reg[18]$_SDFF_PN0__577  (.L_HI(net577));
 sg13g2_tiehi \rando_generator.lfsr_reg[19]$_SDFF_PN0__578  (.L_HI(net578));
 sg13g2_tiehi \rando_generator.lfsr_reg[1]$_SDFF_PN0__579  (.L_HI(net579));
 sg13g2_tiehi \rando_generator.lfsr_reg[20]$_SDFF_PN0__580  (.L_HI(net580));
 sg13g2_tiehi \rando_generator.lfsr_reg[21]$_SDFF_PN0__581  (.L_HI(net581));
 sg13g2_tiehi \rando_generator.lfsr_reg[22]$_SDFF_PN0__582  (.L_HI(net582));
 sg13g2_tiehi \rando_generator.lfsr_reg[23]$_SDFF_PN0__583  (.L_HI(net583));
 sg13g2_tiehi \rando_generator.lfsr_reg[24]$_SDFF_PN0__584  (.L_HI(net584));
 sg13g2_tiehi \rando_generator.lfsr_reg[25]$_SDFF_PN0__585  (.L_HI(net585));
 sg13g2_tiehi \rando_generator.lfsr_reg[26]$_SDFF_PN0__586  (.L_HI(net586));
 sg13g2_tiehi \rando_generator.lfsr_reg[27]$_SDFF_PN0__587  (.L_HI(net587));
 sg13g2_tiehi \rando_generator.lfsr_reg[28]$_SDFF_PN0__588  (.L_HI(net588));
 sg13g2_tiehi \rando_generator.lfsr_reg[29]$_SDFF_PN0__589  (.L_HI(net589));
 sg13g2_tiehi \rando_generator.lfsr_reg[2]$_SDFF_PN0__590  (.L_HI(net590));
 sg13g2_tiehi \rando_generator.lfsr_reg[30]$_SDFF_PN0__591  (.L_HI(net591));
 sg13g2_tiehi \rando_generator.lfsr_reg[3]$_SDFF_PN0__592  (.L_HI(net592));
 sg13g2_tiehi \rando_generator.lfsr_reg[4]$_SDFF_PN0__593  (.L_HI(net593));
 sg13g2_tiehi \rando_generator.lfsr_reg[5]$_SDFF_PN0__594  (.L_HI(net594));
 sg13g2_tiehi \rando_generator.lfsr_reg[6]$_SDFF_PN0__595  (.L_HI(net595));
 sg13g2_tiehi \rando_generator.lfsr_reg[7]$_SDFF_PN0__596  (.L_HI(net596));
 sg13g2_tiehi \rando_generator.lfsr_reg[8]$_SDFF_PN0__597  (.L_HI(net597));
 sg13g2_tiehi \rando_generator.lfsr_reg[9]$_SDFF_PN0__598  (.L_HI(net598));
 sg13g2_tiehi \shift_storage.storage[0]$_SDFFE_PN0P__599  (.L_HI(net599));
 sg13g2_tiehi \shift_storage.storage[1000]$_SDFFE_PN0P__600  (.L_HI(net600));
 sg13g2_tiehi \shift_storage.storage[1001]$_SDFFE_PN0P__601  (.L_HI(net601));
 sg13g2_tiehi \shift_storage.storage[1002]$_SDFFE_PN0P__602  (.L_HI(net602));
 sg13g2_tiehi \shift_storage.storage[1003]$_SDFFE_PN0P__603  (.L_HI(net603));
 sg13g2_tiehi \shift_storage.storage[1004]$_SDFFE_PN0P__604  (.L_HI(net604));
 sg13g2_tiehi \shift_storage.storage[1005]$_SDFFE_PN0P__605  (.L_HI(net605));
 sg13g2_tiehi \shift_storage.storage[1006]$_SDFFE_PN0P__606  (.L_HI(net606));
 sg13g2_tiehi \shift_storage.storage[1007]$_SDFFE_PN0P__607  (.L_HI(net607));
 sg13g2_tiehi \shift_storage.storage[1008]$_SDFFE_PN0P__608  (.L_HI(net608));
 sg13g2_tiehi \shift_storage.storage[1009]$_SDFFE_PN0P__609  (.L_HI(net609));
 sg13g2_tiehi \shift_storage.storage[100]$_SDFFE_PN0P__610  (.L_HI(net610));
 sg13g2_tiehi \shift_storage.storage[1010]$_SDFFE_PN0P__611  (.L_HI(net611));
 sg13g2_tiehi \shift_storage.storage[1011]$_SDFFE_PN0P__612  (.L_HI(net612));
 sg13g2_tiehi \shift_storage.storage[1012]$_SDFFE_PN0P__613  (.L_HI(net613));
 sg13g2_tiehi \shift_storage.storage[1013]$_SDFFE_PN0P__614  (.L_HI(net614));
 sg13g2_tiehi \shift_storage.storage[1014]$_SDFFE_PN0P__615  (.L_HI(net615));
 sg13g2_tiehi \shift_storage.storage[1015]$_SDFFE_PN0P__616  (.L_HI(net616));
 sg13g2_tiehi \shift_storage.storage[1016]$_SDFFE_PN0P__617  (.L_HI(net617));
 sg13g2_tiehi \shift_storage.storage[1017]$_SDFFE_PN0P__618  (.L_HI(net618));
 sg13g2_tiehi \shift_storage.storage[1018]$_SDFFE_PN0P__619  (.L_HI(net619));
 sg13g2_tiehi \shift_storage.storage[1019]$_SDFFE_PN0P__620  (.L_HI(net620));
 sg13g2_tiehi \shift_storage.storage[101]$_SDFFE_PN0P__621  (.L_HI(net621));
 sg13g2_tiehi \shift_storage.storage[1020]$_SDFFE_PN0P__622  (.L_HI(net622));
 sg13g2_tiehi \shift_storage.storage[1021]$_SDFFE_PN0P__623  (.L_HI(net623));
 sg13g2_tiehi \shift_storage.storage[1022]$_SDFFE_PN0P__624  (.L_HI(net624));
 sg13g2_tiehi \shift_storage.storage[1023]$_SDFFE_PN0P__625  (.L_HI(net625));
 sg13g2_tiehi \shift_storage.storage[1024]$_SDFFE_PN0P__626  (.L_HI(net626));
 sg13g2_tiehi \shift_storage.storage[1025]$_SDFFE_PN0P__627  (.L_HI(net627));
 sg13g2_tiehi \shift_storage.storage[1026]$_SDFFE_PN0P__628  (.L_HI(net628));
 sg13g2_tiehi \shift_storage.storage[1027]$_SDFFE_PN0P__629  (.L_HI(net629));
 sg13g2_tiehi \shift_storage.storage[1028]$_SDFFE_PN0P__630  (.L_HI(net630));
 sg13g2_tiehi \shift_storage.storage[1029]$_SDFFE_PN0P__631  (.L_HI(net631));
 sg13g2_tiehi \shift_storage.storage[102]$_SDFFE_PN0P__632  (.L_HI(net632));
 sg13g2_tiehi \shift_storage.storage[1030]$_SDFFE_PN0P__633  (.L_HI(net633));
 sg13g2_tiehi \shift_storage.storage[1031]$_SDFFE_PN0P__634  (.L_HI(net634));
 sg13g2_tiehi \shift_storage.storage[1032]$_SDFFE_PN0P__635  (.L_HI(net635));
 sg13g2_tiehi \shift_storage.storage[1033]$_SDFFE_PN0P__636  (.L_HI(net636));
 sg13g2_tiehi \shift_storage.storage[1034]$_SDFFE_PN0P__637  (.L_HI(net637));
 sg13g2_tiehi \shift_storage.storage[1035]$_SDFFE_PN0P__638  (.L_HI(net638));
 sg13g2_tiehi \shift_storage.storage[1036]$_SDFFE_PN0P__639  (.L_HI(net639));
 sg13g2_tiehi \shift_storage.storage[1037]$_SDFFE_PN0P__640  (.L_HI(net640));
 sg13g2_tiehi \shift_storage.storage[1038]$_SDFFE_PN0P__641  (.L_HI(net641));
 sg13g2_tiehi \shift_storage.storage[1039]$_SDFFE_PN0P__642  (.L_HI(net642));
 sg13g2_tiehi \shift_storage.storage[103]$_SDFFE_PN0P__643  (.L_HI(net643));
 sg13g2_tiehi \shift_storage.storage[1040]$_SDFFE_PN0P__644  (.L_HI(net644));
 sg13g2_tiehi \shift_storage.storage[1041]$_SDFFE_PN0P__645  (.L_HI(net645));
 sg13g2_tiehi \shift_storage.storage[1042]$_SDFFE_PN0P__646  (.L_HI(net646));
 sg13g2_tiehi \shift_storage.storage[1043]$_SDFFE_PN0P__647  (.L_HI(net647));
 sg13g2_tiehi \shift_storage.storage[1044]$_SDFFE_PN0P__648  (.L_HI(net648));
 sg13g2_tiehi \shift_storage.storage[1045]$_SDFFE_PN0P__649  (.L_HI(net649));
 sg13g2_tiehi \shift_storage.storage[1046]$_SDFFE_PN0P__650  (.L_HI(net650));
 sg13g2_tiehi \shift_storage.storage[1047]$_SDFFE_PN0P__651  (.L_HI(net651));
 sg13g2_tiehi \shift_storage.storage[1048]$_SDFFE_PN0P__652  (.L_HI(net652));
 sg13g2_tiehi \shift_storage.storage[1049]$_SDFFE_PN0P__653  (.L_HI(net653));
 sg13g2_tiehi \shift_storage.storage[104]$_SDFFE_PN0P__654  (.L_HI(net654));
 sg13g2_tiehi \shift_storage.storage[1050]$_SDFFE_PN0P__655  (.L_HI(net655));
 sg13g2_tiehi \shift_storage.storage[1051]$_SDFFE_PN0P__656  (.L_HI(net656));
 sg13g2_tiehi \shift_storage.storage[1052]$_SDFFE_PN0P__657  (.L_HI(net657));
 sg13g2_tiehi \shift_storage.storage[1053]$_SDFFE_PN0P__658  (.L_HI(net658));
 sg13g2_tiehi \shift_storage.storage[1054]$_SDFFE_PN0P__659  (.L_HI(net659));
 sg13g2_tiehi \shift_storage.storage[1055]$_SDFFE_PN0P__660  (.L_HI(net660));
 sg13g2_tiehi \shift_storage.storage[1056]$_SDFFE_PN0P__661  (.L_HI(net661));
 sg13g2_tiehi \shift_storage.storage[1057]$_SDFFE_PN0P__662  (.L_HI(net662));
 sg13g2_tiehi \shift_storage.storage[1058]$_SDFFE_PN0P__663  (.L_HI(net663));
 sg13g2_tiehi \shift_storage.storage[1059]$_SDFFE_PN0P__664  (.L_HI(net664));
 sg13g2_tiehi \shift_storage.storage[105]$_SDFFE_PN0P__665  (.L_HI(net665));
 sg13g2_tiehi \shift_storage.storage[1060]$_SDFFE_PN0P__666  (.L_HI(net666));
 sg13g2_tiehi \shift_storage.storage[1061]$_SDFFE_PN0P__667  (.L_HI(net667));
 sg13g2_tiehi \shift_storage.storage[1062]$_SDFFE_PN0P__668  (.L_HI(net668));
 sg13g2_tiehi \shift_storage.storage[1063]$_SDFFE_PN0P__669  (.L_HI(net669));
 sg13g2_tiehi \shift_storage.storage[1064]$_SDFFE_PN0P__670  (.L_HI(net670));
 sg13g2_tiehi \shift_storage.storage[1065]$_SDFFE_PN0P__671  (.L_HI(net671));
 sg13g2_tiehi \shift_storage.storage[1066]$_SDFFE_PN0P__672  (.L_HI(net672));
 sg13g2_tiehi \shift_storage.storage[1067]$_SDFFE_PN0P__673  (.L_HI(net673));
 sg13g2_tiehi \shift_storage.storage[1068]$_SDFFE_PN0P__674  (.L_HI(net674));
 sg13g2_tiehi \shift_storage.storage[1069]$_SDFFE_PN0P__675  (.L_HI(net675));
 sg13g2_tiehi \shift_storage.storage[106]$_SDFFE_PN0P__676  (.L_HI(net676));
 sg13g2_tiehi \shift_storage.storage[1070]$_SDFFE_PN0P__677  (.L_HI(net677));
 sg13g2_tiehi \shift_storage.storage[1071]$_SDFFE_PN0P__678  (.L_HI(net678));
 sg13g2_tiehi \shift_storage.storage[1072]$_SDFFE_PN0P__679  (.L_HI(net679));
 sg13g2_tiehi \shift_storage.storage[1073]$_SDFFE_PN0P__680  (.L_HI(net680));
 sg13g2_tiehi \shift_storage.storage[1074]$_SDFFE_PN0P__681  (.L_HI(net681));
 sg13g2_tiehi \shift_storage.storage[1075]$_SDFFE_PN0P__682  (.L_HI(net682));
 sg13g2_tiehi \shift_storage.storage[1076]$_SDFFE_PN0P__683  (.L_HI(net683));
 sg13g2_tiehi \shift_storage.storage[1077]$_SDFFE_PN0P__684  (.L_HI(net684));
 sg13g2_tiehi \shift_storage.storage[1078]$_SDFFE_PN0P__685  (.L_HI(net685));
 sg13g2_tiehi \shift_storage.storage[1079]$_SDFFE_PN0P__686  (.L_HI(net686));
 sg13g2_tiehi \shift_storage.storage[107]$_SDFFE_PN0P__687  (.L_HI(net687));
 sg13g2_tiehi \shift_storage.storage[1080]$_SDFFE_PN0P__688  (.L_HI(net688));
 sg13g2_tiehi \shift_storage.storage[1081]$_SDFFE_PN0P__689  (.L_HI(net689));
 sg13g2_tiehi \shift_storage.storage[1082]$_SDFFE_PN0P__690  (.L_HI(net690));
 sg13g2_tiehi \shift_storage.storage[1083]$_SDFFE_PN0P__691  (.L_HI(net691));
 sg13g2_tiehi \shift_storage.storage[1084]$_SDFFE_PN0P__692  (.L_HI(net692));
 sg13g2_tiehi \shift_storage.storage[1085]$_SDFFE_PN0P__693  (.L_HI(net693));
 sg13g2_tiehi \shift_storage.storage[1086]$_SDFFE_PN0P__694  (.L_HI(net694));
 sg13g2_tiehi \shift_storage.storage[1087]$_SDFFE_PN0P__695  (.L_HI(net695));
 sg13g2_tiehi \shift_storage.storage[1088]$_SDFFE_PN0P__696  (.L_HI(net696));
 sg13g2_tiehi \shift_storage.storage[1089]$_SDFFE_PN0P__697  (.L_HI(net697));
 sg13g2_tiehi \shift_storage.storage[108]$_SDFFE_PN0P__698  (.L_HI(net698));
 sg13g2_tiehi \shift_storage.storage[1090]$_SDFFE_PN0P__699  (.L_HI(net699));
 sg13g2_tiehi \shift_storage.storage[1091]$_SDFFE_PN0P__700  (.L_HI(net700));
 sg13g2_tiehi \shift_storage.storage[1092]$_SDFFE_PN0P__701  (.L_HI(net701));
 sg13g2_tiehi \shift_storage.storage[1093]$_SDFFE_PN0P__702  (.L_HI(net702));
 sg13g2_tiehi \shift_storage.storage[1094]$_SDFFE_PN0P__703  (.L_HI(net703));
 sg13g2_tiehi \shift_storage.storage[1095]$_SDFFE_PN0P__704  (.L_HI(net704));
 sg13g2_tiehi \shift_storage.storage[1096]$_SDFFE_PN0P__705  (.L_HI(net705));
 sg13g2_tiehi \shift_storage.storage[1097]$_SDFFE_PN0P__706  (.L_HI(net706));
 sg13g2_tiehi \shift_storage.storage[1098]$_SDFFE_PN0P__707  (.L_HI(net707));
 sg13g2_tiehi \shift_storage.storage[1099]$_SDFFE_PN0P__708  (.L_HI(net708));
 sg13g2_tiehi \shift_storage.storage[109]$_SDFFE_PN0P__709  (.L_HI(net709));
 sg13g2_tiehi \shift_storage.storage[10]$_SDFFE_PN0P__710  (.L_HI(net710));
 sg13g2_tiehi \shift_storage.storage[1100]$_SDFFE_PN0P__711  (.L_HI(net711));
 sg13g2_tiehi \shift_storage.storage[1101]$_SDFFE_PN0P__712  (.L_HI(net712));
 sg13g2_tiehi \shift_storage.storage[1102]$_SDFFE_PN0P__713  (.L_HI(net713));
 sg13g2_tiehi \shift_storage.storage[1103]$_SDFFE_PN0P__714  (.L_HI(net714));
 sg13g2_tiehi \shift_storage.storage[1104]$_SDFFE_PN0P__715  (.L_HI(net715));
 sg13g2_tiehi \shift_storage.storage[1105]$_SDFFE_PN0P__716  (.L_HI(net716));
 sg13g2_tiehi \shift_storage.storage[1106]$_SDFFE_PN0P__717  (.L_HI(net717));
 sg13g2_tiehi \shift_storage.storage[1107]$_SDFFE_PN0P__718  (.L_HI(net718));
 sg13g2_tiehi \shift_storage.storage[1108]$_SDFFE_PN0P__719  (.L_HI(net719));
 sg13g2_tiehi \shift_storage.storage[1109]$_SDFFE_PN0P__720  (.L_HI(net720));
 sg13g2_tiehi \shift_storage.storage[110]$_SDFFE_PN0P__721  (.L_HI(net721));
 sg13g2_tiehi \shift_storage.storage[1110]$_SDFFE_PN0P__722  (.L_HI(net722));
 sg13g2_tiehi \shift_storage.storage[1111]$_SDFFE_PN0P__723  (.L_HI(net723));
 sg13g2_tiehi \shift_storage.storage[1112]$_SDFFE_PN0P__724  (.L_HI(net724));
 sg13g2_tiehi \shift_storage.storage[1113]$_SDFFE_PN0P__725  (.L_HI(net725));
 sg13g2_tiehi \shift_storage.storage[1114]$_SDFFE_PN0P__726  (.L_HI(net726));
 sg13g2_tiehi \shift_storage.storage[1115]$_SDFFE_PN0P__727  (.L_HI(net727));
 sg13g2_tiehi \shift_storage.storage[1116]$_SDFFE_PN0P__728  (.L_HI(net728));
 sg13g2_tiehi \shift_storage.storage[1117]$_SDFFE_PN0P__729  (.L_HI(net729));
 sg13g2_tiehi \shift_storage.storage[1118]$_SDFFE_PN0P__730  (.L_HI(net730));
 sg13g2_tiehi \shift_storage.storage[1119]$_SDFFE_PN0P__731  (.L_HI(net731));
 sg13g2_tiehi \shift_storage.storage[111]$_SDFFE_PN0P__732  (.L_HI(net732));
 sg13g2_tiehi \shift_storage.storage[1120]$_SDFFE_PN0P__733  (.L_HI(net733));
 sg13g2_tiehi \shift_storage.storage[1121]$_SDFFE_PN0P__734  (.L_HI(net734));
 sg13g2_tiehi \shift_storage.storage[1122]$_SDFFE_PN0P__735  (.L_HI(net735));
 sg13g2_tiehi \shift_storage.storage[1123]$_SDFFE_PN0P__736  (.L_HI(net736));
 sg13g2_tiehi \shift_storage.storage[1124]$_SDFFE_PN0P__737  (.L_HI(net737));
 sg13g2_tiehi \shift_storage.storage[1125]$_SDFFE_PN0P__738  (.L_HI(net738));
 sg13g2_tiehi \shift_storage.storage[1126]$_SDFFE_PN0P__739  (.L_HI(net739));
 sg13g2_tiehi \shift_storage.storage[1127]$_SDFFE_PN0P__740  (.L_HI(net740));
 sg13g2_tiehi \shift_storage.storage[1128]$_SDFFE_PN0P__741  (.L_HI(net741));
 sg13g2_tiehi \shift_storage.storage[1129]$_SDFFE_PN0P__742  (.L_HI(net742));
 sg13g2_tiehi \shift_storage.storage[112]$_SDFFE_PN0P__743  (.L_HI(net743));
 sg13g2_tiehi \shift_storage.storage[1130]$_SDFFE_PN0P__744  (.L_HI(net744));
 sg13g2_tiehi \shift_storage.storage[1131]$_SDFFE_PN0P__745  (.L_HI(net745));
 sg13g2_tiehi \shift_storage.storage[1132]$_SDFFE_PN0P__746  (.L_HI(net746));
 sg13g2_tiehi \shift_storage.storage[1133]$_SDFFE_PN0P__747  (.L_HI(net747));
 sg13g2_tiehi \shift_storage.storage[1134]$_SDFFE_PN0P__748  (.L_HI(net748));
 sg13g2_tiehi \shift_storage.storage[1135]$_SDFFE_PN0P__749  (.L_HI(net749));
 sg13g2_tiehi \shift_storage.storage[1136]$_SDFFE_PN0P__750  (.L_HI(net750));
 sg13g2_tiehi \shift_storage.storage[1137]$_SDFFE_PN0P__751  (.L_HI(net751));
 sg13g2_tiehi \shift_storage.storage[1138]$_SDFFE_PN0P__752  (.L_HI(net752));
 sg13g2_tiehi \shift_storage.storage[1139]$_SDFFE_PN0P__753  (.L_HI(net753));
 sg13g2_tiehi \shift_storage.storage[113]$_SDFFE_PN0P__754  (.L_HI(net754));
 sg13g2_tiehi \shift_storage.storage[1140]$_SDFFE_PN0P__755  (.L_HI(net755));
 sg13g2_tiehi \shift_storage.storage[1141]$_SDFFE_PN0P__756  (.L_HI(net756));
 sg13g2_tiehi \shift_storage.storage[1142]$_SDFFE_PN0P__757  (.L_HI(net757));
 sg13g2_tiehi \shift_storage.storage[1143]$_SDFFE_PN0P__758  (.L_HI(net758));
 sg13g2_tiehi \shift_storage.storage[1144]$_SDFFE_PN0P__759  (.L_HI(net759));
 sg13g2_tiehi \shift_storage.storage[1145]$_SDFFE_PN0P__760  (.L_HI(net760));
 sg13g2_tiehi \shift_storage.storage[1146]$_SDFFE_PN0P__761  (.L_HI(net761));
 sg13g2_tiehi \shift_storage.storage[1147]$_SDFFE_PN0P__762  (.L_HI(net762));
 sg13g2_tiehi \shift_storage.storage[1148]$_SDFFE_PN0P__763  (.L_HI(net763));
 sg13g2_tiehi \shift_storage.storage[1149]$_SDFFE_PN0P__764  (.L_HI(net764));
 sg13g2_tiehi \shift_storage.storage[114]$_SDFFE_PN0P__765  (.L_HI(net765));
 sg13g2_tiehi \shift_storage.storage[1150]$_SDFFE_PN0P__766  (.L_HI(net766));
 sg13g2_tiehi \shift_storage.storage[1151]$_SDFFE_PN0P__767  (.L_HI(net767));
 sg13g2_tiehi \shift_storage.storage[1152]$_SDFFE_PN0P__768  (.L_HI(net768));
 sg13g2_tiehi \shift_storage.storage[1153]$_SDFFE_PN0P__769  (.L_HI(net769));
 sg13g2_tiehi \shift_storage.storage[1154]$_SDFFE_PN0P__770  (.L_HI(net770));
 sg13g2_tiehi \shift_storage.storage[1155]$_SDFFE_PN0P__771  (.L_HI(net771));
 sg13g2_tiehi \shift_storage.storage[1156]$_SDFFE_PN0P__772  (.L_HI(net772));
 sg13g2_tiehi \shift_storage.storage[1157]$_SDFFE_PN0P__773  (.L_HI(net773));
 sg13g2_tiehi \shift_storage.storage[1158]$_SDFFE_PN0P__774  (.L_HI(net774));
 sg13g2_tiehi \shift_storage.storage[1159]$_SDFFE_PN0P__775  (.L_HI(net775));
 sg13g2_tiehi \shift_storage.storage[115]$_SDFFE_PN0P__776  (.L_HI(net776));
 sg13g2_tiehi \shift_storage.storage[1160]$_SDFFE_PN0P__777  (.L_HI(net777));
 sg13g2_tiehi \shift_storage.storage[1161]$_SDFFE_PN0P__778  (.L_HI(net778));
 sg13g2_tiehi \shift_storage.storage[1162]$_SDFFE_PN0P__779  (.L_HI(net779));
 sg13g2_tiehi \shift_storage.storage[1163]$_SDFFE_PN0P__780  (.L_HI(net780));
 sg13g2_tiehi \shift_storage.storage[1164]$_SDFFE_PN0P__781  (.L_HI(net781));
 sg13g2_tiehi \shift_storage.storage[1165]$_SDFFE_PN0P__782  (.L_HI(net782));
 sg13g2_tiehi \shift_storage.storage[1166]$_SDFFE_PN0P__783  (.L_HI(net783));
 sg13g2_tiehi \shift_storage.storage[1167]$_SDFFE_PN0P__784  (.L_HI(net784));
 sg13g2_tiehi \shift_storage.storage[1168]$_SDFFE_PN0P__785  (.L_HI(net785));
 sg13g2_tiehi \shift_storage.storage[1169]$_SDFFE_PN0P__786  (.L_HI(net786));
 sg13g2_tiehi \shift_storage.storage[116]$_SDFFE_PN0P__787  (.L_HI(net787));
 sg13g2_tiehi \shift_storage.storage[1170]$_SDFFE_PN0P__788  (.L_HI(net788));
 sg13g2_tiehi \shift_storage.storage[1171]$_SDFFE_PN0P__789  (.L_HI(net789));
 sg13g2_tiehi \shift_storage.storage[1172]$_SDFFE_PN0P__790  (.L_HI(net790));
 sg13g2_tiehi \shift_storage.storage[1173]$_SDFFE_PN0P__791  (.L_HI(net791));
 sg13g2_tiehi \shift_storage.storage[1174]$_SDFFE_PN0P__792  (.L_HI(net792));
 sg13g2_tiehi \shift_storage.storage[1175]$_SDFFE_PN0P__793  (.L_HI(net793));
 sg13g2_tiehi \shift_storage.storage[1176]$_SDFFE_PN0P__794  (.L_HI(net794));
 sg13g2_tiehi \shift_storage.storage[1177]$_SDFFE_PN0P__795  (.L_HI(net795));
 sg13g2_tiehi \shift_storage.storage[1178]$_SDFFE_PN0P__796  (.L_HI(net796));
 sg13g2_tiehi \shift_storage.storage[1179]$_SDFFE_PN0P__797  (.L_HI(net797));
 sg13g2_tiehi \shift_storage.storage[117]$_SDFFE_PN0P__798  (.L_HI(net798));
 sg13g2_tiehi \shift_storage.storage[1180]$_SDFFE_PN0P__799  (.L_HI(net799));
 sg13g2_tiehi \shift_storage.storage[1181]$_SDFFE_PN0P__800  (.L_HI(net800));
 sg13g2_tiehi \shift_storage.storage[1182]$_SDFFE_PN0P__801  (.L_HI(net801));
 sg13g2_tiehi \shift_storage.storage[1183]$_SDFFE_PN0P__802  (.L_HI(net802));
 sg13g2_tiehi \shift_storage.storage[1184]$_SDFFE_PN0P__803  (.L_HI(net803));
 sg13g2_tiehi \shift_storage.storage[1185]$_SDFFE_PN0P__804  (.L_HI(net804));
 sg13g2_tiehi \shift_storage.storage[1186]$_SDFFE_PN0P__805  (.L_HI(net805));
 sg13g2_tiehi \shift_storage.storage[1187]$_SDFFE_PN0P__806  (.L_HI(net806));
 sg13g2_tiehi \shift_storage.storage[1188]$_SDFFE_PN0P__807  (.L_HI(net807));
 sg13g2_tiehi \shift_storage.storage[1189]$_SDFFE_PN0P__808  (.L_HI(net808));
 sg13g2_tiehi \shift_storage.storage[118]$_SDFFE_PN0P__809  (.L_HI(net809));
 sg13g2_tiehi \shift_storage.storage[1190]$_SDFFE_PN0P__810  (.L_HI(net810));
 sg13g2_tiehi \shift_storage.storage[1191]$_SDFFE_PN0P__811  (.L_HI(net811));
 sg13g2_tiehi \shift_storage.storage[1192]$_SDFFE_PN0P__812  (.L_HI(net812));
 sg13g2_tiehi \shift_storage.storage[1193]$_SDFFE_PN0P__813  (.L_HI(net813));
 sg13g2_tiehi \shift_storage.storage[1194]$_SDFFE_PN0P__814  (.L_HI(net814));
 sg13g2_tiehi \shift_storage.storage[1195]$_SDFFE_PN0P__815  (.L_HI(net815));
 sg13g2_tiehi \shift_storage.storage[1196]$_SDFFE_PN0P__816  (.L_HI(net816));
 sg13g2_tiehi \shift_storage.storage[1197]$_SDFFE_PN0P__817  (.L_HI(net817));
 sg13g2_tiehi \shift_storage.storage[1198]$_SDFFE_PN0P__818  (.L_HI(net818));
 sg13g2_tiehi \shift_storage.storage[1199]$_SDFFE_PN0P__819  (.L_HI(net819));
 sg13g2_tiehi \shift_storage.storage[119]$_SDFFE_PN0P__820  (.L_HI(net820));
 sg13g2_tiehi \shift_storage.storage[11]$_SDFFE_PN0P__821  (.L_HI(net821));
 sg13g2_tiehi \shift_storage.storage[1200]$_SDFFE_PN0P__822  (.L_HI(net822));
 sg13g2_tiehi \shift_storage.storage[1201]$_SDFFE_PN0P__823  (.L_HI(net823));
 sg13g2_tiehi \shift_storage.storage[1202]$_SDFFE_PN0P__824  (.L_HI(net824));
 sg13g2_tiehi \shift_storage.storage[1203]$_SDFFE_PN0P__825  (.L_HI(net825));
 sg13g2_tiehi \shift_storage.storage[1204]$_SDFFE_PN0P__826  (.L_HI(net826));
 sg13g2_tiehi \shift_storage.storage[1205]$_SDFFE_PN0P__827  (.L_HI(net827));
 sg13g2_tiehi \shift_storage.storage[1206]$_SDFFE_PN0P__828  (.L_HI(net828));
 sg13g2_tiehi \shift_storage.storage[1207]$_SDFFE_PN0P__829  (.L_HI(net829));
 sg13g2_tiehi \shift_storage.storage[1208]$_SDFFE_PN0P__830  (.L_HI(net830));
 sg13g2_tiehi \shift_storage.storage[1209]$_SDFFE_PN0P__831  (.L_HI(net831));
 sg13g2_tiehi \shift_storage.storage[120]$_SDFFE_PN0P__832  (.L_HI(net832));
 sg13g2_tiehi \shift_storage.storage[1210]$_SDFFE_PN0P__833  (.L_HI(net833));
 sg13g2_tiehi \shift_storage.storage[1211]$_SDFFE_PN0P__834  (.L_HI(net834));
 sg13g2_tiehi \shift_storage.storage[1212]$_SDFFE_PN0P__835  (.L_HI(net835));
 sg13g2_tiehi \shift_storage.storage[1213]$_SDFFE_PN0P__836  (.L_HI(net836));
 sg13g2_tiehi \shift_storage.storage[1214]$_SDFFE_PN0P__837  (.L_HI(net837));
 sg13g2_tiehi \shift_storage.storage[1215]$_SDFFE_PN0P__838  (.L_HI(net838));
 sg13g2_tiehi \shift_storage.storage[1216]$_SDFFE_PN0P__839  (.L_HI(net839));
 sg13g2_tiehi \shift_storage.storage[1217]$_SDFFE_PN0P__840  (.L_HI(net840));
 sg13g2_tiehi \shift_storage.storage[1218]$_SDFFE_PN0P__841  (.L_HI(net841));
 sg13g2_tiehi \shift_storage.storage[1219]$_SDFFE_PN0P__842  (.L_HI(net842));
 sg13g2_tiehi \shift_storage.storage[121]$_SDFFE_PN0P__843  (.L_HI(net843));
 sg13g2_tiehi \shift_storage.storage[1220]$_SDFFE_PN0P__844  (.L_HI(net844));
 sg13g2_tiehi \shift_storage.storage[1221]$_SDFFE_PN0P__845  (.L_HI(net845));
 sg13g2_tiehi \shift_storage.storage[1222]$_SDFFE_PN0P__846  (.L_HI(net846));
 sg13g2_tiehi \shift_storage.storage[1223]$_SDFFE_PN0P__847  (.L_HI(net847));
 sg13g2_tiehi \shift_storage.storage[1224]$_SDFFE_PN0P__848  (.L_HI(net848));
 sg13g2_tiehi \shift_storage.storage[1225]$_SDFFE_PN0P__849  (.L_HI(net849));
 sg13g2_tiehi \shift_storage.storage[1226]$_SDFFE_PN0P__850  (.L_HI(net850));
 sg13g2_tiehi \shift_storage.storage[1227]$_SDFFE_PN0P__851  (.L_HI(net851));
 sg13g2_tiehi \shift_storage.storage[1228]$_SDFFE_PN0P__852  (.L_HI(net852));
 sg13g2_tiehi \shift_storage.storage[1229]$_SDFFE_PN0P__853  (.L_HI(net853));
 sg13g2_tiehi \shift_storage.storage[122]$_SDFFE_PN0P__854  (.L_HI(net854));
 sg13g2_tiehi \shift_storage.storage[1230]$_SDFFE_PN0P__855  (.L_HI(net855));
 sg13g2_tiehi \shift_storage.storage[1231]$_SDFFE_PN0P__856  (.L_HI(net856));
 sg13g2_tiehi \shift_storage.storage[1232]$_SDFFE_PN0P__857  (.L_HI(net857));
 sg13g2_tiehi \shift_storage.storage[1233]$_SDFFE_PN0P__858  (.L_HI(net858));
 sg13g2_tiehi \shift_storage.storage[1234]$_SDFFE_PN0P__859  (.L_HI(net859));
 sg13g2_tiehi \shift_storage.storage[1235]$_SDFFE_PN0P__860  (.L_HI(net860));
 sg13g2_tiehi \shift_storage.storage[1236]$_SDFFE_PN0P__861  (.L_HI(net861));
 sg13g2_tiehi \shift_storage.storage[1237]$_SDFFE_PN0P__862  (.L_HI(net862));
 sg13g2_tiehi \shift_storage.storage[1238]$_SDFFE_PN0P__863  (.L_HI(net863));
 sg13g2_tiehi \shift_storage.storage[1239]$_SDFFE_PN0P__864  (.L_HI(net864));
 sg13g2_tiehi \shift_storage.storage[123]$_SDFFE_PN0P__865  (.L_HI(net865));
 sg13g2_tiehi \shift_storage.storage[1240]$_SDFFE_PN0P__866  (.L_HI(net866));
 sg13g2_tiehi \shift_storage.storage[1241]$_SDFFE_PN0P__867  (.L_HI(net867));
 sg13g2_tiehi \shift_storage.storage[1242]$_SDFFE_PN0P__868  (.L_HI(net868));
 sg13g2_tiehi \shift_storage.storage[1243]$_SDFFE_PN0P__869  (.L_HI(net869));
 sg13g2_tiehi \shift_storage.storage[1244]$_SDFFE_PN0P__870  (.L_HI(net870));
 sg13g2_tiehi \shift_storage.storage[1245]$_SDFFE_PN0P__871  (.L_HI(net871));
 sg13g2_tiehi \shift_storage.storage[1246]$_SDFFE_PN0P__872  (.L_HI(net872));
 sg13g2_tiehi \shift_storage.storage[1247]$_SDFFE_PN0P__873  (.L_HI(net873));
 sg13g2_tiehi \shift_storage.storage[1248]$_SDFFE_PN0P__874  (.L_HI(net874));
 sg13g2_tiehi \shift_storage.storage[1249]$_SDFFE_PN0P__875  (.L_HI(net875));
 sg13g2_tiehi \shift_storage.storage[124]$_SDFFE_PN0P__876  (.L_HI(net876));
 sg13g2_tiehi \shift_storage.storage[1250]$_SDFFE_PN0P__877  (.L_HI(net877));
 sg13g2_tiehi \shift_storage.storage[1251]$_SDFFE_PN0P__878  (.L_HI(net878));
 sg13g2_tiehi \shift_storage.storage[1252]$_SDFFE_PN0P__879  (.L_HI(net879));
 sg13g2_tiehi \shift_storage.storage[1253]$_SDFFE_PN0P__880  (.L_HI(net880));
 sg13g2_tiehi \shift_storage.storage[1254]$_SDFFE_PN0P__881  (.L_HI(net881));
 sg13g2_tiehi \shift_storage.storage[1255]$_SDFFE_PN0P__882  (.L_HI(net882));
 sg13g2_tiehi \shift_storage.storage[1256]$_SDFFE_PN0P__883  (.L_HI(net883));
 sg13g2_tiehi \shift_storage.storage[1257]$_SDFFE_PN0P__884  (.L_HI(net884));
 sg13g2_tiehi \shift_storage.storage[1258]$_SDFFE_PN0P__885  (.L_HI(net885));
 sg13g2_tiehi \shift_storage.storage[1259]$_SDFFE_PN0P__886  (.L_HI(net886));
 sg13g2_tiehi \shift_storage.storage[125]$_SDFFE_PN0P__887  (.L_HI(net887));
 sg13g2_tiehi \shift_storage.storage[1260]$_SDFFE_PN0P__888  (.L_HI(net888));
 sg13g2_tiehi \shift_storage.storage[1261]$_SDFFE_PN0P__889  (.L_HI(net889));
 sg13g2_tiehi \shift_storage.storage[1262]$_SDFFE_PN0P__890  (.L_HI(net890));
 sg13g2_tiehi \shift_storage.storage[1263]$_SDFFE_PN0P__891  (.L_HI(net891));
 sg13g2_tiehi \shift_storage.storage[1264]$_SDFFE_PN0P__892  (.L_HI(net892));
 sg13g2_tiehi \shift_storage.storage[1265]$_SDFFE_PN0P__893  (.L_HI(net893));
 sg13g2_tiehi \shift_storage.storage[1266]$_SDFFE_PN0P__894  (.L_HI(net894));
 sg13g2_tiehi \shift_storage.storage[1267]$_SDFFE_PN0P__895  (.L_HI(net895));
 sg13g2_tiehi \shift_storage.storage[1268]$_SDFFE_PN0P__896  (.L_HI(net896));
 sg13g2_tiehi \shift_storage.storage[1269]$_SDFFE_PN0P__897  (.L_HI(net897));
 sg13g2_tiehi \shift_storage.storage[126]$_SDFFE_PN0P__898  (.L_HI(net898));
 sg13g2_tiehi \shift_storage.storage[1270]$_SDFFE_PN0P__899  (.L_HI(net899));
 sg13g2_tiehi \shift_storage.storage[1271]$_SDFFE_PN0P__900  (.L_HI(net900));
 sg13g2_tiehi \shift_storage.storage[1272]$_SDFFE_PN0P__901  (.L_HI(net901));
 sg13g2_tiehi \shift_storage.storage[1273]$_SDFFE_PN0P__902  (.L_HI(net902));
 sg13g2_tiehi \shift_storage.storage[1274]$_SDFFE_PN0P__903  (.L_HI(net903));
 sg13g2_tiehi \shift_storage.storage[1275]$_SDFFE_PN0P__904  (.L_HI(net904));
 sg13g2_tiehi \shift_storage.storage[1276]$_SDFFE_PN0P__905  (.L_HI(net905));
 sg13g2_tiehi \shift_storage.storage[1277]$_SDFFE_PN0P__906  (.L_HI(net906));
 sg13g2_tiehi \shift_storage.storage[1278]$_SDFFE_PN0P__907  (.L_HI(net907));
 sg13g2_tiehi \shift_storage.storage[1279]$_SDFFE_PN0P__908  (.L_HI(net908));
 sg13g2_tiehi \shift_storage.storage[127]$_SDFFE_PN0P__909  (.L_HI(net909));
 sg13g2_tiehi \shift_storage.storage[1280]$_SDFFE_PN0P__910  (.L_HI(net910));
 sg13g2_tiehi \shift_storage.storage[1281]$_SDFFE_PN0P__911  (.L_HI(net911));
 sg13g2_tiehi \shift_storage.storage[1282]$_SDFFE_PN0P__912  (.L_HI(net912));
 sg13g2_tiehi \shift_storage.storage[1283]$_SDFFE_PN0P__913  (.L_HI(net913));
 sg13g2_tiehi \shift_storage.storage[1284]$_SDFFE_PN0P__914  (.L_HI(net914));
 sg13g2_tiehi \shift_storage.storage[1285]$_SDFFE_PN0P__915  (.L_HI(net915));
 sg13g2_tiehi \shift_storage.storage[1286]$_SDFFE_PN0P__916  (.L_HI(net916));
 sg13g2_tiehi \shift_storage.storage[1287]$_SDFFE_PN0P__917  (.L_HI(net917));
 sg13g2_tiehi \shift_storage.storage[1288]$_SDFFE_PN0P__918  (.L_HI(net918));
 sg13g2_tiehi \shift_storage.storage[1289]$_SDFFE_PN0P__919  (.L_HI(net919));
 sg13g2_tiehi \shift_storage.storage[128]$_SDFFE_PN0P__920  (.L_HI(net920));
 sg13g2_tiehi \shift_storage.storage[1290]$_SDFFE_PN0P__921  (.L_HI(net921));
 sg13g2_tiehi \shift_storage.storage[1291]$_SDFFE_PN0P__922  (.L_HI(net922));
 sg13g2_tiehi \shift_storage.storage[1292]$_SDFFE_PN0P__923  (.L_HI(net923));
 sg13g2_tiehi \shift_storage.storage[1293]$_SDFFE_PN0P__924  (.L_HI(net924));
 sg13g2_tiehi \shift_storage.storage[1294]$_SDFFE_PN0P__925  (.L_HI(net925));
 sg13g2_tiehi \shift_storage.storage[1295]$_SDFFE_PN0P__926  (.L_HI(net926));
 sg13g2_tiehi \shift_storage.storage[1296]$_SDFFE_PN0P__927  (.L_HI(net927));
 sg13g2_tiehi \shift_storage.storage[1297]$_SDFFE_PN0P__928  (.L_HI(net928));
 sg13g2_tiehi \shift_storage.storage[1298]$_SDFFE_PN0P__929  (.L_HI(net929));
 sg13g2_tiehi \shift_storage.storage[1299]$_SDFFE_PN0P__930  (.L_HI(net930));
 sg13g2_tiehi \shift_storage.storage[129]$_SDFFE_PN0P__931  (.L_HI(net931));
 sg13g2_tiehi \shift_storage.storage[12]$_SDFFE_PN0P__932  (.L_HI(net932));
 sg13g2_tiehi \shift_storage.storage[1300]$_SDFFE_PN0P__933  (.L_HI(net933));
 sg13g2_tiehi \shift_storage.storage[1301]$_SDFFE_PN0P__934  (.L_HI(net934));
 sg13g2_tiehi \shift_storage.storage[1302]$_SDFFE_PN0P__935  (.L_HI(net935));
 sg13g2_tiehi \shift_storage.storage[1303]$_SDFFE_PN0P__936  (.L_HI(net936));
 sg13g2_tiehi \shift_storage.storage[1304]$_SDFFE_PN0P__937  (.L_HI(net937));
 sg13g2_tiehi \shift_storage.storage[1305]$_SDFFE_PN0P__938  (.L_HI(net938));
 sg13g2_tiehi \shift_storage.storage[1306]$_SDFFE_PN0P__939  (.L_HI(net939));
 sg13g2_tiehi \shift_storage.storage[1307]$_SDFFE_PN0P__940  (.L_HI(net940));
 sg13g2_tiehi \shift_storage.storage[1308]$_SDFFE_PN0P__941  (.L_HI(net941));
 sg13g2_tiehi \shift_storage.storage[1309]$_SDFFE_PN0P__942  (.L_HI(net942));
 sg13g2_tiehi \shift_storage.storage[130]$_SDFFE_PN0P__943  (.L_HI(net943));
 sg13g2_tiehi \shift_storage.storage[1310]$_SDFFE_PN0P__944  (.L_HI(net944));
 sg13g2_tiehi \shift_storage.storage[1311]$_SDFFE_PN0P__945  (.L_HI(net945));
 sg13g2_tiehi \shift_storage.storage[1312]$_SDFFE_PN0P__946  (.L_HI(net946));
 sg13g2_tiehi \shift_storage.storage[1313]$_SDFFE_PN0P__947  (.L_HI(net947));
 sg13g2_tiehi \shift_storage.storage[1314]$_SDFFE_PN0P__948  (.L_HI(net948));
 sg13g2_tiehi \shift_storage.storage[1315]$_SDFFE_PN0P__949  (.L_HI(net949));
 sg13g2_tiehi \shift_storage.storage[1316]$_SDFFE_PN0P__950  (.L_HI(net950));
 sg13g2_tiehi \shift_storage.storage[1317]$_SDFFE_PN0P__951  (.L_HI(net951));
 sg13g2_tiehi \shift_storage.storage[1318]$_SDFFE_PN0P__952  (.L_HI(net952));
 sg13g2_tiehi \shift_storage.storage[1319]$_SDFFE_PN0P__953  (.L_HI(net953));
 sg13g2_tiehi \shift_storage.storage[131]$_SDFFE_PN0P__954  (.L_HI(net954));
 sg13g2_tiehi \shift_storage.storage[1320]$_SDFFE_PN0P__955  (.L_HI(net955));
 sg13g2_tiehi \shift_storage.storage[1321]$_SDFFE_PN0P__956  (.L_HI(net956));
 sg13g2_tiehi \shift_storage.storage[1322]$_SDFFE_PN0P__957  (.L_HI(net957));
 sg13g2_tiehi \shift_storage.storage[1323]$_SDFFE_PN0P__958  (.L_HI(net958));
 sg13g2_tiehi \shift_storage.storage[1324]$_SDFFE_PN0P__959  (.L_HI(net959));
 sg13g2_tiehi \shift_storage.storage[1325]$_SDFFE_PN0P__960  (.L_HI(net960));
 sg13g2_tiehi \shift_storage.storage[1326]$_SDFFE_PN0P__961  (.L_HI(net961));
 sg13g2_tiehi \shift_storage.storage[1327]$_SDFFE_PN0P__962  (.L_HI(net962));
 sg13g2_tiehi \shift_storage.storage[1328]$_SDFFE_PN0P__963  (.L_HI(net963));
 sg13g2_tiehi \shift_storage.storage[1329]$_SDFFE_PN0P__964  (.L_HI(net964));
 sg13g2_tiehi \shift_storage.storage[132]$_SDFFE_PN0P__965  (.L_HI(net965));
 sg13g2_tiehi \shift_storage.storage[1330]$_SDFFE_PN0P__966  (.L_HI(net966));
 sg13g2_tiehi \shift_storage.storage[1331]$_SDFFE_PN0P__967  (.L_HI(net967));
 sg13g2_tiehi \shift_storage.storage[1332]$_SDFFE_PN0P__968  (.L_HI(net968));
 sg13g2_tiehi \shift_storage.storage[1333]$_SDFFE_PN0P__969  (.L_HI(net969));
 sg13g2_tiehi \shift_storage.storage[1334]$_SDFFE_PN0P__970  (.L_HI(net970));
 sg13g2_tiehi \shift_storage.storage[1335]$_SDFFE_PN0P__971  (.L_HI(net971));
 sg13g2_tiehi \shift_storage.storage[1336]$_SDFFE_PN0P__972  (.L_HI(net972));
 sg13g2_tiehi \shift_storage.storage[1337]$_SDFFE_PN0P__973  (.L_HI(net973));
 sg13g2_tiehi \shift_storage.storage[1338]$_SDFFE_PN0P__974  (.L_HI(net974));
 sg13g2_tiehi \shift_storage.storage[1339]$_SDFFE_PN0P__975  (.L_HI(net975));
 sg13g2_tiehi \shift_storage.storage[133]$_SDFFE_PN0P__976  (.L_HI(net976));
 sg13g2_tiehi \shift_storage.storage[1340]$_SDFFE_PN0P__977  (.L_HI(net977));
 sg13g2_tiehi \shift_storage.storage[1341]$_SDFFE_PN0P__978  (.L_HI(net978));
 sg13g2_tiehi \shift_storage.storage[1342]$_SDFFE_PN0P__979  (.L_HI(net979));
 sg13g2_tiehi \shift_storage.storage[1343]$_SDFFE_PN0P__980  (.L_HI(net980));
 sg13g2_tiehi \shift_storage.storage[1344]$_SDFFE_PN0P__981  (.L_HI(net981));
 sg13g2_tiehi \shift_storage.storage[1345]$_SDFFE_PN0P__982  (.L_HI(net982));
 sg13g2_tiehi \shift_storage.storage[1346]$_SDFFE_PN0P__983  (.L_HI(net983));
 sg13g2_tiehi \shift_storage.storage[1347]$_SDFFE_PN0P__984  (.L_HI(net984));
 sg13g2_tiehi \shift_storage.storage[1348]$_SDFFE_PN0P__985  (.L_HI(net985));
 sg13g2_tiehi \shift_storage.storage[1349]$_SDFFE_PN0P__986  (.L_HI(net986));
 sg13g2_tiehi \shift_storage.storage[134]$_SDFFE_PN0P__987  (.L_HI(net987));
 sg13g2_tiehi \shift_storage.storage[1350]$_SDFFE_PN0P__988  (.L_HI(net988));
 sg13g2_tiehi \shift_storage.storage[1351]$_SDFFE_PN0P__989  (.L_HI(net989));
 sg13g2_tiehi \shift_storage.storage[1352]$_SDFFE_PN0P__990  (.L_HI(net990));
 sg13g2_tiehi \shift_storage.storage[1353]$_SDFFE_PN0P__991  (.L_HI(net991));
 sg13g2_tiehi \shift_storage.storage[1354]$_SDFFE_PN0P__992  (.L_HI(net992));
 sg13g2_tiehi \shift_storage.storage[1355]$_SDFFE_PN0P__993  (.L_HI(net993));
 sg13g2_tiehi \shift_storage.storage[1356]$_SDFFE_PN0P__994  (.L_HI(net994));
 sg13g2_tiehi \shift_storage.storage[1357]$_SDFFE_PN0P__995  (.L_HI(net995));
 sg13g2_tiehi \shift_storage.storage[1358]$_SDFFE_PN0P__996  (.L_HI(net996));
 sg13g2_tiehi \shift_storage.storage[1359]$_SDFFE_PN0P__997  (.L_HI(net997));
 sg13g2_tiehi \shift_storage.storage[135]$_SDFFE_PN0P__998  (.L_HI(net998));
 sg13g2_tiehi \shift_storage.storage[1360]$_SDFFE_PN0P__999  (.L_HI(net999));
 sg13g2_tiehi \shift_storage.storage[1361]$_SDFFE_PN0P__1000  (.L_HI(net1000));
 sg13g2_tiehi \shift_storage.storage[1362]$_SDFFE_PN0P__1001  (.L_HI(net1001));
 sg13g2_tiehi \shift_storage.storage[1363]$_SDFFE_PN0P__1002  (.L_HI(net1002));
 sg13g2_tiehi \shift_storage.storage[1364]$_SDFFE_PN0P__1003  (.L_HI(net1003));
 sg13g2_tiehi \shift_storage.storage[1365]$_SDFFE_PN0P__1004  (.L_HI(net1004));
 sg13g2_tiehi \shift_storage.storage[1366]$_SDFFE_PN0P__1005  (.L_HI(net1005));
 sg13g2_tiehi \shift_storage.storage[1367]$_SDFFE_PN0P__1006  (.L_HI(net1006));
 sg13g2_tiehi \shift_storage.storage[1368]$_SDFFE_PN0P__1007  (.L_HI(net1007));
 sg13g2_tiehi \shift_storage.storage[1369]$_SDFFE_PN0P__1008  (.L_HI(net1008));
 sg13g2_tiehi \shift_storage.storage[136]$_SDFFE_PN0P__1009  (.L_HI(net1009));
 sg13g2_tiehi \shift_storage.storage[1370]$_SDFFE_PN0P__1010  (.L_HI(net1010));
 sg13g2_tiehi \shift_storage.storage[1371]$_SDFFE_PN0P__1011  (.L_HI(net1011));
 sg13g2_tiehi \shift_storage.storage[1372]$_SDFFE_PN0P__1012  (.L_HI(net1012));
 sg13g2_tiehi \shift_storage.storage[1373]$_SDFFE_PN0P__1013  (.L_HI(net1013));
 sg13g2_tiehi \shift_storage.storage[1374]$_SDFFE_PN0P__1014  (.L_HI(net1014));
 sg13g2_tiehi \shift_storage.storage[1375]$_SDFFE_PN0P__1015  (.L_HI(net1015));
 sg13g2_tiehi \shift_storage.storage[1376]$_SDFFE_PN0P__1016  (.L_HI(net1016));
 sg13g2_tiehi \shift_storage.storage[1377]$_SDFFE_PN0P__1017  (.L_HI(net1017));
 sg13g2_tiehi \shift_storage.storage[1378]$_SDFFE_PN0P__1018  (.L_HI(net1018));
 sg13g2_tiehi \shift_storage.storage[1379]$_SDFFE_PN0P__1019  (.L_HI(net1019));
 sg13g2_tiehi \shift_storage.storage[137]$_SDFFE_PN0P__1020  (.L_HI(net1020));
 sg13g2_tiehi \shift_storage.storage[1380]$_SDFFE_PN0P__1021  (.L_HI(net1021));
 sg13g2_tiehi \shift_storage.storage[1381]$_SDFFE_PN0P__1022  (.L_HI(net1022));
 sg13g2_tiehi \shift_storage.storage[1382]$_SDFFE_PN0P__1023  (.L_HI(net1023));
 sg13g2_tiehi \shift_storage.storage[1383]$_SDFFE_PN0P__1024  (.L_HI(net1024));
 sg13g2_tiehi \shift_storage.storage[1384]$_SDFFE_PN0P__1025  (.L_HI(net1025));
 sg13g2_tiehi \shift_storage.storage[1385]$_SDFFE_PN0P__1026  (.L_HI(net1026));
 sg13g2_tiehi \shift_storage.storage[1386]$_SDFFE_PN0P__1027  (.L_HI(net1027));
 sg13g2_tiehi \shift_storage.storage[1387]$_SDFFE_PN0P__1028  (.L_HI(net1028));
 sg13g2_tiehi \shift_storage.storage[1388]$_SDFFE_PN0P__1029  (.L_HI(net1029));
 sg13g2_tiehi \shift_storage.storage[1389]$_SDFFE_PN0P__1030  (.L_HI(net1030));
 sg13g2_tiehi \shift_storage.storage[138]$_SDFFE_PN0P__1031  (.L_HI(net1031));
 sg13g2_tiehi \shift_storage.storage[1390]$_SDFFE_PN0P__1032  (.L_HI(net1032));
 sg13g2_tiehi \shift_storage.storage[1391]$_SDFFE_PN0P__1033  (.L_HI(net1033));
 sg13g2_tiehi \shift_storage.storage[1392]$_SDFFE_PN0P__1034  (.L_HI(net1034));
 sg13g2_tiehi \shift_storage.storage[1393]$_SDFFE_PN0P__1035  (.L_HI(net1035));
 sg13g2_tiehi \shift_storage.storage[1394]$_SDFFE_PN0P__1036  (.L_HI(net1036));
 sg13g2_tiehi \shift_storage.storage[1395]$_SDFFE_PN0P__1037  (.L_HI(net1037));
 sg13g2_tiehi \shift_storage.storage[1396]$_SDFFE_PN0P__1038  (.L_HI(net1038));
 sg13g2_tiehi \shift_storage.storage[1397]$_SDFFE_PN0P__1039  (.L_HI(net1039));
 sg13g2_tiehi \shift_storage.storage[1398]$_SDFFE_PN0P__1040  (.L_HI(net1040));
 sg13g2_tiehi \shift_storage.storage[1399]$_SDFFE_PN0P__1041  (.L_HI(net1041));
 sg13g2_tiehi \shift_storage.storage[139]$_SDFFE_PN0P__1042  (.L_HI(net1042));
 sg13g2_tiehi \shift_storage.storage[13]$_SDFFE_PN0P__1043  (.L_HI(net1043));
 sg13g2_tiehi \shift_storage.storage[1400]$_SDFFE_PN0P__1044  (.L_HI(net1044));
 sg13g2_tiehi \shift_storage.storage[1401]$_SDFFE_PN0P__1045  (.L_HI(net1045));
 sg13g2_tiehi \shift_storage.storage[1402]$_SDFFE_PN0P__1046  (.L_HI(net1046));
 sg13g2_tiehi \shift_storage.storage[1403]$_SDFFE_PN0P__1047  (.L_HI(net1047));
 sg13g2_tiehi \shift_storage.storage[1404]$_SDFFE_PN0P__1048  (.L_HI(net1048));
 sg13g2_tiehi \shift_storage.storage[1405]$_SDFFE_PN0P__1049  (.L_HI(net1049));
 sg13g2_tiehi \shift_storage.storage[1406]$_SDFFE_PN0P__1050  (.L_HI(net1050));
 sg13g2_tiehi \shift_storage.storage[1407]$_SDFFE_PN0P__1051  (.L_HI(net1051));
 sg13g2_tiehi \shift_storage.storage[1408]$_SDFFE_PN0P__1052  (.L_HI(net1052));
 sg13g2_tiehi \shift_storage.storage[1409]$_SDFFE_PN0P__1053  (.L_HI(net1053));
 sg13g2_tiehi \shift_storage.storage[140]$_SDFFE_PN0P__1054  (.L_HI(net1054));
 sg13g2_tiehi \shift_storage.storage[1410]$_SDFFE_PN0P__1055  (.L_HI(net1055));
 sg13g2_tiehi \shift_storage.storage[1411]$_SDFFE_PN0P__1056  (.L_HI(net1056));
 sg13g2_tiehi \shift_storage.storage[1412]$_SDFFE_PN0P__1057  (.L_HI(net1057));
 sg13g2_tiehi \shift_storage.storage[1413]$_SDFFE_PN0P__1058  (.L_HI(net1058));
 sg13g2_tiehi \shift_storage.storage[1414]$_SDFFE_PN0P__1059  (.L_HI(net1059));
 sg13g2_tiehi \shift_storage.storage[1415]$_SDFFE_PN0P__1060  (.L_HI(net1060));
 sg13g2_tiehi \shift_storage.storage[1416]$_SDFFE_PN0P__1061  (.L_HI(net1061));
 sg13g2_tiehi \shift_storage.storage[1417]$_SDFFE_PN0P__1062  (.L_HI(net1062));
 sg13g2_tiehi \shift_storage.storage[1418]$_SDFFE_PN0P__1063  (.L_HI(net1063));
 sg13g2_tiehi \shift_storage.storage[1419]$_SDFFE_PN0P__1064  (.L_HI(net1064));
 sg13g2_tiehi \shift_storage.storage[141]$_SDFFE_PN0P__1065  (.L_HI(net1065));
 sg13g2_tiehi \shift_storage.storage[1420]$_SDFFE_PN0P__1066  (.L_HI(net1066));
 sg13g2_tiehi \shift_storage.storage[1421]$_SDFFE_PN0P__1067  (.L_HI(net1067));
 sg13g2_tiehi \shift_storage.storage[1422]$_SDFFE_PN0P__1068  (.L_HI(net1068));
 sg13g2_tiehi \shift_storage.storage[1423]$_SDFFE_PN0P__1069  (.L_HI(net1069));
 sg13g2_tiehi \shift_storage.storage[1424]$_SDFFE_PN0P__1070  (.L_HI(net1070));
 sg13g2_tiehi \shift_storage.storage[1425]$_SDFFE_PN0P__1071  (.L_HI(net1071));
 sg13g2_tiehi \shift_storage.storage[1426]$_SDFFE_PN0P__1072  (.L_HI(net1072));
 sg13g2_tiehi \shift_storage.storage[1427]$_SDFFE_PN0P__1073  (.L_HI(net1073));
 sg13g2_tiehi \shift_storage.storage[1428]$_SDFFE_PN0P__1074  (.L_HI(net1074));
 sg13g2_tiehi \shift_storage.storage[1429]$_SDFFE_PN0P__1075  (.L_HI(net1075));
 sg13g2_tiehi \shift_storage.storage[142]$_SDFFE_PN0P__1076  (.L_HI(net1076));
 sg13g2_tiehi \shift_storage.storage[1430]$_SDFFE_PN0P__1077  (.L_HI(net1077));
 sg13g2_tiehi \shift_storage.storage[1431]$_SDFFE_PN0P__1078  (.L_HI(net1078));
 sg13g2_tiehi \shift_storage.storage[1432]$_SDFFE_PN0P__1079  (.L_HI(net1079));
 sg13g2_tiehi \shift_storage.storage[1433]$_SDFFE_PN0P__1080  (.L_HI(net1080));
 sg13g2_tiehi \shift_storage.storage[1434]$_SDFFE_PN0P__1081  (.L_HI(net1081));
 sg13g2_tiehi \shift_storage.storage[1435]$_SDFFE_PN0P__1082  (.L_HI(net1082));
 sg13g2_tiehi \shift_storage.storage[1436]$_SDFFE_PN0P__1083  (.L_HI(net1083));
 sg13g2_tiehi \shift_storage.storage[1437]$_SDFFE_PN0P__1084  (.L_HI(net1084));
 sg13g2_tiehi \shift_storage.storage[1438]$_SDFFE_PN0P__1085  (.L_HI(net1085));
 sg13g2_tiehi \shift_storage.storage[1439]$_SDFFE_PN0P__1086  (.L_HI(net1086));
 sg13g2_tiehi \shift_storage.storage[143]$_SDFFE_PN0P__1087  (.L_HI(net1087));
 sg13g2_tiehi \shift_storage.storage[1440]$_SDFFE_PN0P__1088  (.L_HI(net1088));
 sg13g2_tiehi \shift_storage.storage[1441]$_SDFFE_PN0P__1089  (.L_HI(net1089));
 sg13g2_tiehi \shift_storage.storage[1442]$_SDFFE_PN0P__1090  (.L_HI(net1090));
 sg13g2_tiehi \shift_storage.storage[1443]$_SDFFE_PN0P__1091  (.L_HI(net1091));
 sg13g2_tiehi \shift_storage.storage[1444]$_SDFFE_PN0P__1092  (.L_HI(net1092));
 sg13g2_tiehi \shift_storage.storage[1445]$_SDFFE_PN0P__1093  (.L_HI(net1093));
 sg13g2_tiehi \shift_storage.storage[1446]$_SDFFE_PN0P__1094  (.L_HI(net1094));
 sg13g2_tiehi \shift_storage.storage[1447]$_SDFFE_PN0P__1095  (.L_HI(net1095));
 sg13g2_tiehi \shift_storage.storage[1448]$_SDFFE_PN0P__1096  (.L_HI(net1096));
 sg13g2_tiehi \shift_storage.storage[1449]$_SDFFE_PN0P__1097  (.L_HI(net1097));
 sg13g2_tiehi \shift_storage.storage[144]$_SDFFE_PN0P__1098  (.L_HI(net1098));
 sg13g2_tiehi \shift_storage.storage[1450]$_SDFFE_PN0P__1099  (.L_HI(net1099));
 sg13g2_tiehi \shift_storage.storage[1451]$_SDFFE_PN0P__1100  (.L_HI(net1100));
 sg13g2_tiehi \shift_storage.storage[1452]$_SDFFE_PN0P__1101  (.L_HI(net1101));
 sg13g2_tiehi \shift_storage.storage[1453]$_SDFFE_PN0P__1102  (.L_HI(net1102));
 sg13g2_tiehi \shift_storage.storage[1454]$_SDFFE_PN0P__1103  (.L_HI(net1103));
 sg13g2_tiehi \shift_storage.storage[1455]$_SDFFE_PN0P__1104  (.L_HI(net1104));
 sg13g2_tiehi \shift_storage.storage[1456]$_SDFFE_PN0P__1105  (.L_HI(net1105));
 sg13g2_tiehi \shift_storage.storage[1457]$_SDFFE_PN0P__1106  (.L_HI(net1106));
 sg13g2_tiehi \shift_storage.storage[1458]$_SDFFE_PN0P__1107  (.L_HI(net1107));
 sg13g2_tiehi \shift_storage.storage[1459]$_SDFFE_PN0P__1108  (.L_HI(net1108));
 sg13g2_tiehi \shift_storage.storage[145]$_SDFFE_PN0P__1109  (.L_HI(net1109));
 sg13g2_tiehi \shift_storage.storage[1460]$_SDFFE_PN0P__1110  (.L_HI(net1110));
 sg13g2_tiehi \shift_storage.storage[1461]$_SDFFE_PN0P__1111  (.L_HI(net1111));
 sg13g2_tiehi \shift_storage.storage[1462]$_SDFFE_PN0P__1112  (.L_HI(net1112));
 sg13g2_tiehi \shift_storage.storage[1463]$_SDFFE_PN0P__1113  (.L_HI(net1113));
 sg13g2_tiehi \shift_storage.storage[1464]$_SDFFE_PN0P__1114  (.L_HI(net1114));
 sg13g2_tiehi \shift_storage.storage[1465]$_SDFFE_PN0P__1115  (.L_HI(net1115));
 sg13g2_tiehi \shift_storage.storage[1466]$_SDFFE_PN0P__1116  (.L_HI(net1116));
 sg13g2_tiehi \shift_storage.storage[1467]$_SDFFE_PN0P__1117  (.L_HI(net1117));
 sg13g2_tiehi \shift_storage.storage[1468]$_SDFFE_PN0P__1118  (.L_HI(net1118));
 sg13g2_tiehi \shift_storage.storage[1469]$_SDFFE_PN0P__1119  (.L_HI(net1119));
 sg13g2_tiehi \shift_storage.storage[146]$_SDFFE_PN0P__1120  (.L_HI(net1120));
 sg13g2_tiehi \shift_storage.storage[1470]$_SDFFE_PN0P__1121  (.L_HI(net1121));
 sg13g2_tiehi \shift_storage.storage[1471]$_SDFFE_PN0P__1122  (.L_HI(net1122));
 sg13g2_tiehi \shift_storage.storage[1472]$_SDFFE_PN0P__1123  (.L_HI(net1123));
 sg13g2_tiehi \shift_storage.storage[1473]$_SDFFE_PN0P__1124  (.L_HI(net1124));
 sg13g2_tiehi \shift_storage.storage[1474]$_SDFFE_PN0P__1125  (.L_HI(net1125));
 sg13g2_tiehi \shift_storage.storage[1475]$_SDFFE_PN0P__1126  (.L_HI(net1126));
 sg13g2_tiehi \shift_storage.storage[1476]$_SDFFE_PN0P__1127  (.L_HI(net1127));
 sg13g2_tiehi \shift_storage.storage[1477]$_SDFFE_PN0P__1128  (.L_HI(net1128));
 sg13g2_tiehi \shift_storage.storage[1478]$_SDFFE_PN0P__1129  (.L_HI(net1129));
 sg13g2_tiehi \shift_storage.storage[1479]$_SDFFE_PN0P__1130  (.L_HI(net1130));
 sg13g2_tiehi \shift_storage.storage[147]$_SDFFE_PN0P__1131  (.L_HI(net1131));
 sg13g2_tiehi \shift_storage.storage[1480]$_SDFFE_PN0P__1132  (.L_HI(net1132));
 sg13g2_tiehi \shift_storage.storage[1481]$_SDFFE_PN0P__1133  (.L_HI(net1133));
 sg13g2_tiehi \shift_storage.storage[1482]$_SDFFE_PN0P__1134  (.L_HI(net1134));
 sg13g2_tiehi \shift_storage.storage[1483]$_SDFFE_PN0P__1135  (.L_HI(net1135));
 sg13g2_tiehi \shift_storage.storage[1484]$_SDFFE_PN0P__1136  (.L_HI(net1136));
 sg13g2_tiehi \shift_storage.storage[1485]$_SDFFE_PN0P__1137  (.L_HI(net1137));
 sg13g2_tiehi \shift_storage.storage[1486]$_SDFFE_PN0P__1138  (.L_HI(net1138));
 sg13g2_tiehi \shift_storage.storage[1487]$_SDFFE_PN0P__1139  (.L_HI(net1139));
 sg13g2_tiehi \shift_storage.storage[1488]$_SDFFE_PN0P__1140  (.L_HI(net1140));
 sg13g2_tiehi \shift_storage.storage[1489]$_SDFFE_PN0P__1141  (.L_HI(net1141));
 sg13g2_tiehi \shift_storage.storage[148]$_SDFFE_PN0P__1142  (.L_HI(net1142));
 sg13g2_tiehi \shift_storage.storage[1490]$_SDFFE_PN0P__1143  (.L_HI(net1143));
 sg13g2_tiehi \shift_storage.storage[1491]$_SDFFE_PN0P__1144  (.L_HI(net1144));
 sg13g2_tiehi \shift_storage.storage[1492]$_SDFFE_PN0P__1145  (.L_HI(net1145));
 sg13g2_tiehi \shift_storage.storage[1493]$_SDFFE_PN0P__1146  (.L_HI(net1146));
 sg13g2_tiehi \shift_storage.storage[1494]$_SDFFE_PN0P__1147  (.L_HI(net1147));
 sg13g2_tiehi \shift_storage.storage[1495]$_SDFFE_PN0P__1148  (.L_HI(net1148));
 sg13g2_tiehi \shift_storage.storage[1496]$_SDFFE_PN0P__1149  (.L_HI(net1149));
 sg13g2_tiehi \shift_storage.storage[1497]$_SDFFE_PN0P__1150  (.L_HI(net1150));
 sg13g2_tiehi \shift_storage.storage[1498]$_SDFFE_PN0P__1151  (.L_HI(net1151));
 sg13g2_tiehi \shift_storage.storage[1499]$_SDFFE_PN0P__1152  (.L_HI(net1152));
 sg13g2_tiehi \shift_storage.storage[149]$_SDFFE_PN0P__1153  (.L_HI(net1153));
 sg13g2_tiehi \shift_storage.storage[14]$_SDFFE_PN0P__1154  (.L_HI(net1154));
 sg13g2_tiehi \shift_storage.storage[1500]$_SDFFE_PN0P__1155  (.L_HI(net1155));
 sg13g2_tiehi \shift_storage.storage[1501]$_SDFFE_PN0P__1156  (.L_HI(net1156));
 sg13g2_tiehi \shift_storage.storage[1502]$_SDFFE_PN0P__1157  (.L_HI(net1157));
 sg13g2_tiehi \shift_storage.storage[1503]$_SDFFE_PN0P__1158  (.L_HI(net1158));
 sg13g2_tiehi \shift_storage.storage[1504]$_SDFFE_PN0P__1159  (.L_HI(net1159));
 sg13g2_tiehi \shift_storage.storage[1505]$_SDFFE_PN0P__1160  (.L_HI(net1160));
 sg13g2_tiehi \shift_storage.storage[1506]$_SDFFE_PN0P__1161  (.L_HI(net1161));
 sg13g2_tiehi \shift_storage.storage[1507]$_SDFFE_PN0P__1162  (.L_HI(net1162));
 sg13g2_tiehi \shift_storage.storage[1508]$_SDFFE_PN0P__1163  (.L_HI(net1163));
 sg13g2_tiehi \shift_storage.storage[1509]$_SDFFE_PN0P__1164  (.L_HI(net1164));
 sg13g2_tiehi \shift_storage.storage[150]$_SDFFE_PN0P__1165  (.L_HI(net1165));
 sg13g2_tiehi \shift_storage.storage[1510]$_SDFFE_PN0P__1166  (.L_HI(net1166));
 sg13g2_tiehi \shift_storage.storage[1511]$_SDFFE_PN0P__1167  (.L_HI(net1167));
 sg13g2_tiehi \shift_storage.storage[1512]$_SDFFE_PN0P__1168  (.L_HI(net1168));
 sg13g2_tiehi \shift_storage.storage[1513]$_SDFFE_PN0P__1169  (.L_HI(net1169));
 sg13g2_tiehi \shift_storage.storage[1514]$_SDFFE_PN0P__1170  (.L_HI(net1170));
 sg13g2_tiehi \shift_storage.storage[1515]$_SDFFE_PN0P__1171  (.L_HI(net1171));
 sg13g2_tiehi \shift_storage.storage[1516]$_SDFFE_PN0P__1172  (.L_HI(net1172));
 sg13g2_tiehi \shift_storage.storage[1517]$_SDFFE_PN0P__1173  (.L_HI(net1173));
 sg13g2_tiehi \shift_storage.storage[1518]$_SDFFE_PN0P__1174  (.L_HI(net1174));
 sg13g2_tiehi \shift_storage.storage[1519]$_SDFFE_PN0P__1175  (.L_HI(net1175));
 sg13g2_tiehi \shift_storage.storage[151]$_SDFFE_PN0P__1176  (.L_HI(net1176));
 sg13g2_tiehi \shift_storage.storage[1520]$_SDFFE_PN0P__1177  (.L_HI(net1177));
 sg13g2_tiehi \shift_storage.storage[1521]$_SDFFE_PN0P__1178  (.L_HI(net1178));
 sg13g2_tiehi \shift_storage.storage[1522]$_SDFFE_PN0P__1179  (.L_HI(net1179));
 sg13g2_tiehi \shift_storage.storage[1523]$_SDFFE_PN0P__1180  (.L_HI(net1180));
 sg13g2_tiehi \shift_storage.storage[1524]$_SDFFE_PN0P__1181  (.L_HI(net1181));
 sg13g2_tiehi \shift_storage.storage[1525]$_SDFFE_PN0P__1182  (.L_HI(net1182));
 sg13g2_tiehi \shift_storage.storage[1526]$_SDFFE_PN0P__1183  (.L_HI(net1183));
 sg13g2_tiehi \shift_storage.storage[1527]$_SDFFE_PN0P__1184  (.L_HI(net1184));
 sg13g2_tiehi \shift_storage.storage[1528]$_SDFFE_PN0P__1185  (.L_HI(net1185));
 sg13g2_tiehi \shift_storage.storage[1529]$_SDFFE_PN0P__1186  (.L_HI(net1186));
 sg13g2_tiehi \shift_storage.storage[152]$_SDFFE_PN0P__1187  (.L_HI(net1187));
 sg13g2_tiehi \shift_storage.storage[1530]$_SDFFE_PN0P__1188  (.L_HI(net1188));
 sg13g2_tiehi \shift_storage.storage[1531]$_SDFFE_PN0P__1189  (.L_HI(net1189));
 sg13g2_tiehi \shift_storage.storage[1532]$_SDFFE_PN0P__1190  (.L_HI(net1190));
 sg13g2_tiehi \shift_storage.storage[1533]$_SDFFE_PN0P__1191  (.L_HI(net1191));
 sg13g2_tiehi \shift_storage.storage[1534]$_SDFFE_PN0P__1192  (.L_HI(net1192));
 sg13g2_tiehi \shift_storage.storage[1535]$_SDFFE_PN0P__1193  (.L_HI(net1193));
 sg13g2_tiehi \shift_storage.storage[1536]$_SDFFE_PN0P__1194  (.L_HI(net1194));
 sg13g2_tiehi \shift_storage.storage[1537]$_SDFFE_PN0P__1195  (.L_HI(net1195));
 sg13g2_tiehi \shift_storage.storage[1538]$_SDFFE_PN0P__1196  (.L_HI(net1196));
 sg13g2_tiehi \shift_storage.storage[1539]$_SDFFE_PN0P__1197  (.L_HI(net1197));
 sg13g2_tiehi \shift_storage.storage[153]$_SDFFE_PN0P__1198  (.L_HI(net1198));
 sg13g2_tiehi \shift_storage.storage[1540]$_SDFFE_PN0P__1199  (.L_HI(net1199));
 sg13g2_tiehi \shift_storage.storage[1541]$_SDFFE_PN0P__1200  (.L_HI(net1200));
 sg13g2_tiehi \shift_storage.storage[1542]$_SDFFE_PN0P__1201  (.L_HI(net1201));
 sg13g2_tiehi \shift_storage.storage[1543]$_SDFFE_PN0P__1202  (.L_HI(net1202));
 sg13g2_tiehi \shift_storage.storage[1544]$_SDFFE_PN0P__1203  (.L_HI(net1203));
 sg13g2_tiehi \shift_storage.storage[1545]$_SDFFE_PN0P__1204  (.L_HI(net1204));
 sg13g2_tiehi \shift_storage.storage[1546]$_SDFFE_PN0P__1205  (.L_HI(net1205));
 sg13g2_tiehi \shift_storage.storage[1547]$_SDFFE_PN0P__1206  (.L_HI(net1206));
 sg13g2_tiehi \shift_storage.storage[1548]$_SDFFE_PN0P__1207  (.L_HI(net1207));
 sg13g2_tiehi \shift_storage.storage[1549]$_SDFFE_PN0P__1208  (.L_HI(net1208));
 sg13g2_tiehi \shift_storage.storage[154]$_SDFFE_PN0P__1209  (.L_HI(net1209));
 sg13g2_tiehi \shift_storage.storage[1550]$_SDFFE_PN0P__1210  (.L_HI(net1210));
 sg13g2_tiehi \shift_storage.storage[1551]$_SDFFE_PN0P__1211  (.L_HI(net1211));
 sg13g2_tiehi \shift_storage.storage[1552]$_SDFFE_PN0P__1212  (.L_HI(net1212));
 sg13g2_tiehi \shift_storage.storage[1553]$_SDFFE_PN0P__1213  (.L_HI(net1213));
 sg13g2_tiehi \shift_storage.storage[1554]$_SDFFE_PN0P__1214  (.L_HI(net1214));
 sg13g2_tiehi \shift_storage.storage[1555]$_SDFFE_PN0P__1215  (.L_HI(net1215));
 sg13g2_tiehi \shift_storage.storage[1556]$_SDFFE_PN0P__1216  (.L_HI(net1216));
 sg13g2_tiehi \shift_storage.storage[1557]$_SDFFE_PN0P__1217  (.L_HI(net1217));
 sg13g2_tiehi \shift_storage.storage[1558]$_SDFFE_PN0P__1218  (.L_HI(net1218));
 sg13g2_tiehi \shift_storage.storage[1559]$_SDFFE_PN0P__1219  (.L_HI(net1219));
 sg13g2_tiehi \shift_storage.storage[155]$_SDFFE_PN0P__1220  (.L_HI(net1220));
 sg13g2_tiehi \shift_storage.storage[1560]$_SDFFE_PN0P__1221  (.L_HI(net1221));
 sg13g2_tiehi \shift_storage.storage[1561]$_SDFFE_PN0P__1222  (.L_HI(net1222));
 sg13g2_tiehi \shift_storage.storage[1562]$_SDFFE_PN0P__1223  (.L_HI(net1223));
 sg13g2_tiehi \shift_storage.storage[1563]$_SDFFE_PN0P__1224  (.L_HI(net1224));
 sg13g2_tiehi \shift_storage.storage[1564]$_SDFFE_PN0P__1225  (.L_HI(net1225));
 sg13g2_tiehi \shift_storage.storage[1565]$_SDFFE_PN0P__1226  (.L_HI(net1226));
 sg13g2_tiehi \shift_storage.storage[1566]$_SDFFE_PN0P__1227  (.L_HI(net1227));
 sg13g2_tiehi \shift_storage.storage[1567]$_SDFFE_PN0P__1228  (.L_HI(net1228));
 sg13g2_tiehi \shift_storage.storage[1568]$_SDFFE_PN0P__1229  (.L_HI(net1229));
 sg13g2_tiehi \shift_storage.storage[1569]$_SDFFE_PN0P__1230  (.L_HI(net1230));
 sg13g2_tiehi \shift_storage.storage[156]$_SDFFE_PN0P__1231  (.L_HI(net1231));
 sg13g2_tiehi \shift_storage.storage[1570]$_SDFFE_PN0P__1232  (.L_HI(net1232));
 sg13g2_tiehi \shift_storage.storage[1571]$_SDFFE_PN0P__1233  (.L_HI(net1233));
 sg13g2_tiehi \shift_storage.storage[1572]$_SDFFE_PN0P__1234  (.L_HI(net1234));
 sg13g2_tiehi \shift_storage.storage[1573]$_SDFFE_PN0P__1235  (.L_HI(net1235));
 sg13g2_tiehi \shift_storage.storage[1574]$_SDFFE_PN0P__1236  (.L_HI(net1236));
 sg13g2_tiehi \shift_storage.storage[1575]$_SDFFE_PN0P__1237  (.L_HI(net1237));
 sg13g2_tiehi \shift_storage.storage[1576]$_SDFFE_PN0P__1238  (.L_HI(net1238));
 sg13g2_tiehi \shift_storage.storage[1577]$_SDFFE_PN0P__1239  (.L_HI(net1239));
 sg13g2_tiehi \shift_storage.storage[1578]$_SDFFE_PN0P__1240  (.L_HI(net1240));
 sg13g2_tiehi \shift_storage.storage[1579]$_SDFFE_PN0P__1241  (.L_HI(net1241));
 sg13g2_tiehi \shift_storage.storage[157]$_SDFFE_PN0P__1242  (.L_HI(net1242));
 sg13g2_tiehi \shift_storage.storage[1580]$_SDFFE_PN0P__1243  (.L_HI(net1243));
 sg13g2_tiehi \shift_storage.storage[1581]$_SDFFE_PN0P__1244  (.L_HI(net1244));
 sg13g2_tiehi \shift_storage.storage[1582]$_SDFFE_PN0P__1245  (.L_HI(net1245));
 sg13g2_tiehi \shift_storage.storage[1583]$_SDFFE_PN0P__1246  (.L_HI(net1246));
 sg13g2_tiehi \shift_storage.storage[1584]$_SDFFE_PN0P__1247  (.L_HI(net1247));
 sg13g2_tiehi \shift_storage.storage[1585]$_SDFFE_PN0P__1248  (.L_HI(net1248));
 sg13g2_tiehi \shift_storage.storage[1586]$_SDFFE_PN0P__1249  (.L_HI(net1249));
 sg13g2_tiehi \shift_storage.storage[1587]$_SDFFE_PN0P__1250  (.L_HI(net1250));
 sg13g2_tiehi \shift_storage.storage[1588]$_SDFFE_PN0P__1251  (.L_HI(net1251));
 sg13g2_tiehi \shift_storage.storage[1589]$_SDFFE_PN0P__1252  (.L_HI(net1252));
 sg13g2_tiehi \shift_storage.storage[158]$_SDFFE_PN0P__1253  (.L_HI(net1253));
 sg13g2_tiehi \shift_storage.storage[1590]$_SDFFE_PN0P__1254  (.L_HI(net1254));
 sg13g2_tiehi \shift_storage.storage[1591]$_SDFFE_PN0P__1255  (.L_HI(net1255));
 sg13g2_tiehi \shift_storage.storage[1592]$_SDFFE_PN0P__1256  (.L_HI(net1256));
 sg13g2_tiehi \shift_storage.storage[1593]$_SDFFE_PN0P__1257  (.L_HI(net1257));
 sg13g2_tiehi \shift_storage.storage[1594]$_SDFFE_PN0P__1258  (.L_HI(net1258));
 sg13g2_tiehi \shift_storage.storage[1595]$_SDFFE_PN0P__1259  (.L_HI(net1259));
 sg13g2_tiehi \shift_storage.storage[1596]$_SDFFE_PN0P__1260  (.L_HI(net1260));
 sg13g2_tiehi \shift_storage.storage[1597]$_SDFFE_PN0P__1261  (.L_HI(net1261));
 sg13g2_tiehi \shift_storage.storage[1598]$_SDFFE_PN0P__1262  (.L_HI(net1262));
 sg13g2_tiehi \shift_storage.storage[1599]$_SDFFE_PN0P__1263  (.L_HI(net1263));
 sg13g2_tiehi \shift_storage.storage[159]$_SDFFE_PN0P__1264  (.L_HI(net1264));
 sg13g2_tiehi \shift_storage.storage[15]$_SDFFE_PN0P__1265  (.L_HI(net1265));
 sg13g2_tiehi \shift_storage.storage[160]$_SDFFE_PN0P__1266  (.L_HI(net1266));
 sg13g2_tiehi \shift_storage.storage[161]$_SDFFE_PN0P__1267  (.L_HI(net1267));
 sg13g2_tiehi \shift_storage.storage[162]$_SDFFE_PN0P__1268  (.L_HI(net1268));
 sg13g2_tiehi \shift_storage.storage[163]$_SDFFE_PN0P__1269  (.L_HI(net1269));
 sg13g2_tiehi \shift_storage.storage[164]$_SDFFE_PN0P__1270  (.L_HI(net1270));
 sg13g2_tiehi \shift_storage.storage[165]$_SDFFE_PN0P__1271  (.L_HI(net1271));
 sg13g2_tiehi \shift_storage.storage[166]$_SDFFE_PN0P__1272  (.L_HI(net1272));
 sg13g2_tiehi \shift_storage.storage[167]$_SDFFE_PN0P__1273  (.L_HI(net1273));
 sg13g2_tiehi \shift_storage.storage[168]$_SDFFE_PN0P__1274  (.L_HI(net1274));
 sg13g2_tiehi \shift_storage.storage[169]$_SDFFE_PN0P__1275  (.L_HI(net1275));
 sg13g2_tiehi \shift_storage.storage[16]$_SDFFE_PN0P__1276  (.L_HI(net1276));
 sg13g2_tiehi \shift_storage.storage[170]$_SDFFE_PN0P__1277  (.L_HI(net1277));
 sg13g2_tiehi \shift_storage.storage[171]$_SDFFE_PN0P__1278  (.L_HI(net1278));
 sg13g2_tiehi \shift_storage.storage[172]$_SDFFE_PN0P__1279  (.L_HI(net1279));
 sg13g2_tiehi \shift_storage.storage[173]$_SDFFE_PN0P__1280  (.L_HI(net1280));
 sg13g2_tiehi \shift_storage.storage[174]$_SDFFE_PN0P__1281  (.L_HI(net1281));
 sg13g2_tiehi \shift_storage.storage[175]$_SDFFE_PN0P__1282  (.L_HI(net1282));
 sg13g2_tiehi \shift_storage.storage[176]$_SDFFE_PN0P__1283  (.L_HI(net1283));
 sg13g2_tiehi \shift_storage.storage[177]$_SDFFE_PN0P__1284  (.L_HI(net1284));
 sg13g2_tiehi \shift_storage.storage[178]$_SDFFE_PN0P__1285  (.L_HI(net1285));
 sg13g2_tiehi \shift_storage.storage[179]$_SDFFE_PN0P__1286  (.L_HI(net1286));
 sg13g2_tiehi \shift_storage.storage[17]$_SDFFE_PN0P__1287  (.L_HI(net1287));
 sg13g2_tiehi \shift_storage.storage[180]$_SDFFE_PN0P__1288  (.L_HI(net1288));
 sg13g2_tiehi \shift_storage.storage[181]$_SDFFE_PN0P__1289  (.L_HI(net1289));
 sg13g2_tiehi \shift_storage.storage[182]$_SDFFE_PN0P__1290  (.L_HI(net1290));
 sg13g2_tiehi \shift_storage.storage[183]$_SDFFE_PN0P__1291  (.L_HI(net1291));
 sg13g2_tiehi \shift_storage.storage[184]$_SDFFE_PN0P__1292  (.L_HI(net1292));
 sg13g2_tiehi \shift_storage.storage[185]$_SDFFE_PN0P__1293  (.L_HI(net1293));
 sg13g2_tiehi \shift_storage.storage[186]$_SDFFE_PN0P__1294  (.L_HI(net1294));
 sg13g2_tiehi \shift_storage.storage[187]$_SDFFE_PN0P__1295  (.L_HI(net1295));
 sg13g2_tiehi \shift_storage.storage[188]$_SDFFE_PN0P__1296  (.L_HI(net1296));
 sg13g2_tiehi \shift_storage.storage[189]$_SDFFE_PN0P__1297  (.L_HI(net1297));
 sg13g2_tiehi \shift_storage.storage[18]$_SDFFE_PN0P__1298  (.L_HI(net1298));
 sg13g2_tiehi \shift_storage.storage[190]$_SDFFE_PN0P__1299  (.L_HI(net1299));
 sg13g2_tiehi \shift_storage.storage[191]$_SDFFE_PN0P__1300  (.L_HI(net1300));
 sg13g2_tiehi \shift_storage.storage[192]$_SDFFE_PN0P__1301  (.L_HI(net1301));
 sg13g2_tiehi \shift_storage.storage[193]$_SDFFE_PN0P__1302  (.L_HI(net1302));
 sg13g2_tiehi \shift_storage.storage[194]$_SDFFE_PN0P__1303  (.L_HI(net1303));
 sg13g2_tiehi \shift_storage.storage[195]$_SDFFE_PN0P__1304  (.L_HI(net1304));
 sg13g2_tiehi \shift_storage.storage[196]$_SDFFE_PN0P__1305  (.L_HI(net1305));
 sg13g2_tiehi \shift_storage.storage[197]$_SDFFE_PN0P__1306  (.L_HI(net1306));
 sg13g2_tiehi \shift_storage.storage[198]$_SDFFE_PN0P__1307  (.L_HI(net1307));
 sg13g2_tiehi \shift_storage.storage[199]$_SDFFE_PN0P__1308  (.L_HI(net1308));
 sg13g2_tiehi \shift_storage.storage[19]$_SDFFE_PN0P__1309  (.L_HI(net1309));
 sg13g2_tiehi \shift_storage.storage[1]$_SDFFE_PN0P__1310  (.L_HI(net1310));
 sg13g2_tiehi \shift_storage.storage[200]$_SDFFE_PN0P__1311  (.L_HI(net1311));
 sg13g2_tiehi \shift_storage.storage[201]$_SDFFE_PN0P__1312  (.L_HI(net1312));
 sg13g2_tiehi \shift_storage.storage[202]$_SDFFE_PN0P__1313  (.L_HI(net1313));
 sg13g2_tiehi \shift_storage.storage[203]$_SDFFE_PN0P__1314  (.L_HI(net1314));
 sg13g2_tiehi \shift_storage.storage[204]$_SDFFE_PN0P__1315  (.L_HI(net1315));
 sg13g2_tiehi \shift_storage.storage[205]$_SDFFE_PN0P__1316  (.L_HI(net1316));
 sg13g2_tiehi \shift_storage.storage[206]$_SDFFE_PN0P__1317  (.L_HI(net1317));
 sg13g2_tiehi \shift_storage.storage[207]$_SDFFE_PN0P__1318  (.L_HI(net1318));
 sg13g2_tiehi \shift_storage.storage[208]$_SDFFE_PN0P__1319  (.L_HI(net1319));
 sg13g2_tiehi \shift_storage.storage[209]$_SDFFE_PN0P__1320  (.L_HI(net1320));
 sg13g2_tiehi \shift_storage.storage[20]$_SDFFE_PN0P__1321  (.L_HI(net1321));
 sg13g2_tiehi \shift_storage.storage[210]$_SDFFE_PN0P__1322  (.L_HI(net1322));
 sg13g2_tiehi \shift_storage.storage[211]$_SDFFE_PN0P__1323  (.L_HI(net1323));
 sg13g2_tiehi \shift_storage.storage[212]$_SDFFE_PN0P__1324  (.L_HI(net1324));
 sg13g2_tiehi \shift_storage.storage[213]$_SDFFE_PN0P__1325  (.L_HI(net1325));
 sg13g2_tiehi \shift_storage.storage[214]$_SDFFE_PN0P__1326  (.L_HI(net1326));
 sg13g2_tiehi \shift_storage.storage[215]$_SDFFE_PN0P__1327  (.L_HI(net1327));
 sg13g2_tiehi \shift_storage.storage[216]$_SDFFE_PN0P__1328  (.L_HI(net1328));
 sg13g2_tiehi \shift_storage.storage[217]$_SDFFE_PN0P__1329  (.L_HI(net1329));
 sg13g2_tiehi \shift_storage.storage[218]$_SDFFE_PN0P__1330  (.L_HI(net1330));
 sg13g2_tiehi \shift_storage.storage[219]$_SDFFE_PN0P__1331  (.L_HI(net1331));
 sg13g2_tiehi \shift_storage.storage[21]$_SDFFE_PN0P__1332  (.L_HI(net1332));
 sg13g2_tiehi \shift_storage.storage[220]$_SDFFE_PN0P__1333  (.L_HI(net1333));
 sg13g2_tiehi \shift_storage.storage[221]$_SDFFE_PN0P__1334  (.L_HI(net1334));
 sg13g2_tiehi \shift_storage.storage[222]$_SDFFE_PN0P__1335  (.L_HI(net1335));
 sg13g2_tiehi \shift_storage.storage[223]$_SDFFE_PN0P__1336  (.L_HI(net1336));
 sg13g2_tiehi \shift_storage.storage[224]$_SDFFE_PN0P__1337  (.L_HI(net1337));
 sg13g2_tiehi \shift_storage.storage[225]$_SDFFE_PN0P__1338  (.L_HI(net1338));
 sg13g2_tiehi \shift_storage.storage[226]$_SDFFE_PN0P__1339  (.L_HI(net1339));
 sg13g2_tiehi \shift_storage.storage[227]$_SDFFE_PN0P__1340  (.L_HI(net1340));
 sg13g2_tiehi \shift_storage.storage[228]$_SDFFE_PN0P__1341  (.L_HI(net1341));
 sg13g2_tiehi \shift_storage.storage[229]$_SDFFE_PN0P__1342  (.L_HI(net1342));
 sg13g2_tiehi \shift_storage.storage[22]$_SDFFE_PN0P__1343  (.L_HI(net1343));
 sg13g2_tiehi \shift_storage.storage[230]$_SDFFE_PN0P__1344  (.L_HI(net1344));
 sg13g2_tiehi \shift_storage.storage[231]$_SDFFE_PN0P__1345  (.L_HI(net1345));
 sg13g2_tiehi \shift_storage.storage[232]$_SDFFE_PN0P__1346  (.L_HI(net1346));
 sg13g2_tiehi \shift_storage.storage[233]$_SDFFE_PN0P__1347  (.L_HI(net1347));
 sg13g2_tiehi \shift_storage.storage[234]$_SDFFE_PN0P__1348  (.L_HI(net1348));
 sg13g2_tiehi \shift_storage.storage[235]$_SDFFE_PN0P__1349  (.L_HI(net1349));
 sg13g2_tiehi \shift_storage.storage[236]$_SDFFE_PN0P__1350  (.L_HI(net1350));
 sg13g2_tiehi \shift_storage.storage[237]$_SDFFE_PN0P__1351  (.L_HI(net1351));
 sg13g2_tiehi \shift_storage.storage[238]$_SDFFE_PN0P__1352  (.L_HI(net1352));
 sg13g2_tiehi \shift_storage.storage[239]$_SDFFE_PN0P__1353  (.L_HI(net1353));
 sg13g2_tiehi \shift_storage.storage[23]$_SDFFE_PN0P__1354  (.L_HI(net1354));
 sg13g2_tiehi \shift_storage.storage[240]$_SDFFE_PN0P__1355  (.L_HI(net1355));
 sg13g2_tiehi \shift_storage.storage[241]$_SDFFE_PN0P__1356  (.L_HI(net1356));
 sg13g2_tiehi \shift_storage.storage[242]$_SDFFE_PN0P__1357  (.L_HI(net1357));
 sg13g2_tiehi \shift_storage.storage[243]$_SDFFE_PN0P__1358  (.L_HI(net1358));
 sg13g2_tiehi \shift_storage.storage[244]$_SDFFE_PN0P__1359  (.L_HI(net1359));
 sg13g2_tiehi \shift_storage.storage[245]$_SDFFE_PN0P__1360  (.L_HI(net1360));
 sg13g2_tiehi \shift_storage.storage[246]$_SDFFE_PN0P__1361  (.L_HI(net1361));
 sg13g2_tiehi \shift_storage.storage[247]$_SDFFE_PN0P__1362  (.L_HI(net1362));
 sg13g2_tiehi \shift_storage.storage[248]$_SDFFE_PN0P__1363  (.L_HI(net1363));
 sg13g2_tiehi \shift_storage.storage[249]$_SDFFE_PN0P__1364  (.L_HI(net1364));
 sg13g2_tiehi \shift_storage.storage[24]$_SDFFE_PN0P__1365  (.L_HI(net1365));
 sg13g2_tiehi \shift_storage.storage[250]$_SDFFE_PN0P__1366  (.L_HI(net1366));
 sg13g2_tiehi \shift_storage.storage[251]$_SDFFE_PN0P__1367  (.L_HI(net1367));
 sg13g2_tiehi \shift_storage.storage[252]$_SDFFE_PN0P__1368  (.L_HI(net1368));
 sg13g2_tiehi \shift_storage.storage[253]$_SDFFE_PN0P__1369  (.L_HI(net1369));
 sg13g2_tiehi \shift_storage.storage[254]$_SDFFE_PN0P__1370  (.L_HI(net1370));
 sg13g2_tiehi \shift_storage.storage[255]$_SDFFE_PN0P__1371  (.L_HI(net1371));
 sg13g2_tiehi \shift_storage.storage[256]$_SDFFE_PN0P__1372  (.L_HI(net1372));
 sg13g2_tiehi \shift_storage.storage[257]$_SDFFE_PN0P__1373  (.L_HI(net1373));
 sg13g2_tiehi \shift_storage.storage[258]$_SDFFE_PN0P__1374  (.L_HI(net1374));
 sg13g2_tiehi \shift_storage.storage[259]$_SDFFE_PN0P__1375  (.L_HI(net1375));
 sg13g2_tiehi \shift_storage.storage[25]$_SDFFE_PN0P__1376  (.L_HI(net1376));
 sg13g2_tiehi \shift_storage.storage[260]$_SDFFE_PN0P__1377  (.L_HI(net1377));
 sg13g2_tiehi \shift_storage.storage[261]$_SDFFE_PN0P__1378  (.L_HI(net1378));
 sg13g2_tiehi \shift_storage.storage[262]$_SDFFE_PN0P__1379  (.L_HI(net1379));
 sg13g2_tiehi \shift_storage.storage[263]$_SDFFE_PN0P__1380  (.L_HI(net1380));
 sg13g2_tiehi \shift_storage.storage[264]$_SDFFE_PN0P__1381  (.L_HI(net1381));
 sg13g2_tiehi \shift_storage.storage[265]$_SDFFE_PN0P__1382  (.L_HI(net1382));
 sg13g2_tiehi \shift_storage.storage[266]$_SDFFE_PN0P__1383  (.L_HI(net1383));
 sg13g2_tiehi \shift_storage.storage[267]$_SDFFE_PN0P__1384  (.L_HI(net1384));
 sg13g2_tiehi \shift_storage.storage[268]$_SDFFE_PN0P__1385  (.L_HI(net1385));
 sg13g2_tiehi \shift_storage.storage[269]$_SDFFE_PN0P__1386  (.L_HI(net1386));
 sg13g2_tiehi \shift_storage.storage[26]$_SDFFE_PN0P__1387  (.L_HI(net1387));
 sg13g2_tiehi \shift_storage.storage[270]$_SDFFE_PN0P__1388  (.L_HI(net1388));
 sg13g2_tiehi \shift_storage.storage[271]$_SDFFE_PN0P__1389  (.L_HI(net1389));
 sg13g2_tiehi \shift_storage.storage[272]$_SDFFE_PN0P__1390  (.L_HI(net1390));
 sg13g2_tiehi \shift_storage.storage[273]$_SDFFE_PN0P__1391  (.L_HI(net1391));
 sg13g2_tiehi \shift_storage.storage[274]$_SDFFE_PN0P__1392  (.L_HI(net1392));
 sg13g2_tiehi \shift_storage.storage[275]$_SDFFE_PN0P__1393  (.L_HI(net1393));
 sg13g2_tiehi \shift_storage.storage[276]$_SDFFE_PN0P__1394  (.L_HI(net1394));
 sg13g2_tiehi \shift_storage.storage[277]$_SDFFE_PN0P__1395  (.L_HI(net1395));
 sg13g2_tiehi \shift_storage.storage[278]$_SDFFE_PN0P__1396  (.L_HI(net1396));
 sg13g2_tiehi \shift_storage.storage[279]$_SDFFE_PN0P__1397  (.L_HI(net1397));
 sg13g2_tiehi \shift_storage.storage[27]$_SDFFE_PN0P__1398  (.L_HI(net1398));
 sg13g2_tiehi \shift_storage.storage[280]$_SDFFE_PN0P__1399  (.L_HI(net1399));
 sg13g2_tiehi \shift_storage.storage[281]$_SDFFE_PN0P__1400  (.L_HI(net1400));
 sg13g2_tiehi \shift_storage.storage[282]$_SDFFE_PN0P__1401  (.L_HI(net1401));
 sg13g2_tiehi \shift_storage.storage[283]$_SDFFE_PN0P__1402  (.L_HI(net1402));
 sg13g2_tiehi \shift_storage.storage[284]$_SDFFE_PN0P__1403  (.L_HI(net1403));
 sg13g2_tiehi \shift_storage.storage[285]$_SDFFE_PN0P__1404  (.L_HI(net1404));
 sg13g2_tiehi \shift_storage.storage[286]$_SDFFE_PN0P__1405  (.L_HI(net1405));
 sg13g2_tiehi \shift_storage.storage[287]$_SDFFE_PN0P__1406  (.L_HI(net1406));
 sg13g2_tiehi \shift_storage.storage[288]$_SDFFE_PN0P__1407  (.L_HI(net1407));
 sg13g2_tiehi \shift_storage.storage[289]$_SDFFE_PN0P__1408  (.L_HI(net1408));
 sg13g2_tiehi \shift_storage.storage[28]$_SDFFE_PN0P__1409  (.L_HI(net1409));
 sg13g2_tiehi \shift_storage.storage[290]$_SDFFE_PN0P__1410  (.L_HI(net1410));
 sg13g2_tiehi \shift_storage.storage[291]$_SDFFE_PN0P__1411  (.L_HI(net1411));
 sg13g2_tiehi \shift_storage.storage[292]$_SDFFE_PN0P__1412  (.L_HI(net1412));
 sg13g2_tiehi \shift_storage.storage[293]$_SDFFE_PN0P__1413  (.L_HI(net1413));
 sg13g2_tiehi \shift_storage.storage[294]$_SDFFE_PN0P__1414  (.L_HI(net1414));
 sg13g2_tiehi \shift_storage.storage[295]$_SDFFE_PN0P__1415  (.L_HI(net1415));
 sg13g2_tiehi \shift_storage.storage[296]$_SDFFE_PN0P__1416  (.L_HI(net1416));
 sg13g2_tiehi \shift_storage.storage[297]$_SDFFE_PN0P__1417  (.L_HI(net1417));
 sg13g2_tiehi \shift_storage.storage[298]$_SDFFE_PN0P__1418  (.L_HI(net1418));
 sg13g2_tiehi \shift_storage.storage[299]$_SDFFE_PN0P__1419  (.L_HI(net1419));
 sg13g2_tiehi \shift_storage.storage[29]$_SDFFE_PN0P__1420  (.L_HI(net1420));
 sg13g2_tiehi \shift_storage.storage[2]$_SDFFE_PN0P__1421  (.L_HI(net1421));
 sg13g2_tiehi \shift_storage.storage[300]$_SDFFE_PN0P__1422  (.L_HI(net1422));
 sg13g2_tiehi \shift_storage.storage[301]$_SDFFE_PN0P__1423  (.L_HI(net1423));
 sg13g2_tiehi \shift_storage.storage[302]$_SDFFE_PN0P__1424  (.L_HI(net1424));
 sg13g2_tiehi \shift_storage.storage[303]$_SDFFE_PN0P__1425  (.L_HI(net1425));
 sg13g2_tiehi \shift_storage.storage[304]$_SDFFE_PN0P__1426  (.L_HI(net1426));
 sg13g2_tiehi \shift_storage.storage[305]$_SDFFE_PN0P__1427  (.L_HI(net1427));
 sg13g2_tiehi \shift_storage.storage[306]$_SDFFE_PN0P__1428  (.L_HI(net1428));
 sg13g2_tiehi \shift_storage.storage[307]$_SDFFE_PN0P__1429  (.L_HI(net1429));
 sg13g2_tiehi \shift_storage.storage[308]$_SDFFE_PN0P__1430  (.L_HI(net1430));
 sg13g2_tiehi \shift_storage.storage[309]$_SDFFE_PN0P__1431  (.L_HI(net1431));
 sg13g2_tiehi \shift_storage.storage[30]$_SDFFE_PN0P__1432  (.L_HI(net1432));
 sg13g2_tiehi \shift_storage.storage[310]$_SDFFE_PN0P__1433  (.L_HI(net1433));
 sg13g2_tiehi \shift_storage.storage[311]$_SDFFE_PN0P__1434  (.L_HI(net1434));
 sg13g2_tiehi \shift_storage.storage[312]$_SDFFE_PN0P__1435  (.L_HI(net1435));
 sg13g2_tiehi \shift_storage.storage[313]$_SDFFE_PN0P__1436  (.L_HI(net1436));
 sg13g2_tiehi \shift_storage.storage[314]$_SDFFE_PN0P__1437  (.L_HI(net1437));
 sg13g2_tiehi \shift_storage.storage[315]$_SDFFE_PN0P__1438  (.L_HI(net1438));
 sg13g2_tiehi \shift_storage.storage[316]$_SDFFE_PN0P__1439  (.L_HI(net1439));
 sg13g2_tiehi \shift_storage.storage[317]$_SDFFE_PN0P__1440  (.L_HI(net1440));
 sg13g2_tiehi \shift_storage.storage[318]$_SDFFE_PN0P__1441  (.L_HI(net1441));
 sg13g2_tiehi \shift_storage.storage[319]$_SDFFE_PN0P__1442  (.L_HI(net1442));
 sg13g2_tiehi \shift_storage.storage[31]$_SDFFE_PN0P__1443  (.L_HI(net1443));
 sg13g2_tiehi \shift_storage.storage[320]$_SDFFE_PN0P__1444  (.L_HI(net1444));
 sg13g2_tiehi \shift_storage.storage[321]$_SDFFE_PN0P__1445  (.L_HI(net1445));
 sg13g2_tiehi \shift_storage.storage[322]$_SDFFE_PN0P__1446  (.L_HI(net1446));
 sg13g2_tiehi \shift_storage.storage[323]$_SDFFE_PN0P__1447  (.L_HI(net1447));
 sg13g2_tiehi \shift_storage.storage[324]$_SDFFE_PN0P__1448  (.L_HI(net1448));
 sg13g2_tiehi \shift_storage.storage[325]$_SDFFE_PN0P__1449  (.L_HI(net1449));
 sg13g2_tiehi \shift_storage.storage[326]$_SDFFE_PN0P__1450  (.L_HI(net1450));
 sg13g2_tiehi \shift_storage.storage[327]$_SDFFE_PN0P__1451  (.L_HI(net1451));
 sg13g2_tiehi \shift_storage.storage[328]$_SDFFE_PN0P__1452  (.L_HI(net1452));
 sg13g2_tiehi \shift_storage.storage[329]$_SDFFE_PN0P__1453  (.L_HI(net1453));
 sg13g2_tiehi \shift_storage.storage[32]$_SDFFE_PN0P__1454  (.L_HI(net1454));
 sg13g2_tiehi \shift_storage.storage[330]$_SDFFE_PN0P__1455  (.L_HI(net1455));
 sg13g2_tiehi \shift_storage.storage[331]$_SDFFE_PN0P__1456  (.L_HI(net1456));
 sg13g2_tiehi \shift_storage.storage[332]$_SDFFE_PN0P__1457  (.L_HI(net1457));
 sg13g2_tiehi \shift_storage.storage[333]$_SDFFE_PN0P__1458  (.L_HI(net1458));
 sg13g2_tiehi \shift_storage.storage[334]$_SDFFE_PN0P__1459  (.L_HI(net1459));
 sg13g2_tiehi \shift_storage.storage[335]$_SDFFE_PN0P__1460  (.L_HI(net1460));
 sg13g2_tiehi \shift_storage.storage[336]$_SDFFE_PN0P__1461  (.L_HI(net1461));
 sg13g2_tiehi \shift_storage.storage[337]$_SDFFE_PN0P__1462  (.L_HI(net1462));
 sg13g2_tiehi \shift_storage.storage[338]$_SDFFE_PN0P__1463  (.L_HI(net1463));
 sg13g2_tiehi \shift_storage.storage[339]$_SDFFE_PN0P__1464  (.L_HI(net1464));
 sg13g2_tiehi \shift_storage.storage[33]$_SDFFE_PN0P__1465  (.L_HI(net1465));
 sg13g2_tiehi \shift_storage.storage[340]$_SDFFE_PN0P__1466  (.L_HI(net1466));
 sg13g2_tiehi \shift_storage.storage[341]$_SDFFE_PN0P__1467  (.L_HI(net1467));
 sg13g2_tiehi \shift_storage.storage[342]$_SDFFE_PN0P__1468  (.L_HI(net1468));
 sg13g2_tiehi \shift_storage.storage[343]$_SDFFE_PN0P__1469  (.L_HI(net1469));
 sg13g2_tiehi \shift_storage.storage[344]$_SDFFE_PN0P__1470  (.L_HI(net1470));
 sg13g2_tiehi \shift_storage.storage[345]$_SDFFE_PN0P__1471  (.L_HI(net1471));
 sg13g2_tiehi \shift_storage.storage[346]$_SDFFE_PN0P__1472  (.L_HI(net1472));
 sg13g2_tiehi \shift_storage.storage[347]$_SDFFE_PN0P__1473  (.L_HI(net1473));
 sg13g2_tiehi \shift_storage.storage[348]$_SDFFE_PN0P__1474  (.L_HI(net1474));
 sg13g2_tiehi \shift_storage.storage[349]$_SDFFE_PN0P__1475  (.L_HI(net1475));
 sg13g2_tiehi \shift_storage.storage[34]$_SDFFE_PN0P__1476  (.L_HI(net1476));
 sg13g2_tiehi \shift_storage.storage[350]$_SDFFE_PN0P__1477  (.L_HI(net1477));
 sg13g2_tiehi \shift_storage.storage[351]$_SDFFE_PN0P__1478  (.L_HI(net1478));
 sg13g2_tiehi \shift_storage.storage[352]$_SDFFE_PN0P__1479  (.L_HI(net1479));
 sg13g2_tiehi \shift_storage.storage[353]$_SDFFE_PN0P__1480  (.L_HI(net1480));
 sg13g2_tiehi \shift_storage.storage[354]$_SDFFE_PN0P__1481  (.L_HI(net1481));
 sg13g2_tiehi \shift_storage.storage[355]$_SDFFE_PN0P__1482  (.L_HI(net1482));
 sg13g2_tiehi \shift_storage.storage[356]$_SDFFE_PN0P__1483  (.L_HI(net1483));
 sg13g2_tiehi \shift_storage.storage[357]$_SDFFE_PN0P__1484  (.L_HI(net1484));
 sg13g2_tiehi \shift_storage.storage[358]$_SDFFE_PN0P__1485  (.L_HI(net1485));
 sg13g2_tiehi \shift_storage.storage[359]$_SDFFE_PN0P__1486  (.L_HI(net1486));
 sg13g2_tiehi \shift_storage.storage[35]$_SDFFE_PN0P__1487  (.L_HI(net1487));
 sg13g2_tiehi \shift_storage.storage[360]$_SDFFE_PN0P__1488  (.L_HI(net1488));
 sg13g2_tiehi \shift_storage.storage[361]$_SDFFE_PN0P__1489  (.L_HI(net1489));
 sg13g2_tiehi \shift_storage.storage[362]$_SDFFE_PN0P__1490  (.L_HI(net1490));
 sg13g2_tiehi \shift_storage.storage[363]$_SDFFE_PN0P__1491  (.L_HI(net1491));
 sg13g2_tiehi \shift_storage.storage[364]$_SDFFE_PN0P__1492  (.L_HI(net1492));
 sg13g2_tiehi \shift_storage.storage[365]$_SDFFE_PN0P__1493  (.L_HI(net1493));
 sg13g2_tiehi \shift_storage.storage[366]$_SDFFE_PN0P__1494  (.L_HI(net1494));
 sg13g2_tiehi \shift_storage.storage[367]$_SDFFE_PN0P__1495  (.L_HI(net1495));
 sg13g2_tiehi \shift_storage.storage[368]$_SDFFE_PN0P__1496  (.L_HI(net1496));
 sg13g2_tiehi \shift_storage.storage[369]$_SDFFE_PN0P__1497  (.L_HI(net1497));
 sg13g2_tiehi \shift_storage.storage[36]$_SDFFE_PN0P__1498  (.L_HI(net1498));
 sg13g2_tiehi \shift_storage.storage[370]$_SDFFE_PN0P__1499  (.L_HI(net1499));
 sg13g2_tiehi \shift_storage.storage[371]$_SDFFE_PN0P__1500  (.L_HI(net1500));
 sg13g2_tiehi \shift_storage.storage[372]$_SDFFE_PN0P__1501  (.L_HI(net1501));
 sg13g2_tiehi \shift_storage.storage[373]$_SDFFE_PN0P__1502  (.L_HI(net1502));
 sg13g2_tiehi \shift_storage.storage[374]$_SDFFE_PN0P__1503  (.L_HI(net1503));
 sg13g2_tiehi \shift_storage.storage[375]$_SDFFE_PN0P__1504  (.L_HI(net1504));
 sg13g2_tiehi \shift_storage.storage[376]$_SDFFE_PN0P__1505  (.L_HI(net1505));
 sg13g2_tiehi \shift_storage.storage[377]$_SDFFE_PN0P__1506  (.L_HI(net1506));
 sg13g2_tiehi \shift_storage.storage[378]$_SDFFE_PN0P__1507  (.L_HI(net1507));
 sg13g2_tiehi \shift_storage.storage[379]$_SDFFE_PN0P__1508  (.L_HI(net1508));
 sg13g2_tiehi \shift_storage.storage[37]$_SDFFE_PN0P__1509  (.L_HI(net1509));
 sg13g2_tiehi \shift_storage.storage[380]$_SDFFE_PN0P__1510  (.L_HI(net1510));
 sg13g2_tiehi \shift_storage.storage[381]$_SDFFE_PN0P__1511  (.L_HI(net1511));
 sg13g2_tiehi \shift_storage.storage[382]$_SDFFE_PN0P__1512  (.L_HI(net1512));
 sg13g2_tiehi \shift_storage.storage[383]$_SDFFE_PN0P__1513  (.L_HI(net1513));
 sg13g2_tiehi \shift_storage.storage[384]$_SDFFE_PN0P__1514  (.L_HI(net1514));
 sg13g2_tiehi \shift_storage.storage[385]$_SDFFE_PN0P__1515  (.L_HI(net1515));
 sg13g2_tiehi \shift_storage.storage[386]$_SDFFE_PN0P__1516  (.L_HI(net1516));
 sg13g2_tiehi \shift_storage.storage[387]$_SDFFE_PN0P__1517  (.L_HI(net1517));
 sg13g2_tiehi \shift_storage.storage[388]$_SDFFE_PN0P__1518  (.L_HI(net1518));
 sg13g2_tiehi \shift_storage.storage[389]$_SDFFE_PN0P__1519  (.L_HI(net1519));
 sg13g2_tiehi \shift_storage.storage[38]$_SDFFE_PN0P__1520  (.L_HI(net1520));
 sg13g2_tiehi \shift_storage.storage[390]$_SDFFE_PN0P__1521  (.L_HI(net1521));
 sg13g2_tiehi \shift_storage.storage[391]$_SDFFE_PN0P__1522  (.L_HI(net1522));
 sg13g2_tiehi \shift_storage.storage[392]$_SDFFE_PN0P__1523  (.L_HI(net1523));
 sg13g2_tiehi \shift_storage.storage[393]$_SDFFE_PN0P__1524  (.L_HI(net1524));
 sg13g2_tiehi \shift_storage.storage[394]$_SDFFE_PN0P__1525  (.L_HI(net1525));
 sg13g2_tiehi \shift_storage.storage[395]$_SDFFE_PN0P__1526  (.L_HI(net1526));
 sg13g2_tiehi \shift_storage.storage[396]$_SDFFE_PN0P__1527  (.L_HI(net1527));
 sg13g2_tiehi \shift_storage.storage[397]$_SDFFE_PN0P__1528  (.L_HI(net1528));
 sg13g2_tiehi \shift_storage.storage[398]$_SDFFE_PN0P__1529  (.L_HI(net1529));
 sg13g2_tiehi \shift_storage.storage[399]$_SDFFE_PN0P__1530  (.L_HI(net1530));
 sg13g2_tiehi \shift_storage.storage[39]$_SDFFE_PN0P__1531  (.L_HI(net1531));
 sg13g2_tiehi \shift_storage.storage[3]$_SDFFE_PN0P__1532  (.L_HI(net1532));
 sg13g2_tiehi \shift_storage.storage[400]$_SDFFE_PN0P__1533  (.L_HI(net1533));
 sg13g2_tiehi \shift_storage.storage[401]$_SDFFE_PN0P__1534  (.L_HI(net1534));
 sg13g2_tiehi \shift_storage.storage[402]$_SDFFE_PN0P__1535  (.L_HI(net1535));
 sg13g2_tiehi \shift_storage.storage[403]$_SDFFE_PN0P__1536  (.L_HI(net1536));
 sg13g2_tiehi \shift_storage.storage[404]$_SDFFE_PN0P__1537  (.L_HI(net1537));
 sg13g2_tiehi \shift_storage.storage[405]$_SDFFE_PN0P__1538  (.L_HI(net1538));
 sg13g2_tiehi \shift_storage.storage[406]$_SDFFE_PN0P__1539  (.L_HI(net1539));
 sg13g2_tiehi \shift_storage.storage[407]$_SDFFE_PN0P__1540  (.L_HI(net1540));
 sg13g2_tiehi \shift_storage.storage[408]$_SDFFE_PN0P__1541  (.L_HI(net1541));
 sg13g2_tiehi \shift_storage.storage[409]$_SDFFE_PN0P__1542  (.L_HI(net1542));
 sg13g2_tiehi \shift_storage.storage[40]$_SDFFE_PN0P__1543  (.L_HI(net1543));
 sg13g2_tiehi \shift_storage.storage[410]$_SDFFE_PN0P__1544  (.L_HI(net1544));
 sg13g2_tiehi \shift_storage.storage[411]$_SDFFE_PN0P__1545  (.L_HI(net1545));
 sg13g2_tiehi \shift_storage.storage[412]$_SDFFE_PN0P__1546  (.L_HI(net1546));
 sg13g2_tiehi \shift_storage.storage[413]$_SDFFE_PN0P__1547  (.L_HI(net1547));
 sg13g2_tiehi \shift_storage.storage[414]$_SDFFE_PN0P__1548  (.L_HI(net1548));
 sg13g2_tiehi \shift_storage.storage[415]$_SDFFE_PN0P__1549  (.L_HI(net1549));
 sg13g2_tiehi \shift_storage.storage[416]$_SDFFE_PN0P__1550  (.L_HI(net1550));
 sg13g2_tiehi \shift_storage.storage[417]$_SDFFE_PN0P__1551  (.L_HI(net1551));
 sg13g2_tiehi \shift_storage.storage[418]$_SDFFE_PN0P__1552  (.L_HI(net1552));
 sg13g2_tiehi \shift_storage.storage[419]$_SDFFE_PN0P__1553  (.L_HI(net1553));
 sg13g2_tiehi \shift_storage.storage[41]$_SDFFE_PN0P__1554  (.L_HI(net1554));
 sg13g2_tiehi \shift_storage.storage[420]$_SDFFE_PN0P__1555  (.L_HI(net1555));
 sg13g2_tiehi \shift_storage.storage[421]$_SDFFE_PN0P__1556  (.L_HI(net1556));
 sg13g2_tiehi \shift_storage.storage[422]$_SDFFE_PN0P__1557  (.L_HI(net1557));
 sg13g2_tiehi \shift_storage.storage[423]$_SDFFE_PN0P__1558  (.L_HI(net1558));
 sg13g2_tiehi \shift_storage.storage[424]$_SDFFE_PN0P__1559  (.L_HI(net1559));
 sg13g2_tiehi \shift_storage.storage[425]$_SDFFE_PN0P__1560  (.L_HI(net1560));
 sg13g2_tiehi \shift_storage.storage[426]$_SDFFE_PN0P__1561  (.L_HI(net1561));
 sg13g2_tiehi \shift_storage.storage[427]$_SDFFE_PN0P__1562  (.L_HI(net1562));
 sg13g2_tiehi \shift_storage.storage[428]$_SDFFE_PN0P__1563  (.L_HI(net1563));
 sg13g2_tiehi \shift_storage.storage[429]$_SDFFE_PN0P__1564  (.L_HI(net1564));
 sg13g2_tiehi \shift_storage.storage[42]$_SDFFE_PN0P__1565  (.L_HI(net1565));
 sg13g2_tiehi \shift_storage.storage[430]$_SDFFE_PN0P__1566  (.L_HI(net1566));
 sg13g2_tiehi \shift_storage.storage[431]$_SDFFE_PN0P__1567  (.L_HI(net1567));
 sg13g2_tiehi \shift_storage.storage[432]$_SDFFE_PN0P__1568  (.L_HI(net1568));
 sg13g2_tiehi \shift_storage.storage[433]$_SDFFE_PN0P__1569  (.L_HI(net1569));
 sg13g2_tiehi \shift_storage.storage[434]$_SDFFE_PN0P__1570  (.L_HI(net1570));
 sg13g2_tiehi \shift_storage.storage[435]$_SDFFE_PN0P__1571  (.L_HI(net1571));
 sg13g2_tiehi \shift_storage.storage[436]$_SDFFE_PN0P__1572  (.L_HI(net1572));
 sg13g2_tiehi \shift_storage.storage[437]$_SDFFE_PN0P__1573  (.L_HI(net1573));
 sg13g2_tiehi \shift_storage.storage[438]$_SDFFE_PN0P__1574  (.L_HI(net1574));
 sg13g2_tiehi \shift_storage.storage[439]$_SDFFE_PN0P__1575  (.L_HI(net1575));
 sg13g2_tiehi \shift_storage.storage[43]$_SDFFE_PN0P__1576  (.L_HI(net1576));
 sg13g2_tiehi \shift_storage.storage[440]$_SDFFE_PN0P__1577  (.L_HI(net1577));
 sg13g2_tiehi \shift_storage.storage[441]$_SDFFE_PN0P__1578  (.L_HI(net1578));
 sg13g2_tiehi \shift_storage.storage[442]$_SDFFE_PN0P__1579  (.L_HI(net1579));
 sg13g2_tiehi \shift_storage.storage[443]$_SDFFE_PN0P__1580  (.L_HI(net1580));
 sg13g2_tiehi \shift_storage.storage[444]$_SDFFE_PN0P__1581  (.L_HI(net1581));
 sg13g2_tiehi \shift_storage.storage[445]$_SDFFE_PN0P__1582  (.L_HI(net1582));
 sg13g2_tiehi \shift_storage.storage[446]$_SDFFE_PN0P__1583  (.L_HI(net1583));
 sg13g2_tiehi \shift_storage.storage[447]$_SDFFE_PN0P__1584  (.L_HI(net1584));
 sg13g2_tiehi \shift_storage.storage[448]$_SDFFE_PN0P__1585  (.L_HI(net1585));
 sg13g2_tiehi \shift_storage.storage[449]$_SDFFE_PN0P__1586  (.L_HI(net1586));
 sg13g2_tiehi \shift_storage.storage[44]$_SDFFE_PN0P__1587  (.L_HI(net1587));
 sg13g2_tiehi \shift_storage.storage[450]$_SDFFE_PN0P__1588  (.L_HI(net1588));
 sg13g2_tiehi \shift_storage.storage[451]$_SDFFE_PN0P__1589  (.L_HI(net1589));
 sg13g2_tiehi \shift_storage.storage[452]$_SDFFE_PN0P__1590  (.L_HI(net1590));
 sg13g2_tiehi \shift_storage.storage[453]$_SDFFE_PN0P__1591  (.L_HI(net1591));
 sg13g2_tiehi \shift_storage.storage[454]$_SDFFE_PN0P__1592  (.L_HI(net1592));
 sg13g2_tiehi \shift_storage.storage[455]$_SDFFE_PN0P__1593  (.L_HI(net1593));
 sg13g2_tiehi \shift_storage.storage[456]$_SDFFE_PN0P__1594  (.L_HI(net1594));
 sg13g2_tiehi \shift_storage.storage[457]$_SDFFE_PN0P__1595  (.L_HI(net1595));
 sg13g2_tiehi \shift_storage.storage[458]$_SDFFE_PN0P__1596  (.L_HI(net1596));
 sg13g2_tiehi \shift_storage.storage[459]$_SDFFE_PN0P__1597  (.L_HI(net1597));
 sg13g2_tiehi \shift_storage.storage[45]$_SDFFE_PN0P__1598  (.L_HI(net1598));
 sg13g2_tiehi \shift_storage.storage[460]$_SDFFE_PN0P__1599  (.L_HI(net1599));
 sg13g2_tiehi \shift_storage.storage[461]$_SDFFE_PN0P__1600  (.L_HI(net1600));
 sg13g2_tiehi \shift_storage.storage[462]$_SDFFE_PN0P__1601  (.L_HI(net1601));
 sg13g2_tiehi \shift_storage.storage[463]$_SDFFE_PN0P__1602  (.L_HI(net1602));
 sg13g2_tiehi \shift_storage.storage[464]$_SDFFE_PN0P__1603  (.L_HI(net1603));
 sg13g2_tiehi \shift_storage.storage[465]$_SDFFE_PN0P__1604  (.L_HI(net1604));
 sg13g2_tiehi \shift_storage.storage[466]$_SDFFE_PN0P__1605  (.L_HI(net1605));
 sg13g2_tiehi \shift_storage.storage[467]$_SDFFE_PN0P__1606  (.L_HI(net1606));
 sg13g2_tiehi \shift_storage.storage[468]$_SDFFE_PN0P__1607  (.L_HI(net1607));
 sg13g2_tiehi \shift_storage.storage[469]$_SDFFE_PN0P__1608  (.L_HI(net1608));
 sg13g2_tiehi \shift_storage.storage[46]$_SDFFE_PN0P__1609  (.L_HI(net1609));
 sg13g2_tiehi \shift_storage.storage[470]$_SDFFE_PN0P__1610  (.L_HI(net1610));
 sg13g2_tiehi \shift_storage.storage[471]$_SDFFE_PN0P__1611  (.L_HI(net1611));
 sg13g2_tiehi \shift_storage.storage[472]$_SDFFE_PN0P__1612  (.L_HI(net1612));
 sg13g2_tiehi \shift_storage.storage[473]$_SDFFE_PN0P__1613  (.L_HI(net1613));
 sg13g2_tiehi \shift_storage.storage[474]$_SDFFE_PN0P__1614  (.L_HI(net1614));
 sg13g2_tiehi \shift_storage.storage[475]$_SDFFE_PN0P__1615  (.L_HI(net1615));
 sg13g2_tiehi \shift_storage.storage[476]$_SDFFE_PN0P__1616  (.L_HI(net1616));
 sg13g2_tiehi \shift_storage.storage[477]$_SDFFE_PN0P__1617  (.L_HI(net1617));
 sg13g2_tiehi \shift_storage.storage[478]$_SDFFE_PN0P__1618  (.L_HI(net1618));
 sg13g2_tiehi \shift_storage.storage[479]$_SDFFE_PN0P__1619  (.L_HI(net1619));
 sg13g2_tiehi \shift_storage.storage[47]$_SDFFE_PN0P__1620  (.L_HI(net1620));
 sg13g2_tiehi \shift_storage.storage[480]$_SDFFE_PN0P__1621  (.L_HI(net1621));
 sg13g2_tiehi \shift_storage.storage[481]$_SDFFE_PN0P__1622  (.L_HI(net1622));
 sg13g2_tiehi \shift_storage.storage[482]$_SDFFE_PN0P__1623  (.L_HI(net1623));
 sg13g2_tiehi \shift_storage.storage[483]$_SDFFE_PN0P__1624  (.L_HI(net1624));
 sg13g2_tiehi \shift_storage.storage[484]$_SDFFE_PN0P__1625  (.L_HI(net1625));
 sg13g2_tiehi \shift_storage.storage[485]$_SDFFE_PN0P__1626  (.L_HI(net1626));
 sg13g2_tiehi \shift_storage.storage[486]$_SDFFE_PN0P__1627  (.L_HI(net1627));
 sg13g2_tiehi \shift_storage.storage[487]$_SDFFE_PN0P__1628  (.L_HI(net1628));
 sg13g2_tiehi \shift_storage.storage[488]$_SDFFE_PN0P__1629  (.L_HI(net1629));
 sg13g2_tiehi \shift_storage.storage[489]$_SDFFE_PN0P__1630  (.L_HI(net1630));
 sg13g2_tiehi \shift_storage.storage[48]$_SDFFE_PN0P__1631  (.L_HI(net1631));
 sg13g2_tiehi \shift_storage.storage[490]$_SDFFE_PN0P__1632  (.L_HI(net1632));
 sg13g2_tiehi \shift_storage.storage[491]$_SDFFE_PN0P__1633  (.L_HI(net1633));
 sg13g2_tiehi \shift_storage.storage[492]$_SDFFE_PN0P__1634  (.L_HI(net1634));
 sg13g2_tiehi \shift_storage.storage[493]$_SDFFE_PN0P__1635  (.L_HI(net1635));
 sg13g2_tiehi \shift_storage.storage[494]$_SDFFE_PN0P__1636  (.L_HI(net1636));
 sg13g2_tiehi \shift_storage.storage[495]$_SDFFE_PN0P__1637  (.L_HI(net1637));
 sg13g2_tiehi \shift_storage.storage[496]$_SDFFE_PN0P__1638  (.L_HI(net1638));
 sg13g2_tiehi \shift_storage.storage[497]$_SDFFE_PN0P__1639  (.L_HI(net1639));
 sg13g2_tiehi \shift_storage.storage[498]$_SDFFE_PN0P__1640  (.L_HI(net1640));
 sg13g2_tiehi \shift_storage.storage[499]$_SDFFE_PN0P__1641  (.L_HI(net1641));
 sg13g2_tiehi \shift_storage.storage[49]$_SDFFE_PN0P__1642  (.L_HI(net1642));
 sg13g2_tiehi \shift_storage.storage[4]$_SDFFE_PN0P__1643  (.L_HI(net1643));
 sg13g2_tiehi \shift_storage.storage[500]$_SDFFE_PN0P__1644  (.L_HI(net1644));
 sg13g2_tiehi \shift_storage.storage[501]$_SDFFE_PN0P__1645  (.L_HI(net1645));
 sg13g2_tiehi \shift_storage.storage[502]$_SDFFE_PN0P__1646  (.L_HI(net1646));
 sg13g2_tiehi \shift_storage.storage[503]$_SDFFE_PN0P__1647  (.L_HI(net1647));
 sg13g2_tiehi \shift_storage.storage[504]$_SDFFE_PN0P__1648  (.L_HI(net1648));
 sg13g2_tiehi \shift_storage.storage[505]$_SDFFE_PN0P__1649  (.L_HI(net1649));
 sg13g2_tiehi \shift_storage.storage[506]$_SDFFE_PN0P__1650  (.L_HI(net1650));
 sg13g2_tiehi \shift_storage.storage[507]$_SDFFE_PN0P__1651  (.L_HI(net1651));
 sg13g2_tiehi \shift_storage.storage[508]$_SDFFE_PN0P__1652  (.L_HI(net1652));
 sg13g2_tiehi \shift_storage.storage[509]$_SDFFE_PN0P__1653  (.L_HI(net1653));
 sg13g2_tiehi \shift_storage.storage[50]$_SDFFE_PN0P__1654  (.L_HI(net1654));
 sg13g2_tiehi \shift_storage.storage[510]$_SDFFE_PN0P__1655  (.L_HI(net1655));
 sg13g2_tiehi \shift_storage.storage[511]$_SDFFE_PN0P__1656  (.L_HI(net1656));
 sg13g2_tiehi \shift_storage.storage[512]$_SDFFE_PN0P__1657  (.L_HI(net1657));
 sg13g2_tiehi \shift_storage.storage[513]$_SDFFE_PN0P__1658  (.L_HI(net1658));
 sg13g2_tiehi \shift_storage.storage[514]$_SDFFE_PN0P__1659  (.L_HI(net1659));
 sg13g2_tiehi \shift_storage.storage[515]$_SDFFE_PN0P__1660  (.L_HI(net1660));
 sg13g2_tiehi \shift_storage.storage[516]$_SDFFE_PN0P__1661  (.L_HI(net1661));
 sg13g2_tiehi \shift_storage.storage[517]$_SDFFE_PN0P__1662  (.L_HI(net1662));
 sg13g2_tiehi \shift_storage.storage[518]$_SDFFE_PN0P__1663  (.L_HI(net1663));
 sg13g2_tiehi \shift_storage.storage[519]$_SDFFE_PN0P__1664  (.L_HI(net1664));
 sg13g2_tiehi \shift_storage.storage[51]$_SDFFE_PN0P__1665  (.L_HI(net1665));
 sg13g2_tiehi \shift_storage.storage[520]$_SDFFE_PN0P__1666  (.L_HI(net1666));
 sg13g2_tiehi \shift_storage.storage[521]$_SDFFE_PN0P__1667  (.L_HI(net1667));
 sg13g2_tiehi \shift_storage.storage[522]$_SDFFE_PN0P__1668  (.L_HI(net1668));
 sg13g2_tiehi \shift_storage.storage[523]$_SDFFE_PN0P__1669  (.L_HI(net1669));
 sg13g2_tiehi \shift_storage.storage[524]$_SDFFE_PN0P__1670  (.L_HI(net1670));
 sg13g2_tiehi \shift_storage.storage[525]$_SDFFE_PN0P__1671  (.L_HI(net1671));
 sg13g2_tiehi \shift_storage.storage[526]$_SDFFE_PN0P__1672  (.L_HI(net1672));
 sg13g2_tiehi \shift_storage.storage[527]$_SDFFE_PN0P__1673  (.L_HI(net1673));
 sg13g2_tiehi \shift_storage.storage[528]$_SDFFE_PN0P__1674  (.L_HI(net1674));
 sg13g2_tiehi \shift_storage.storage[529]$_SDFFE_PN0P__1675  (.L_HI(net1675));
 sg13g2_tiehi \shift_storage.storage[52]$_SDFFE_PN0P__1676  (.L_HI(net1676));
 sg13g2_tiehi \shift_storage.storage[530]$_SDFFE_PN0P__1677  (.L_HI(net1677));
 sg13g2_tiehi \shift_storage.storage[531]$_SDFFE_PN0P__1678  (.L_HI(net1678));
 sg13g2_tiehi \shift_storage.storage[532]$_SDFFE_PN0P__1679  (.L_HI(net1679));
 sg13g2_tiehi \shift_storage.storage[533]$_SDFFE_PN0P__1680  (.L_HI(net1680));
 sg13g2_tiehi \shift_storage.storage[534]$_SDFFE_PN0P__1681  (.L_HI(net1681));
 sg13g2_tiehi \shift_storage.storage[535]$_SDFFE_PN0P__1682  (.L_HI(net1682));
 sg13g2_tiehi \shift_storage.storage[536]$_SDFFE_PN0P__1683  (.L_HI(net1683));
 sg13g2_tiehi \shift_storage.storage[537]$_SDFFE_PN0P__1684  (.L_HI(net1684));
 sg13g2_tiehi \shift_storage.storage[538]$_SDFFE_PN0P__1685  (.L_HI(net1685));
 sg13g2_tiehi \shift_storage.storage[539]$_SDFFE_PN0P__1686  (.L_HI(net1686));
 sg13g2_tiehi \shift_storage.storage[53]$_SDFFE_PN0P__1687  (.L_HI(net1687));
 sg13g2_tiehi \shift_storage.storage[540]$_SDFFE_PN0P__1688  (.L_HI(net1688));
 sg13g2_tiehi \shift_storage.storage[541]$_SDFFE_PN0P__1689  (.L_HI(net1689));
 sg13g2_tiehi \shift_storage.storage[542]$_SDFFE_PN0P__1690  (.L_HI(net1690));
 sg13g2_tiehi \shift_storage.storage[543]$_SDFFE_PN0P__1691  (.L_HI(net1691));
 sg13g2_tiehi \shift_storage.storage[544]$_SDFFE_PN0P__1692  (.L_HI(net1692));
 sg13g2_tiehi \shift_storage.storage[545]$_SDFFE_PN0P__1693  (.L_HI(net1693));
 sg13g2_tiehi \shift_storage.storage[546]$_SDFFE_PN0P__1694  (.L_HI(net1694));
 sg13g2_tiehi \shift_storage.storage[547]$_SDFFE_PN0P__1695  (.L_HI(net1695));
 sg13g2_tiehi \shift_storage.storage[548]$_SDFFE_PN0P__1696  (.L_HI(net1696));
 sg13g2_tiehi \shift_storage.storage[549]$_SDFFE_PN0P__1697  (.L_HI(net1697));
 sg13g2_tiehi \shift_storage.storage[54]$_SDFFE_PN0P__1698  (.L_HI(net1698));
 sg13g2_tiehi \shift_storage.storage[550]$_SDFFE_PN0P__1699  (.L_HI(net1699));
 sg13g2_tiehi \shift_storage.storage[551]$_SDFFE_PN0P__1700  (.L_HI(net1700));
 sg13g2_tiehi \shift_storage.storage[552]$_SDFFE_PN0P__1701  (.L_HI(net1701));
 sg13g2_tiehi \shift_storage.storage[553]$_SDFFE_PN0P__1702  (.L_HI(net1702));
 sg13g2_tiehi \shift_storage.storage[554]$_SDFFE_PN0P__1703  (.L_HI(net1703));
 sg13g2_tiehi \shift_storage.storage[555]$_SDFFE_PN0P__1704  (.L_HI(net1704));
 sg13g2_tiehi \shift_storage.storage[556]$_SDFFE_PN0P__1705  (.L_HI(net1705));
 sg13g2_tiehi \shift_storage.storage[557]$_SDFFE_PN0P__1706  (.L_HI(net1706));
 sg13g2_tiehi \shift_storage.storage[558]$_SDFFE_PN0P__1707  (.L_HI(net1707));
 sg13g2_tiehi \shift_storage.storage[559]$_SDFFE_PN0P__1708  (.L_HI(net1708));
 sg13g2_tiehi \shift_storage.storage[55]$_SDFFE_PN0P__1709  (.L_HI(net1709));
 sg13g2_tiehi \shift_storage.storage[560]$_SDFFE_PN0P__1710  (.L_HI(net1710));
 sg13g2_tiehi \shift_storage.storage[561]$_SDFFE_PN0P__1711  (.L_HI(net1711));
 sg13g2_tiehi \shift_storage.storage[562]$_SDFFE_PN0P__1712  (.L_HI(net1712));
 sg13g2_tiehi \shift_storage.storage[563]$_SDFFE_PN0P__1713  (.L_HI(net1713));
 sg13g2_tiehi \shift_storage.storage[564]$_SDFFE_PN0P__1714  (.L_HI(net1714));
 sg13g2_tiehi \shift_storage.storage[565]$_SDFFE_PN0P__1715  (.L_HI(net1715));
 sg13g2_tiehi \shift_storage.storage[566]$_SDFFE_PN0P__1716  (.L_HI(net1716));
 sg13g2_tiehi \shift_storage.storage[567]$_SDFFE_PN0P__1717  (.L_HI(net1717));
 sg13g2_tiehi \shift_storage.storage[568]$_SDFFE_PN0P__1718  (.L_HI(net1718));
 sg13g2_tiehi \shift_storage.storage[569]$_SDFFE_PN0P__1719  (.L_HI(net1719));
 sg13g2_tiehi \shift_storage.storage[56]$_SDFFE_PN0P__1720  (.L_HI(net1720));
 sg13g2_tiehi \shift_storage.storage[570]$_SDFFE_PN0P__1721  (.L_HI(net1721));
 sg13g2_tiehi \shift_storage.storage[571]$_SDFFE_PN0P__1722  (.L_HI(net1722));
 sg13g2_tiehi \shift_storage.storage[572]$_SDFFE_PN0P__1723  (.L_HI(net1723));
 sg13g2_tiehi \shift_storage.storage[573]$_SDFFE_PN0P__1724  (.L_HI(net1724));
 sg13g2_tiehi \shift_storage.storage[574]$_SDFFE_PN0P__1725  (.L_HI(net1725));
 sg13g2_tiehi \shift_storage.storage[575]$_SDFFE_PN0P__1726  (.L_HI(net1726));
 sg13g2_tiehi \shift_storage.storage[576]$_SDFFE_PN0P__1727  (.L_HI(net1727));
 sg13g2_tiehi \shift_storage.storage[577]$_SDFFE_PN0P__1728  (.L_HI(net1728));
 sg13g2_tiehi \shift_storage.storage[578]$_SDFFE_PN0P__1729  (.L_HI(net1729));
 sg13g2_tiehi \shift_storage.storage[579]$_SDFFE_PN0P__1730  (.L_HI(net1730));
 sg13g2_tiehi \shift_storage.storage[57]$_SDFFE_PN0P__1731  (.L_HI(net1731));
 sg13g2_tiehi \shift_storage.storage[580]$_SDFFE_PN0P__1732  (.L_HI(net1732));
 sg13g2_tiehi \shift_storage.storage[581]$_SDFFE_PN0P__1733  (.L_HI(net1733));
 sg13g2_tiehi \shift_storage.storage[582]$_SDFFE_PN0P__1734  (.L_HI(net1734));
 sg13g2_tiehi \shift_storage.storage[583]$_SDFFE_PN0P__1735  (.L_HI(net1735));
 sg13g2_tiehi \shift_storage.storage[584]$_SDFFE_PN0P__1736  (.L_HI(net1736));
 sg13g2_tiehi \shift_storage.storage[585]$_SDFFE_PN0P__1737  (.L_HI(net1737));
 sg13g2_tiehi \shift_storage.storage[586]$_SDFFE_PN0P__1738  (.L_HI(net1738));
 sg13g2_tiehi \shift_storage.storage[587]$_SDFFE_PN0P__1739  (.L_HI(net1739));
 sg13g2_tiehi \shift_storage.storage[588]$_SDFFE_PN0P__1740  (.L_HI(net1740));
 sg13g2_tiehi \shift_storage.storage[589]$_SDFFE_PN0P__1741  (.L_HI(net1741));
 sg13g2_tiehi \shift_storage.storage[58]$_SDFFE_PN0P__1742  (.L_HI(net1742));
 sg13g2_tiehi \shift_storage.storage[590]$_SDFFE_PN0P__1743  (.L_HI(net1743));
 sg13g2_tiehi \shift_storage.storage[591]$_SDFFE_PN0P__1744  (.L_HI(net1744));
 sg13g2_tiehi \shift_storage.storage[592]$_SDFFE_PN0P__1745  (.L_HI(net1745));
 sg13g2_tiehi \shift_storage.storage[593]$_SDFFE_PN0P__1746  (.L_HI(net1746));
 sg13g2_tiehi \shift_storage.storage[594]$_SDFFE_PN0P__1747  (.L_HI(net1747));
 sg13g2_tiehi \shift_storage.storage[595]$_SDFFE_PN0P__1748  (.L_HI(net1748));
 sg13g2_tiehi \shift_storage.storage[596]$_SDFFE_PN0P__1749  (.L_HI(net1749));
 sg13g2_tiehi \shift_storage.storage[597]$_SDFFE_PN0P__1750  (.L_HI(net1750));
 sg13g2_tiehi \shift_storage.storage[598]$_SDFFE_PN0P__1751  (.L_HI(net1751));
 sg13g2_tiehi \shift_storage.storage[599]$_SDFFE_PN0P__1752  (.L_HI(net1752));
 sg13g2_tiehi \shift_storage.storage[59]$_SDFFE_PN0P__1753  (.L_HI(net1753));
 sg13g2_tiehi \shift_storage.storage[5]$_SDFFE_PN0P__1754  (.L_HI(net1754));
 sg13g2_tiehi \shift_storage.storage[600]$_SDFFE_PN0P__1755  (.L_HI(net1755));
 sg13g2_tiehi \shift_storage.storage[601]$_SDFFE_PN0P__1756  (.L_HI(net1756));
 sg13g2_tiehi \shift_storage.storage[602]$_SDFFE_PN0P__1757  (.L_HI(net1757));
 sg13g2_tiehi \shift_storage.storage[603]$_SDFFE_PN0P__1758  (.L_HI(net1758));
 sg13g2_tiehi \shift_storage.storage[604]$_SDFFE_PN0P__1759  (.L_HI(net1759));
 sg13g2_tiehi \shift_storage.storage[605]$_SDFFE_PN0P__1760  (.L_HI(net1760));
 sg13g2_tiehi \shift_storage.storage[606]$_SDFFE_PN0P__1761  (.L_HI(net1761));
 sg13g2_tiehi \shift_storage.storage[607]$_SDFFE_PN0P__1762  (.L_HI(net1762));
 sg13g2_tiehi \shift_storage.storage[608]$_SDFFE_PN0P__1763  (.L_HI(net1763));
 sg13g2_tiehi \shift_storage.storage[609]$_SDFFE_PN0P__1764  (.L_HI(net1764));
 sg13g2_tiehi \shift_storage.storage[60]$_SDFFE_PN0P__1765  (.L_HI(net1765));
 sg13g2_tiehi \shift_storage.storage[610]$_SDFFE_PN0P__1766  (.L_HI(net1766));
 sg13g2_tiehi \shift_storage.storage[611]$_SDFFE_PN0P__1767  (.L_HI(net1767));
 sg13g2_tiehi \shift_storage.storage[612]$_SDFFE_PN0P__1768  (.L_HI(net1768));
 sg13g2_tiehi \shift_storage.storage[613]$_SDFFE_PN0P__1769  (.L_HI(net1769));
 sg13g2_tiehi \shift_storage.storage[614]$_SDFFE_PN0P__1770  (.L_HI(net1770));
 sg13g2_tiehi \shift_storage.storage[615]$_SDFFE_PN0P__1771  (.L_HI(net1771));
 sg13g2_tiehi \shift_storage.storage[616]$_SDFFE_PN0P__1772  (.L_HI(net1772));
 sg13g2_tiehi \shift_storage.storage[617]$_SDFFE_PN0P__1773  (.L_HI(net1773));
 sg13g2_tiehi \shift_storage.storage[618]$_SDFFE_PN0P__1774  (.L_HI(net1774));
 sg13g2_tiehi \shift_storage.storage[619]$_SDFFE_PN0P__1775  (.L_HI(net1775));
 sg13g2_tiehi \shift_storage.storage[61]$_SDFFE_PN0P__1776  (.L_HI(net1776));
 sg13g2_tiehi \shift_storage.storage[620]$_SDFFE_PN0P__1777  (.L_HI(net1777));
 sg13g2_tiehi \shift_storage.storage[621]$_SDFFE_PN0P__1778  (.L_HI(net1778));
 sg13g2_tiehi \shift_storage.storage[622]$_SDFFE_PN0P__1779  (.L_HI(net1779));
 sg13g2_tiehi \shift_storage.storage[623]$_SDFFE_PN0P__1780  (.L_HI(net1780));
 sg13g2_tiehi \shift_storage.storage[624]$_SDFFE_PN0P__1781  (.L_HI(net1781));
 sg13g2_tiehi \shift_storage.storage[625]$_SDFFE_PN0P__1782  (.L_HI(net1782));
 sg13g2_tiehi \shift_storage.storage[626]$_SDFFE_PN0P__1783  (.L_HI(net1783));
 sg13g2_tiehi \shift_storage.storage[627]$_SDFFE_PN0P__1784  (.L_HI(net1784));
 sg13g2_tiehi \shift_storage.storage[628]$_SDFFE_PN0P__1785  (.L_HI(net1785));
 sg13g2_tiehi \shift_storage.storage[629]$_SDFFE_PN0P__1786  (.L_HI(net1786));
 sg13g2_tiehi \shift_storage.storage[62]$_SDFFE_PN0P__1787  (.L_HI(net1787));
 sg13g2_tiehi \shift_storage.storage[630]$_SDFFE_PN0P__1788  (.L_HI(net1788));
 sg13g2_tiehi \shift_storage.storage[631]$_SDFFE_PN0P__1789  (.L_HI(net1789));
 sg13g2_tiehi \shift_storage.storage[632]$_SDFFE_PN0P__1790  (.L_HI(net1790));
 sg13g2_tiehi \shift_storage.storage[633]$_SDFFE_PN0P__1791  (.L_HI(net1791));
 sg13g2_tiehi \shift_storage.storage[634]$_SDFFE_PN0P__1792  (.L_HI(net1792));
 sg13g2_tiehi \shift_storage.storage[635]$_SDFFE_PN0P__1793  (.L_HI(net1793));
 sg13g2_tiehi \shift_storage.storage[636]$_SDFFE_PN0P__1794  (.L_HI(net1794));
 sg13g2_tiehi \shift_storage.storage[637]$_SDFFE_PN0P__1795  (.L_HI(net1795));
 sg13g2_tiehi \shift_storage.storage[638]$_SDFFE_PN0P__1796  (.L_HI(net1796));
 sg13g2_tiehi \shift_storage.storage[639]$_SDFFE_PN0P__1797  (.L_HI(net1797));
 sg13g2_tiehi \shift_storage.storage[63]$_SDFFE_PN0P__1798  (.L_HI(net1798));
 sg13g2_tiehi \shift_storage.storage[640]$_SDFFE_PN0P__1799  (.L_HI(net1799));
 sg13g2_tiehi \shift_storage.storage[641]$_SDFFE_PN0P__1800  (.L_HI(net1800));
 sg13g2_tiehi \shift_storage.storage[642]$_SDFFE_PN0P__1801  (.L_HI(net1801));
 sg13g2_tiehi \shift_storage.storage[643]$_SDFFE_PN0P__1802  (.L_HI(net1802));
 sg13g2_tiehi \shift_storage.storage[644]$_SDFFE_PN0P__1803  (.L_HI(net1803));
 sg13g2_tiehi \shift_storage.storage[645]$_SDFFE_PN0P__1804  (.L_HI(net1804));
 sg13g2_tiehi \shift_storage.storage[646]$_SDFFE_PN0P__1805  (.L_HI(net1805));
 sg13g2_tiehi \shift_storage.storage[647]$_SDFFE_PN0P__1806  (.L_HI(net1806));
 sg13g2_tiehi \shift_storage.storage[648]$_SDFFE_PN0P__1807  (.L_HI(net1807));
 sg13g2_tiehi \shift_storage.storage[649]$_SDFFE_PN0P__1808  (.L_HI(net1808));
 sg13g2_tiehi \shift_storage.storage[64]$_SDFFE_PN0P__1809  (.L_HI(net1809));
 sg13g2_tiehi \shift_storage.storage[650]$_SDFFE_PN0P__1810  (.L_HI(net1810));
 sg13g2_tiehi \shift_storage.storage[651]$_SDFFE_PN0P__1811  (.L_HI(net1811));
 sg13g2_tiehi \shift_storage.storage[652]$_SDFFE_PN0P__1812  (.L_HI(net1812));
 sg13g2_tiehi \shift_storage.storage[653]$_SDFFE_PN0P__1813  (.L_HI(net1813));
 sg13g2_tiehi \shift_storage.storage[654]$_SDFFE_PN0P__1814  (.L_HI(net1814));
 sg13g2_tiehi \shift_storage.storage[655]$_SDFFE_PN0P__1815  (.L_HI(net1815));
 sg13g2_tiehi \shift_storage.storage[656]$_SDFFE_PN0P__1816  (.L_HI(net1816));
 sg13g2_tiehi \shift_storage.storage[657]$_SDFFE_PN0P__1817  (.L_HI(net1817));
 sg13g2_tiehi \shift_storage.storage[658]$_SDFFE_PN0P__1818  (.L_HI(net1818));
 sg13g2_tiehi \shift_storage.storage[659]$_SDFFE_PN0P__1819  (.L_HI(net1819));
 sg13g2_tiehi \shift_storage.storage[65]$_SDFFE_PN0P__1820  (.L_HI(net1820));
 sg13g2_tiehi \shift_storage.storage[660]$_SDFFE_PN0P__1821  (.L_HI(net1821));
 sg13g2_tiehi \shift_storage.storage[661]$_SDFFE_PN0P__1822  (.L_HI(net1822));
 sg13g2_tiehi \shift_storage.storage[662]$_SDFFE_PN0P__1823  (.L_HI(net1823));
 sg13g2_tiehi \shift_storage.storage[663]$_SDFFE_PN0P__1824  (.L_HI(net1824));
 sg13g2_tiehi \shift_storage.storage[664]$_SDFFE_PN0P__1825  (.L_HI(net1825));
 sg13g2_tiehi \shift_storage.storage[665]$_SDFFE_PN0P__1826  (.L_HI(net1826));
 sg13g2_tiehi \shift_storage.storage[666]$_SDFFE_PN0P__1827  (.L_HI(net1827));
 sg13g2_tiehi \shift_storage.storage[667]$_SDFFE_PN0P__1828  (.L_HI(net1828));
 sg13g2_tiehi \shift_storage.storage[668]$_SDFFE_PN0P__1829  (.L_HI(net1829));
 sg13g2_tiehi \shift_storage.storage[669]$_SDFFE_PN0P__1830  (.L_HI(net1830));
 sg13g2_tiehi \shift_storage.storage[66]$_SDFFE_PN0P__1831  (.L_HI(net1831));
 sg13g2_tiehi \shift_storage.storage[670]$_SDFFE_PN0P__1832  (.L_HI(net1832));
 sg13g2_tiehi \shift_storage.storage[671]$_SDFFE_PN0P__1833  (.L_HI(net1833));
 sg13g2_tiehi \shift_storage.storage[672]$_SDFFE_PN0P__1834  (.L_HI(net1834));
 sg13g2_tiehi \shift_storage.storage[673]$_SDFFE_PN0P__1835  (.L_HI(net1835));
 sg13g2_tiehi \shift_storage.storage[674]$_SDFFE_PN0P__1836  (.L_HI(net1836));
 sg13g2_tiehi \shift_storage.storage[675]$_SDFFE_PN0P__1837  (.L_HI(net1837));
 sg13g2_tiehi \shift_storage.storage[676]$_SDFFE_PN0P__1838  (.L_HI(net1838));
 sg13g2_tiehi \shift_storage.storage[677]$_SDFFE_PN0P__1839  (.L_HI(net1839));
 sg13g2_tiehi \shift_storage.storage[678]$_SDFFE_PN0P__1840  (.L_HI(net1840));
 sg13g2_tiehi \shift_storage.storage[679]$_SDFFE_PN0P__1841  (.L_HI(net1841));
 sg13g2_tiehi \shift_storage.storage[67]$_SDFFE_PN0P__1842  (.L_HI(net1842));
 sg13g2_tiehi \shift_storage.storage[680]$_SDFFE_PN0P__1843  (.L_HI(net1843));
 sg13g2_tiehi \shift_storage.storage[681]$_SDFFE_PN0P__1844  (.L_HI(net1844));
 sg13g2_tiehi \shift_storage.storage[682]$_SDFFE_PN0P__1845  (.L_HI(net1845));
 sg13g2_tiehi \shift_storage.storage[683]$_SDFFE_PN0P__1846  (.L_HI(net1846));
 sg13g2_tiehi \shift_storage.storage[684]$_SDFFE_PN0P__1847  (.L_HI(net1847));
 sg13g2_tiehi \shift_storage.storage[685]$_SDFFE_PN0P__1848  (.L_HI(net1848));
 sg13g2_tiehi \shift_storage.storage[686]$_SDFFE_PN0P__1849  (.L_HI(net1849));
 sg13g2_tiehi \shift_storage.storage[687]$_SDFFE_PN0P__1850  (.L_HI(net1850));
 sg13g2_tiehi \shift_storage.storage[688]$_SDFFE_PN0P__1851  (.L_HI(net1851));
 sg13g2_tiehi \shift_storage.storage[689]$_SDFFE_PN0P__1852  (.L_HI(net1852));
 sg13g2_tiehi \shift_storage.storage[68]$_SDFFE_PN0P__1853  (.L_HI(net1853));
 sg13g2_tiehi \shift_storage.storage[690]$_SDFFE_PN0P__1854  (.L_HI(net1854));
 sg13g2_tiehi \shift_storage.storage[691]$_SDFFE_PN0P__1855  (.L_HI(net1855));
 sg13g2_tiehi \shift_storage.storage[692]$_SDFFE_PN0P__1856  (.L_HI(net1856));
 sg13g2_tiehi \shift_storage.storage[693]$_SDFFE_PN0P__1857  (.L_HI(net1857));
 sg13g2_tiehi \shift_storage.storage[694]$_SDFFE_PN0P__1858  (.L_HI(net1858));
 sg13g2_tiehi \shift_storage.storage[695]$_SDFFE_PN0P__1859  (.L_HI(net1859));
 sg13g2_tiehi \shift_storage.storage[696]$_SDFFE_PN0P__1860  (.L_HI(net1860));
 sg13g2_tiehi \shift_storage.storage[697]$_SDFFE_PN0P__1861  (.L_HI(net1861));
 sg13g2_tiehi \shift_storage.storage[698]$_SDFFE_PN0P__1862  (.L_HI(net1862));
 sg13g2_tiehi \shift_storage.storage[699]$_SDFFE_PN0P__1863  (.L_HI(net1863));
 sg13g2_tiehi \shift_storage.storage[69]$_SDFFE_PN0P__1864  (.L_HI(net1864));
 sg13g2_tiehi \shift_storage.storage[6]$_SDFFE_PN0P__1865  (.L_HI(net1865));
 sg13g2_tiehi \shift_storage.storage[700]$_SDFFE_PN0P__1866  (.L_HI(net1866));
 sg13g2_tiehi \shift_storage.storage[701]$_SDFFE_PN0P__1867  (.L_HI(net1867));
 sg13g2_tiehi \shift_storage.storage[702]$_SDFFE_PN0P__1868  (.L_HI(net1868));
 sg13g2_tiehi \shift_storage.storage[703]$_SDFFE_PN0P__1869  (.L_HI(net1869));
 sg13g2_tiehi \shift_storage.storage[704]$_SDFFE_PN0P__1870  (.L_HI(net1870));
 sg13g2_tiehi \shift_storage.storage[705]$_SDFFE_PN0P__1871  (.L_HI(net1871));
 sg13g2_tiehi \shift_storage.storage[706]$_SDFFE_PN0P__1872  (.L_HI(net1872));
 sg13g2_tiehi \shift_storage.storage[707]$_SDFFE_PN0P__1873  (.L_HI(net1873));
 sg13g2_tiehi \shift_storage.storage[708]$_SDFFE_PN0P__1874  (.L_HI(net1874));
 sg13g2_tiehi \shift_storage.storage[709]$_SDFFE_PN0P__1875  (.L_HI(net1875));
 sg13g2_tiehi \shift_storage.storage[70]$_SDFFE_PN0P__1876  (.L_HI(net1876));
 sg13g2_tiehi \shift_storage.storage[710]$_SDFFE_PN0P__1877  (.L_HI(net1877));
 sg13g2_tiehi \shift_storage.storage[711]$_SDFFE_PN0P__1878  (.L_HI(net1878));
 sg13g2_tiehi \shift_storage.storage[712]$_SDFFE_PN0P__1879  (.L_HI(net1879));
 sg13g2_tiehi \shift_storage.storage[713]$_SDFFE_PN0P__1880  (.L_HI(net1880));
 sg13g2_tiehi \shift_storage.storage[714]$_SDFFE_PN0P__1881  (.L_HI(net1881));
 sg13g2_tiehi \shift_storage.storage[715]$_SDFFE_PN0P__1882  (.L_HI(net1882));
 sg13g2_tiehi \shift_storage.storage[716]$_SDFFE_PN0P__1883  (.L_HI(net1883));
 sg13g2_tiehi \shift_storage.storage[717]$_SDFFE_PN0P__1884  (.L_HI(net1884));
 sg13g2_tiehi \shift_storage.storage[718]$_SDFFE_PN0P__1885  (.L_HI(net1885));
 sg13g2_tiehi \shift_storage.storage[719]$_SDFFE_PN0P__1886  (.L_HI(net1886));
 sg13g2_tiehi \shift_storage.storage[71]$_SDFFE_PN0P__1887  (.L_HI(net1887));
 sg13g2_tiehi \shift_storage.storage[720]$_SDFFE_PN0P__1888  (.L_HI(net1888));
 sg13g2_tiehi \shift_storage.storage[721]$_SDFFE_PN0P__1889  (.L_HI(net1889));
 sg13g2_tiehi \shift_storage.storage[722]$_SDFFE_PN0P__1890  (.L_HI(net1890));
 sg13g2_tiehi \shift_storage.storage[723]$_SDFFE_PN0P__1891  (.L_HI(net1891));
 sg13g2_tiehi \shift_storage.storage[724]$_SDFFE_PN0P__1892  (.L_HI(net1892));
 sg13g2_tiehi \shift_storage.storage[725]$_SDFFE_PN0P__1893  (.L_HI(net1893));
 sg13g2_tiehi \shift_storage.storage[726]$_SDFFE_PN0P__1894  (.L_HI(net1894));
 sg13g2_tiehi \shift_storage.storage[727]$_SDFFE_PN0P__1895  (.L_HI(net1895));
 sg13g2_tiehi \shift_storage.storage[728]$_SDFFE_PN0P__1896  (.L_HI(net1896));
 sg13g2_tiehi \shift_storage.storage[729]$_SDFFE_PN0P__1897  (.L_HI(net1897));
 sg13g2_tiehi \shift_storage.storage[72]$_SDFFE_PN0P__1898  (.L_HI(net1898));
 sg13g2_tiehi \shift_storage.storage[730]$_SDFFE_PN0P__1899  (.L_HI(net1899));
 sg13g2_tiehi \shift_storage.storage[731]$_SDFFE_PN0P__1900  (.L_HI(net1900));
 sg13g2_tiehi \shift_storage.storage[732]$_SDFFE_PN0P__1901  (.L_HI(net1901));
 sg13g2_tiehi \shift_storage.storage[733]$_SDFFE_PN0P__1902  (.L_HI(net1902));
 sg13g2_tiehi \shift_storage.storage[734]$_SDFFE_PN0P__1903  (.L_HI(net1903));
 sg13g2_tiehi \shift_storage.storage[735]$_SDFFE_PN0P__1904  (.L_HI(net1904));
 sg13g2_tiehi \shift_storage.storage[736]$_SDFFE_PN0P__1905  (.L_HI(net1905));
 sg13g2_tiehi \shift_storage.storage[737]$_SDFFE_PN0P__1906  (.L_HI(net1906));
 sg13g2_tiehi \shift_storage.storage[738]$_SDFFE_PN0P__1907  (.L_HI(net1907));
 sg13g2_tiehi \shift_storage.storage[739]$_SDFFE_PN0P__1908  (.L_HI(net1908));
 sg13g2_tiehi \shift_storage.storage[73]$_SDFFE_PN0P__1909  (.L_HI(net1909));
 sg13g2_tiehi \shift_storage.storage[740]$_SDFFE_PN0P__1910  (.L_HI(net1910));
 sg13g2_tiehi \shift_storage.storage[741]$_SDFFE_PN0P__1911  (.L_HI(net1911));
 sg13g2_tiehi \shift_storage.storage[742]$_SDFFE_PN0P__1912  (.L_HI(net1912));
 sg13g2_tiehi \shift_storage.storage[743]$_SDFFE_PN0P__1913  (.L_HI(net1913));
 sg13g2_tiehi \shift_storage.storage[744]$_SDFFE_PN0P__1914  (.L_HI(net1914));
 sg13g2_tiehi \shift_storage.storage[745]$_SDFFE_PN0P__1915  (.L_HI(net1915));
 sg13g2_tiehi \shift_storage.storage[746]$_SDFFE_PN0P__1916  (.L_HI(net1916));
 sg13g2_tiehi \shift_storage.storage[747]$_SDFFE_PN0P__1917  (.L_HI(net1917));
 sg13g2_tiehi \shift_storage.storage[748]$_SDFFE_PN0P__1918  (.L_HI(net1918));
 sg13g2_tiehi \shift_storage.storage[749]$_SDFFE_PN0P__1919  (.L_HI(net1919));
 sg13g2_tiehi \shift_storage.storage[74]$_SDFFE_PN0P__1920  (.L_HI(net1920));
 sg13g2_tiehi \shift_storage.storage[750]$_SDFFE_PN0P__1921  (.L_HI(net1921));
 sg13g2_tiehi \shift_storage.storage[751]$_SDFFE_PN0P__1922  (.L_HI(net1922));
 sg13g2_tiehi \shift_storage.storage[752]$_SDFFE_PN0P__1923  (.L_HI(net1923));
 sg13g2_tiehi \shift_storage.storage[753]$_SDFFE_PN0P__1924  (.L_HI(net1924));
 sg13g2_tiehi \shift_storage.storage[754]$_SDFFE_PN0P__1925  (.L_HI(net1925));
 sg13g2_tiehi \shift_storage.storage[755]$_SDFFE_PN0P__1926  (.L_HI(net1926));
 sg13g2_tiehi \shift_storage.storage[756]$_SDFFE_PN0P__1927  (.L_HI(net1927));
 sg13g2_tiehi \shift_storage.storage[757]$_SDFFE_PN0P__1928  (.L_HI(net1928));
 sg13g2_tiehi \shift_storage.storage[758]$_SDFFE_PN0P__1929  (.L_HI(net1929));
 sg13g2_tiehi \shift_storage.storage[759]$_SDFFE_PN0P__1930  (.L_HI(net1930));
 sg13g2_tiehi \shift_storage.storage[75]$_SDFFE_PN0P__1931  (.L_HI(net1931));
 sg13g2_tiehi \shift_storage.storage[760]$_SDFFE_PN0P__1932  (.L_HI(net1932));
 sg13g2_tiehi \shift_storage.storage[761]$_SDFFE_PN0P__1933  (.L_HI(net1933));
 sg13g2_tiehi \shift_storage.storage[762]$_SDFFE_PN0P__1934  (.L_HI(net1934));
 sg13g2_tiehi \shift_storage.storage[763]$_SDFFE_PN0P__1935  (.L_HI(net1935));
 sg13g2_tiehi \shift_storage.storage[764]$_SDFFE_PN0P__1936  (.L_HI(net1936));
 sg13g2_tiehi \shift_storage.storage[765]$_SDFFE_PN0P__1937  (.L_HI(net1937));
 sg13g2_tiehi \shift_storage.storage[766]$_SDFFE_PN0P__1938  (.L_HI(net1938));
 sg13g2_tiehi \shift_storage.storage[767]$_SDFFE_PN0P__1939  (.L_HI(net1939));
 sg13g2_tiehi \shift_storage.storage[768]$_SDFFE_PN0P__1940  (.L_HI(net1940));
 sg13g2_tiehi \shift_storage.storage[769]$_SDFFE_PN0P__1941  (.L_HI(net1941));
 sg13g2_tiehi \shift_storage.storage[76]$_SDFFE_PN0P__1942  (.L_HI(net1942));
 sg13g2_tiehi \shift_storage.storage[770]$_SDFFE_PN0P__1943  (.L_HI(net1943));
 sg13g2_tiehi \shift_storage.storage[771]$_SDFFE_PN0P__1944  (.L_HI(net1944));
 sg13g2_tiehi \shift_storage.storage[772]$_SDFFE_PN0P__1945  (.L_HI(net1945));
 sg13g2_tiehi \shift_storage.storage[773]$_SDFFE_PN0P__1946  (.L_HI(net1946));
 sg13g2_tiehi \shift_storage.storage[774]$_SDFFE_PN0P__1947  (.L_HI(net1947));
 sg13g2_tiehi \shift_storage.storage[775]$_SDFFE_PN0P__1948  (.L_HI(net1948));
 sg13g2_tiehi \shift_storage.storage[776]$_SDFFE_PN0P__1949  (.L_HI(net1949));
 sg13g2_tiehi \shift_storage.storage[777]$_SDFFE_PN0P__1950  (.L_HI(net1950));
 sg13g2_tiehi \shift_storage.storage[778]$_SDFFE_PN0P__1951  (.L_HI(net1951));
 sg13g2_tiehi \shift_storage.storage[779]$_SDFFE_PN0P__1952  (.L_HI(net1952));
 sg13g2_tiehi \shift_storage.storage[77]$_SDFFE_PN0P__1953  (.L_HI(net1953));
 sg13g2_tiehi \shift_storage.storage[780]$_SDFFE_PN0P__1954  (.L_HI(net1954));
 sg13g2_tiehi \shift_storage.storage[781]$_SDFFE_PN0P__1955  (.L_HI(net1955));
 sg13g2_tiehi \shift_storage.storage[782]$_SDFFE_PN0P__1956  (.L_HI(net1956));
 sg13g2_tiehi \shift_storage.storage[783]$_SDFFE_PN0P__1957  (.L_HI(net1957));
 sg13g2_tiehi \shift_storage.storage[784]$_SDFFE_PN0P__1958  (.L_HI(net1958));
 sg13g2_tiehi \shift_storage.storage[785]$_SDFFE_PN0P__1959  (.L_HI(net1959));
 sg13g2_tiehi \shift_storage.storage[786]$_SDFFE_PN0P__1960  (.L_HI(net1960));
 sg13g2_tiehi \shift_storage.storage[787]$_SDFFE_PN0P__1961  (.L_HI(net1961));
 sg13g2_tiehi \shift_storage.storage[788]$_SDFFE_PN0P__1962  (.L_HI(net1962));
 sg13g2_tiehi \shift_storage.storage[789]$_SDFFE_PN0P__1963  (.L_HI(net1963));
 sg13g2_tiehi \shift_storage.storage[78]$_SDFFE_PN0P__1964  (.L_HI(net1964));
 sg13g2_tiehi \shift_storage.storage[790]$_SDFFE_PN0P__1965  (.L_HI(net1965));
 sg13g2_tiehi \shift_storage.storage[791]$_SDFFE_PN0P__1966  (.L_HI(net1966));
 sg13g2_tiehi \shift_storage.storage[792]$_SDFFE_PN0P__1967  (.L_HI(net1967));
 sg13g2_tiehi \shift_storage.storage[793]$_SDFFE_PN0P__1968  (.L_HI(net1968));
 sg13g2_tiehi \shift_storage.storage[794]$_SDFFE_PN0P__1969  (.L_HI(net1969));
 sg13g2_tiehi \shift_storage.storage[795]$_SDFFE_PN0P__1970  (.L_HI(net1970));
 sg13g2_tiehi \shift_storage.storage[796]$_SDFFE_PN0P__1971  (.L_HI(net1971));
 sg13g2_tiehi \shift_storage.storage[797]$_SDFFE_PN0P__1972  (.L_HI(net1972));
 sg13g2_tiehi \shift_storage.storage[798]$_SDFFE_PN0P__1973  (.L_HI(net1973));
 sg13g2_tiehi \shift_storage.storage[799]$_SDFFE_PN0P__1974  (.L_HI(net1974));
 sg13g2_tiehi \shift_storage.storage[79]$_SDFFE_PN0P__1975  (.L_HI(net1975));
 sg13g2_tiehi \shift_storage.storage[7]$_SDFFE_PN0P__1976  (.L_HI(net1976));
 sg13g2_tiehi \shift_storage.storage[800]$_SDFFE_PN0P__1977  (.L_HI(net1977));
 sg13g2_tiehi \shift_storage.storage[801]$_SDFFE_PN0P__1978  (.L_HI(net1978));
 sg13g2_tiehi \shift_storage.storage[802]$_SDFFE_PN0P__1979  (.L_HI(net1979));
 sg13g2_tiehi \shift_storage.storage[803]$_SDFFE_PN0P__1980  (.L_HI(net1980));
 sg13g2_tiehi \shift_storage.storage[804]$_SDFFE_PN0P__1981  (.L_HI(net1981));
 sg13g2_tiehi \shift_storage.storage[805]$_SDFFE_PN0P__1982  (.L_HI(net1982));
 sg13g2_tiehi \shift_storage.storage[806]$_SDFFE_PN0P__1983  (.L_HI(net1983));
 sg13g2_tiehi \shift_storage.storage[807]$_SDFFE_PN0P__1984  (.L_HI(net1984));
 sg13g2_tiehi \shift_storage.storage[808]$_SDFFE_PN0P__1985  (.L_HI(net1985));
 sg13g2_tiehi \shift_storage.storage[809]$_SDFFE_PN0P__1986  (.L_HI(net1986));
 sg13g2_tiehi \shift_storage.storage[80]$_SDFFE_PN0P__1987  (.L_HI(net1987));
 sg13g2_tiehi \shift_storage.storage[810]$_SDFFE_PN0P__1988  (.L_HI(net1988));
 sg13g2_tiehi \shift_storage.storage[811]$_SDFFE_PN0P__1989  (.L_HI(net1989));
 sg13g2_tiehi \shift_storage.storage[812]$_SDFFE_PN0P__1990  (.L_HI(net1990));
 sg13g2_tiehi \shift_storage.storage[813]$_SDFFE_PN0P__1991  (.L_HI(net1991));
 sg13g2_tiehi \shift_storage.storage[814]$_SDFFE_PN0P__1992  (.L_HI(net1992));
 sg13g2_tiehi \shift_storage.storage[815]$_SDFFE_PN0P__1993  (.L_HI(net1993));
 sg13g2_tiehi \shift_storage.storage[816]$_SDFFE_PN0P__1994  (.L_HI(net1994));
 sg13g2_tiehi \shift_storage.storage[817]$_SDFFE_PN0P__1995  (.L_HI(net1995));
 sg13g2_tiehi \shift_storage.storage[818]$_SDFFE_PN0P__1996  (.L_HI(net1996));
 sg13g2_tiehi \shift_storage.storage[819]$_SDFFE_PN0P__1997  (.L_HI(net1997));
 sg13g2_tiehi \shift_storage.storage[81]$_SDFFE_PN0P__1998  (.L_HI(net1998));
 sg13g2_tiehi \shift_storage.storage[820]$_SDFFE_PN0P__1999  (.L_HI(net1999));
 sg13g2_tiehi \shift_storage.storage[821]$_SDFFE_PN0P__2000  (.L_HI(net2000));
 sg13g2_tiehi \shift_storage.storage[822]$_SDFFE_PN0P__2001  (.L_HI(net2001));
 sg13g2_tiehi \shift_storage.storage[823]$_SDFFE_PN0P__2002  (.L_HI(net2002));
 sg13g2_tiehi \shift_storage.storage[824]$_SDFFE_PN0P__2003  (.L_HI(net2003));
 sg13g2_tiehi \shift_storage.storage[825]$_SDFFE_PN0P__2004  (.L_HI(net2004));
 sg13g2_tiehi \shift_storage.storage[826]$_SDFFE_PN0P__2005  (.L_HI(net2005));
 sg13g2_tiehi \shift_storage.storage[827]$_SDFFE_PN0P__2006  (.L_HI(net2006));
 sg13g2_tiehi \shift_storage.storage[828]$_SDFFE_PN0P__2007  (.L_HI(net2007));
 sg13g2_tiehi \shift_storage.storage[829]$_SDFFE_PN0P__2008  (.L_HI(net2008));
 sg13g2_tiehi \shift_storage.storage[82]$_SDFFE_PN0P__2009  (.L_HI(net2009));
 sg13g2_tiehi \shift_storage.storage[830]$_SDFFE_PN0P__2010  (.L_HI(net2010));
 sg13g2_tiehi \shift_storage.storage[831]$_SDFFE_PN0P__2011  (.L_HI(net2011));
 sg13g2_tiehi \shift_storage.storage[832]$_SDFFE_PN0P__2012  (.L_HI(net2012));
 sg13g2_tiehi \shift_storage.storage[833]$_SDFFE_PN0P__2013  (.L_HI(net2013));
 sg13g2_tiehi \shift_storage.storage[834]$_SDFFE_PN0P__2014  (.L_HI(net2014));
 sg13g2_tiehi \shift_storage.storage[835]$_SDFFE_PN0P__2015  (.L_HI(net2015));
 sg13g2_tiehi \shift_storage.storage[836]$_SDFFE_PN0P__2016  (.L_HI(net2016));
 sg13g2_tiehi \shift_storage.storage[837]$_SDFFE_PN0P__2017  (.L_HI(net2017));
 sg13g2_tiehi \shift_storage.storage[838]$_SDFFE_PN0P__2018  (.L_HI(net2018));
 sg13g2_tiehi \shift_storage.storage[839]$_SDFFE_PN0P__2019  (.L_HI(net2019));
 sg13g2_tiehi \shift_storage.storage[83]$_SDFFE_PN0P__2020  (.L_HI(net2020));
 sg13g2_tiehi \shift_storage.storage[840]$_SDFFE_PN0P__2021  (.L_HI(net2021));
 sg13g2_tiehi \shift_storage.storage[841]$_SDFFE_PN0P__2022  (.L_HI(net2022));
 sg13g2_tiehi \shift_storage.storage[842]$_SDFFE_PN0P__2023  (.L_HI(net2023));
 sg13g2_tiehi \shift_storage.storage[843]$_SDFFE_PN0P__2024  (.L_HI(net2024));
 sg13g2_tiehi \shift_storage.storage[844]$_SDFFE_PN0P__2025  (.L_HI(net2025));
 sg13g2_tiehi \shift_storage.storage[845]$_SDFFE_PN0P__2026  (.L_HI(net2026));
 sg13g2_tiehi \shift_storage.storage[846]$_SDFFE_PN0P__2027  (.L_HI(net2027));
 sg13g2_tiehi \shift_storage.storage[847]$_SDFFE_PN0P__2028  (.L_HI(net2028));
 sg13g2_tiehi \shift_storage.storage[848]$_SDFFE_PN0P__2029  (.L_HI(net2029));
 sg13g2_tiehi \shift_storage.storage[849]$_SDFFE_PN0P__2030  (.L_HI(net2030));
 sg13g2_tiehi \shift_storage.storage[84]$_SDFFE_PN0P__2031  (.L_HI(net2031));
 sg13g2_tiehi \shift_storage.storage[850]$_SDFFE_PN0P__2032  (.L_HI(net2032));
 sg13g2_tiehi \shift_storage.storage[851]$_SDFFE_PN0P__2033  (.L_HI(net2033));
 sg13g2_tiehi \shift_storage.storage[852]$_SDFFE_PN0P__2034  (.L_HI(net2034));
 sg13g2_tiehi \shift_storage.storage[853]$_SDFFE_PN0P__2035  (.L_HI(net2035));
 sg13g2_tiehi \shift_storage.storage[854]$_SDFFE_PN0P__2036  (.L_HI(net2036));
 sg13g2_tiehi \shift_storage.storage[855]$_SDFFE_PN0P__2037  (.L_HI(net2037));
 sg13g2_tiehi \shift_storage.storage[856]$_SDFFE_PN0P__2038  (.L_HI(net2038));
 sg13g2_tiehi \shift_storage.storage[857]$_SDFFE_PN0P__2039  (.L_HI(net2039));
 sg13g2_tiehi \shift_storage.storage[858]$_SDFFE_PN0P__2040  (.L_HI(net2040));
 sg13g2_tiehi \shift_storage.storage[859]$_SDFFE_PN0P__2041  (.L_HI(net2041));
 sg13g2_tiehi \shift_storage.storage[85]$_SDFFE_PN0P__2042  (.L_HI(net2042));
 sg13g2_tiehi \shift_storage.storage[860]$_SDFFE_PN0P__2043  (.L_HI(net2043));
 sg13g2_tiehi \shift_storage.storage[861]$_SDFFE_PN0P__2044  (.L_HI(net2044));
 sg13g2_tiehi \shift_storage.storage[862]$_SDFFE_PN0P__2045  (.L_HI(net2045));
 sg13g2_tiehi \shift_storage.storage[863]$_SDFFE_PN0P__2046  (.L_HI(net2046));
 sg13g2_tiehi \shift_storage.storage[864]$_SDFFE_PN0P__2047  (.L_HI(net2047));
 sg13g2_tiehi \shift_storage.storage[865]$_SDFFE_PN0P__2048  (.L_HI(net2048));
 sg13g2_tiehi \shift_storage.storage[866]$_SDFFE_PN0P__2049  (.L_HI(net2049));
 sg13g2_tiehi \shift_storage.storage[867]$_SDFFE_PN0P__2050  (.L_HI(net2050));
 sg13g2_tiehi \shift_storage.storage[868]$_SDFFE_PN0P__2051  (.L_HI(net2051));
 sg13g2_tiehi \shift_storage.storage[869]$_SDFFE_PN0P__2052  (.L_HI(net2052));
 sg13g2_tiehi \shift_storage.storage[86]$_SDFFE_PN0P__2053  (.L_HI(net2053));
 sg13g2_tiehi \shift_storage.storage[870]$_SDFFE_PN0P__2054  (.L_HI(net2054));
 sg13g2_tiehi \shift_storage.storage[871]$_SDFFE_PN0P__2055  (.L_HI(net2055));
 sg13g2_tiehi \shift_storage.storage[872]$_SDFFE_PN0P__2056  (.L_HI(net2056));
 sg13g2_tiehi \shift_storage.storage[873]$_SDFFE_PN0P__2057  (.L_HI(net2057));
 sg13g2_tiehi \shift_storage.storage[874]$_SDFFE_PN0P__2058  (.L_HI(net2058));
 sg13g2_tiehi \shift_storage.storage[875]$_SDFFE_PN0P__2059  (.L_HI(net2059));
 sg13g2_tiehi \shift_storage.storage[876]$_SDFFE_PN0P__2060  (.L_HI(net2060));
 sg13g2_tiehi \shift_storage.storage[877]$_SDFFE_PN0P__2061  (.L_HI(net2061));
 sg13g2_tiehi \shift_storage.storage[878]$_SDFFE_PN0P__2062  (.L_HI(net2062));
 sg13g2_tiehi \shift_storage.storage[879]$_SDFFE_PN0P__2063  (.L_HI(net2063));
 sg13g2_tiehi \shift_storage.storage[87]$_SDFFE_PN0P__2064  (.L_HI(net2064));
 sg13g2_tiehi \shift_storage.storage[880]$_SDFFE_PN0P__2065  (.L_HI(net2065));
 sg13g2_tiehi \shift_storage.storage[881]$_SDFFE_PN0P__2066  (.L_HI(net2066));
 sg13g2_tiehi \shift_storage.storage[882]$_SDFFE_PN0P__2067  (.L_HI(net2067));
 sg13g2_tiehi \shift_storage.storage[883]$_SDFFE_PN0P__2068  (.L_HI(net2068));
 sg13g2_tiehi \shift_storage.storage[884]$_SDFFE_PN0P__2069  (.L_HI(net2069));
 sg13g2_tiehi \shift_storage.storage[885]$_SDFFE_PN0P__2070  (.L_HI(net2070));
 sg13g2_tiehi \shift_storage.storage[886]$_SDFFE_PN0P__2071  (.L_HI(net2071));
 sg13g2_tiehi \shift_storage.storage[887]$_SDFFE_PN0P__2072  (.L_HI(net2072));
 sg13g2_tiehi \shift_storage.storage[888]$_SDFFE_PN0P__2073  (.L_HI(net2073));
 sg13g2_tiehi \shift_storage.storage[889]$_SDFFE_PN0P__2074  (.L_HI(net2074));
 sg13g2_tiehi \shift_storage.storage[88]$_SDFFE_PN0P__2075  (.L_HI(net2075));
 sg13g2_tiehi \shift_storage.storage[890]$_SDFFE_PN0P__2076  (.L_HI(net2076));
 sg13g2_tiehi \shift_storage.storage[891]$_SDFFE_PN0P__2077  (.L_HI(net2077));
 sg13g2_tiehi \shift_storage.storage[892]$_SDFFE_PN0P__2078  (.L_HI(net2078));
 sg13g2_tiehi \shift_storage.storage[893]$_SDFFE_PN0P__2079  (.L_HI(net2079));
 sg13g2_tiehi \shift_storage.storage[894]$_SDFFE_PN0P__2080  (.L_HI(net2080));
 sg13g2_tiehi \shift_storage.storage[895]$_SDFFE_PN0P__2081  (.L_HI(net2081));
 sg13g2_tiehi \shift_storage.storage[896]$_SDFFE_PN0P__2082  (.L_HI(net2082));
 sg13g2_tiehi \shift_storage.storage[897]$_SDFFE_PN0P__2083  (.L_HI(net2083));
 sg13g2_tiehi \shift_storage.storage[898]$_SDFFE_PN0P__2084  (.L_HI(net2084));
 sg13g2_tiehi \shift_storage.storage[899]$_SDFFE_PN0P__2085  (.L_HI(net2085));
 sg13g2_tiehi \shift_storage.storage[89]$_SDFFE_PN0P__2086  (.L_HI(net2086));
 sg13g2_tiehi \shift_storage.storage[8]$_SDFFE_PN0P__2087  (.L_HI(net2087));
 sg13g2_tiehi \shift_storage.storage[900]$_SDFFE_PN0P__2088  (.L_HI(net2088));
 sg13g2_tiehi \shift_storage.storage[901]$_SDFFE_PN0P__2089  (.L_HI(net2089));
 sg13g2_tiehi \shift_storage.storage[902]$_SDFFE_PN0P__2090  (.L_HI(net2090));
 sg13g2_tiehi \shift_storage.storage[903]$_SDFFE_PN0P__2091  (.L_HI(net2091));
 sg13g2_tiehi \shift_storage.storage[904]$_SDFFE_PN0P__2092  (.L_HI(net2092));
 sg13g2_tiehi \shift_storage.storage[905]$_SDFFE_PN0P__2093  (.L_HI(net2093));
 sg13g2_tiehi \shift_storage.storage[906]$_SDFFE_PN0P__2094  (.L_HI(net2094));
 sg13g2_tiehi \shift_storage.storage[907]$_SDFFE_PN0P__2095  (.L_HI(net2095));
 sg13g2_tiehi \shift_storage.storage[908]$_SDFFE_PN0P__2096  (.L_HI(net2096));
 sg13g2_tiehi \shift_storage.storage[909]$_SDFFE_PN0P__2097  (.L_HI(net2097));
 sg13g2_tiehi \shift_storage.storage[90]$_SDFFE_PN0P__2098  (.L_HI(net2098));
 sg13g2_tiehi \shift_storage.storage[910]$_SDFFE_PN0P__2099  (.L_HI(net2099));
 sg13g2_tiehi \shift_storage.storage[911]$_SDFFE_PN0P__2100  (.L_HI(net2100));
 sg13g2_tiehi \shift_storage.storage[912]$_SDFFE_PN0P__2101  (.L_HI(net2101));
 sg13g2_tiehi \shift_storage.storage[913]$_SDFFE_PN0P__2102  (.L_HI(net2102));
 sg13g2_tiehi \shift_storage.storage[914]$_SDFFE_PN0P__2103  (.L_HI(net2103));
 sg13g2_tiehi \shift_storage.storage[915]$_SDFFE_PN0P__2104  (.L_HI(net2104));
 sg13g2_tiehi \shift_storage.storage[916]$_SDFFE_PN0P__2105  (.L_HI(net2105));
 sg13g2_tiehi \shift_storage.storage[917]$_SDFFE_PN0P__2106  (.L_HI(net2106));
 sg13g2_tiehi \shift_storage.storage[918]$_SDFFE_PN0P__2107  (.L_HI(net2107));
 sg13g2_tiehi \shift_storage.storage[919]$_SDFFE_PN0P__2108  (.L_HI(net2108));
 sg13g2_tiehi \shift_storage.storage[91]$_SDFFE_PN0P__2109  (.L_HI(net2109));
 sg13g2_tiehi \shift_storage.storage[920]$_SDFFE_PN0P__2110  (.L_HI(net2110));
 sg13g2_tiehi \shift_storage.storage[921]$_SDFFE_PN0P__2111  (.L_HI(net2111));
 sg13g2_tiehi \shift_storage.storage[922]$_SDFFE_PN0P__2112  (.L_HI(net2112));
 sg13g2_tiehi \shift_storage.storage[923]$_SDFFE_PN0P__2113  (.L_HI(net2113));
 sg13g2_tiehi \shift_storage.storage[924]$_SDFFE_PN0P__2114  (.L_HI(net2114));
 sg13g2_tiehi \shift_storage.storage[925]$_SDFFE_PN0P__2115  (.L_HI(net2115));
 sg13g2_tiehi \shift_storage.storage[926]$_SDFFE_PN0P__2116  (.L_HI(net2116));
 sg13g2_tiehi \shift_storage.storage[927]$_SDFFE_PN0P__2117  (.L_HI(net2117));
 sg13g2_tiehi \shift_storage.storage[928]$_SDFFE_PN0P__2118  (.L_HI(net2118));
 sg13g2_tiehi \shift_storage.storage[929]$_SDFFE_PN0P__2119  (.L_HI(net2119));
 sg13g2_tiehi \shift_storage.storage[92]$_SDFFE_PN0P__2120  (.L_HI(net2120));
 sg13g2_tiehi \shift_storage.storage[930]$_SDFFE_PN0P__2121  (.L_HI(net2121));
 sg13g2_tiehi \shift_storage.storage[931]$_SDFFE_PN0P__2122  (.L_HI(net2122));
 sg13g2_tiehi \shift_storage.storage[932]$_SDFFE_PN0P__2123  (.L_HI(net2123));
 sg13g2_tiehi \shift_storage.storage[933]$_SDFFE_PN0P__2124  (.L_HI(net2124));
 sg13g2_tiehi \shift_storage.storage[934]$_SDFFE_PN0P__2125  (.L_HI(net2125));
 sg13g2_tiehi \shift_storage.storage[935]$_SDFFE_PN0P__2126  (.L_HI(net2126));
 sg13g2_tiehi \shift_storage.storage[936]$_SDFFE_PN0P__2127  (.L_HI(net2127));
 sg13g2_tiehi \shift_storage.storage[937]$_SDFFE_PN0P__2128  (.L_HI(net2128));
 sg13g2_tiehi \shift_storage.storage[938]$_SDFFE_PN0P__2129  (.L_HI(net2129));
 sg13g2_tiehi \shift_storage.storage[939]$_SDFFE_PN0P__2130  (.L_HI(net2130));
 sg13g2_tiehi \shift_storage.storage[93]$_SDFFE_PN0P__2131  (.L_HI(net2131));
 sg13g2_tiehi \shift_storage.storage[940]$_SDFFE_PN0P__2132  (.L_HI(net2132));
 sg13g2_tiehi \shift_storage.storage[941]$_SDFFE_PN0P__2133  (.L_HI(net2133));
 sg13g2_tiehi \shift_storage.storage[942]$_SDFFE_PN0P__2134  (.L_HI(net2134));
 sg13g2_tiehi \shift_storage.storage[943]$_SDFFE_PN0P__2135  (.L_HI(net2135));
 sg13g2_tiehi \shift_storage.storage[944]$_SDFFE_PN0P__2136  (.L_HI(net2136));
 sg13g2_tiehi \shift_storage.storage[945]$_SDFFE_PN0P__2137  (.L_HI(net2137));
 sg13g2_tiehi \shift_storage.storage[946]$_SDFFE_PN0P__2138  (.L_HI(net2138));
 sg13g2_tiehi \shift_storage.storage[947]$_SDFFE_PN0P__2139  (.L_HI(net2139));
 sg13g2_tiehi \shift_storage.storage[948]$_SDFFE_PN0P__2140  (.L_HI(net2140));
 sg13g2_tiehi \shift_storage.storage[949]$_SDFFE_PN0P__2141  (.L_HI(net2141));
 sg13g2_tiehi \shift_storage.storage[94]$_SDFFE_PN0P__2142  (.L_HI(net2142));
 sg13g2_tiehi \shift_storage.storage[950]$_SDFFE_PN0P__2143  (.L_HI(net2143));
 sg13g2_tiehi \shift_storage.storage[951]$_SDFFE_PN0P__2144  (.L_HI(net2144));
 sg13g2_tiehi \shift_storage.storage[952]$_SDFFE_PN0P__2145  (.L_HI(net2145));
 sg13g2_tiehi \shift_storage.storage[953]$_SDFFE_PN0P__2146  (.L_HI(net2146));
 sg13g2_tiehi \shift_storage.storage[954]$_SDFFE_PN0P__2147  (.L_HI(net2147));
 sg13g2_tiehi \shift_storage.storage[955]$_SDFFE_PN0P__2148  (.L_HI(net2148));
 sg13g2_tiehi \shift_storage.storage[956]$_SDFFE_PN0P__2149  (.L_HI(net2149));
 sg13g2_tiehi \shift_storage.storage[957]$_SDFFE_PN0P__2150  (.L_HI(net2150));
 sg13g2_tiehi \shift_storage.storage[958]$_SDFFE_PN0P__2151  (.L_HI(net2151));
 sg13g2_tiehi \shift_storage.storage[959]$_SDFFE_PN0P__2152  (.L_HI(net2152));
 sg13g2_tiehi \shift_storage.storage[95]$_SDFFE_PN0P__2153  (.L_HI(net2153));
 sg13g2_tiehi \shift_storage.storage[960]$_SDFFE_PN0P__2154  (.L_HI(net2154));
 sg13g2_tiehi \shift_storage.storage[961]$_SDFFE_PN0P__2155  (.L_HI(net2155));
 sg13g2_tiehi \shift_storage.storage[962]$_SDFFE_PN0P__2156  (.L_HI(net2156));
 sg13g2_tiehi \shift_storage.storage[963]$_SDFFE_PN0P__2157  (.L_HI(net2157));
 sg13g2_tiehi \shift_storage.storage[964]$_SDFFE_PN0P__2158  (.L_HI(net2158));
 sg13g2_tiehi \shift_storage.storage[965]$_SDFFE_PN0P__2159  (.L_HI(net2159));
 sg13g2_tiehi \shift_storage.storage[966]$_SDFFE_PN0P__2160  (.L_HI(net2160));
 sg13g2_tiehi \shift_storage.storage[967]$_SDFFE_PN0P__2161  (.L_HI(net2161));
 sg13g2_tiehi \shift_storage.storage[968]$_SDFFE_PN0P__2162  (.L_HI(net2162));
 sg13g2_tiehi \shift_storage.storage[969]$_SDFFE_PN0P__2163  (.L_HI(net2163));
 sg13g2_tiehi \shift_storage.storage[96]$_SDFFE_PN0P__2164  (.L_HI(net2164));
 sg13g2_tiehi \shift_storage.storage[970]$_SDFFE_PN0P__2165  (.L_HI(net2165));
 sg13g2_tiehi \shift_storage.storage[971]$_SDFFE_PN0P__2166  (.L_HI(net2166));
 sg13g2_tiehi \shift_storage.storage[972]$_SDFFE_PN0P__2167  (.L_HI(net2167));
 sg13g2_tiehi \shift_storage.storage[973]$_SDFFE_PN0P__2168  (.L_HI(net2168));
 sg13g2_tiehi \shift_storage.storage[974]$_SDFFE_PN0P__2169  (.L_HI(net2169));
 sg13g2_tiehi \shift_storage.storage[975]$_SDFFE_PN0P__2170  (.L_HI(net2170));
 sg13g2_tiehi \shift_storage.storage[976]$_SDFFE_PN0P__2171  (.L_HI(net2171));
 sg13g2_tiehi \shift_storage.storage[977]$_SDFFE_PN0P__2172  (.L_HI(net2172));
 sg13g2_tiehi \shift_storage.storage[978]$_SDFFE_PN0P__2173  (.L_HI(net2173));
 sg13g2_tiehi \shift_storage.storage[979]$_SDFFE_PN0P__2174  (.L_HI(net2174));
 sg13g2_tiehi \shift_storage.storage[97]$_SDFFE_PN0P__2175  (.L_HI(net2175));
 sg13g2_tiehi \shift_storage.storage[980]$_SDFFE_PN0P__2176  (.L_HI(net2176));
 sg13g2_tiehi \shift_storage.storage[981]$_SDFFE_PN0P__2177  (.L_HI(net2177));
 sg13g2_tiehi \shift_storage.storage[982]$_SDFFE_PN0P__2178  (.L_HI(net2178));
 sg13g2_tiehi \shift_storage.storage[983]$_SDFFE_PN0P__2179  (.L_HI(net2179));
 sg13g2_tiehi \shift_storage.storage[984]$_SDFFE_PN0P__2180  (.L_HI(net2180));
 sg13g2_tiehi \shift_storage.storage[985]$_SDFFE_PN0P__2181  (.L_HI(net2181));
 sg13g2_tiehi \shift_storage.storage[986]$_SDFFE_PN0P__2182  (.L_HI(net2182));
 sg13g2_tiehi \shift_storage.storage[987]$_SDFFE_PN0P__2183  (.L_HI(net2183));
 sg13g2_tiehi \shift_storage.storage[988]$_SDFFE_PN0P__2184  (.L_HI(net2184));
 sg13g2_tiehi \shift_storage.storage[989]$_SDFFE_PN0P__2185  (.L_HI(net2185));
 sg13g2_tiehi \shift_storage.storage[98]$_SDFFE_PN0P__2186  (.L_HI(net2186));
 sg13g2_tiehi \shift_storage.storage[990]$_SDFFE_PN0P__2187  (.L_HI(net2187));
 sg13g2_tiehi \shift_storage.storage[991]$_SDFFE_PN0P__2188  (.L_HI(net2188));
 sg13g2_tiehi \shift_storage.storage[992]$_SDFFE_PN0P__2189  (.L_HI(net2189));
 sg13g2_tiehi \shift_storage.storage[993]$_SDFFE_PN0P__2190  (.L_HI(net2190));
 sg13g2_tiehi \shift_storage.storage[994]$_SDFFE_PN0P__2191  (.L_HI(net2191));
 sg13g2_tiehi \shift_storage.storage[995]$_SDFFE_PN0P__2192  (.L_HI(net2192));
 sg13g2_tiehi \shift_storage.storage[996]$_SDFFE_PN0P__2193  (.L_HI(net2193));
 sg13g2_tiehi \shift_storage.storage[997]$_SDFFE_PN0P__2194  (.L_HI(net2194));
 sg13g2_tiehi \shift_storage.storage[998]$_SDFFE_PN0P__2195  (.L_HI(net2195));
 sg13g2_tiehi \shift_storage.storage[999]$_SDFFE_PN0P__2196  (.L_HI(net2196));
 sg13g2_tiehi \shift_storage.storage[99]$_SDFFE_PN0P__2197  (.L_HI(net2197));
 sg13g2_tiehi \shift_storage.storage[9]$_SDFFE_PN0P__2198  (.L_HI(net2198));
 sg13g2_buf_4 clkbuf_leaf_1_clk_p2c (.X(clknet_leaf_1_clk_p2c),
    .A(clknet_5_0__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_2_clk_p2c (.X(clknet_leaf_2_clk_p2c),
    .A(clknet_5_0__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_3_clk_p2c (.X(clknet_leaf_3_clk_p2c),
    .A(clknet_5_0__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_4_clk_p2c (.X(clknet_leaf_4_clk_p2c),
    .A(clknet_5_0__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_5_clk_p2c (.X(clknet_leaf_5_clk_p2c),
    .A(clknet_5_0__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_6_clk_p2c (.X(clknet_leaf_6_clk_p2c),
    .A(clknet_5_2__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_7_clk_p2c (.X(clknet_leaf_7_clk_p2c),
    .A(clknet_5_2__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_8_clk_p2c (.X(clknet_leaf_8_clk_p2c),
    .A(clknet_5_0__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_9_clk_p2c (.X(clknet_leaf_9_clk_p2c),
    .A(clknet_5_0__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_10_clk_p2c (.X(clknet_leaf_10_clk_p2c),
    .A(clknet_5_3__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_11_clk_p2c (.X(clknet_leaf_11_clk_p2c),
    .A(clknet_5_3__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_12_clk_p2c (.X(clknet_leaf_12_clk_p2c),
    .A(clknet_5_3__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_13_clk_p2c (.X(clknet_leaf_13_clk_p2c),
    .A(clknet_5_3__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_14_clk_p2c (.X(clknet_leaf_14_clk_p2c),
    .A(clknet_5_3__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_15_clk_p2c (.X(clknet_leaf_15_clk_p2c),
    .A(clknet_5_2__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_16_clk_p2c (.X(clknet_leaf_16_clk_p2c),
    .A(clknet_5_2__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_17_clk_p2c (.X(clknet_leaf_17_clk_p2c),
    .A(clknet_5_2__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_18_clk_p2c (.X(clknet_leaf_18_clk_p2c),
    .A(clknet_5_2__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_19_clk_p2c (.X(clknet_leaf_19_clk_p2c),
    .A(clknet_5_2__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_20_clk_p2c (.X(clknet_leaf_20_clk_p2c),
    .A(clknet_5_2__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_21_clk_p2c (.X(clknet_leaf_21_clk_p2c),
    .A(clknet_5_2__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_22_clk_p2c (.X(clknet_leaf_22_clk_p2c),
    .A(clknet_5_2__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_23_clk_p2c (.X(clknet_leaf_23_clk_p2c),
    .A(clknet_5_8__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_24_clk_p2c (.X(clknet_leaf_24_clk_p2c),
    .A(clknet_5_8__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_25_clk_p2c (.X(clknet_leaf_25_clk_p2c),
    .A(clknet_5_8__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_26_clk_p2c (.X(clknet_leaf_26_clk_p2c),
    .A(clknet_5_2__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_27_clk_p2c (.X(clknet_leaf_27_clk_p2c),
    .A(clknet_5_3__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_28_clk_p2c (.X(clknet_leaf_28_clk_p2c),
    .A(clknet_5_9__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_29_clk_p2c (.X(clknet_leaf_29_clk_p2c),
    .A(clknet_5_9__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_30_clk_p2c (.X(clknet_leaf_30_clk_p2c),
    .A(clknet_5_9__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_31_clk_p2c (.X(clknet_leaf_31_clk_p2c),
    .A(clknet_5_3__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_32_clk_p2c (.X(clknet_leaf_32_clk_p2c),
    .A(clknet_5_3__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_33_clk_p2c (.X(clknet_leaf_33_clk_p2c),
    .A(clknet_5_3__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_34_clk_p2c (.X(clknet_leaf_34_clk_p2c),
    .A(clknet_5_3__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_35_clk_p2c (.X(clknet_leaf_35_clk_p2c),
    .A(clknet_5_3__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_36_clk_p2c (.X(clknet_leaf_36_clk_p2c),
    .A(clknet_5_3__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_37_clk_p2c (.X(clknet_leaf_37_clk_p2c),
    .A(clknet_5_6__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_38_clk_p2c (.X(clknet_leaf_38_clk_p2c),
    .A(clknet_5_6__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_39_clk_p2c (.X(clknet_leaf_39_clk_p2c),
    .A(clknet_5_6__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_40_clk_p2c (.X(clknet_leaf_40_clk_p2c),
    .A(clknet_5_6__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_41_clk_p2c (.X(clknet_leaf_41_clk_p2c),
    .A(clknet_5_12__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_42_clk_p2c (.X(clknet_leaf_42_clk_p2c),
    .A(clknet_5_12__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_43_clk_p2c (.X(clknet_leaf_43_clk_p2c),
    .A(clknet_5_13__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_44_clk_p2c (.X(clknet_leaf_44_clk_p2c),
    .A(clknet_5_6__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_45_clk_p2c (.X(clknet_leaf_45_clk_p2c),
    .A(clknet_5_6__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_46_clk_p2c (.X(clknet_leaf_46_clk_p2c),
    .A(clknet_5_13__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_47_clk_p2c (.X(clknet_leaf_47_clk_p2c),
    .A(clknet_5_13__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_48_clk_p2c (.X(clknet_leaf_48_clk_p2c),
    .A(clknet_5_13__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_49_clk_p2c (.X(clknet_leaf_49_clk_p2c),
    .A(clknet_5_13__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_50_clk_p2c (.X(clknet_leaf_50_clk_p2c),
    .A(clknet_5_13__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_51_clk_p2c (.X(clknet_leaf_51_clk_p2c),
    .A(clknet_5_12__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_52_clk_p2c (.X(clknet_leaf_52_clk_p2c),
    .A(clknet_5_12__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_53_clk_p2c (.X(clknet_leaf_53_clk_p2c),
    .A(clknet_5_12__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_54_clk_p2c (.X(clknet_leaf_54_clk_p2c),
    .A(clknet_5_12__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_55_clk_p2c (.X(clknet_leaf_55_clk_p2c),
    .A(clknet_5_12__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_56_clk_p2c (.X(clknet_leaf_56_clk_p2c),
    .A(clknet_5_12__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_57_clk_p2c (.X(clknet_leaf_57_clk_p2c),
    .A(clknet_5_12__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_58_clk_p2c (.X(clknet_leaf_58_clk_p2c),
    .A(clknet_5_14__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_59_clk_p2c (.X(clknet_leaf_59_clk_p2c),
    .A(clknet_5_14__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_60_clk_p2c (.X(clknet_leaf_60_clk_p2c),
    .A(clknet_5_11__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_61_clk_p2c (.X(clknet_leaf_61_clk_p2c),
    .A(clknet_5_11__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_62_clk_p2c (.X(clknet_leaf_62_clk_p2c),
    .A(clknet_5_9__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_63_clk_p2c (.X(clknet_leaf_63_clk_p2c),
    .A(clknet_5_9__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_64_clk_p2c (.X(clknet_leaf_64_clk_p2c),
    .A(clknet_5_9__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_65_clk_p2c (.X(clknet_leaf_65_clk_p2c),
    .A(clknet_5_9__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_66_clk_p2c (.X(clknet_leaf_66_clk_p2c),
    .A(clknet_5_9__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_67_clk_p2c (.X(clknet_leaf_67_clk_p2c),
    .A(clknet_5_9__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_68_clk_p2c (.X(clknet_leaf_68_clk_p2c),
    .A(clknet_5_9__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_69_clk_p2c (.X(clknet_leaf_69_clk_p2c),
    .A(clknet_5_8__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_70_clk_p2c (.X(clknet_leaf_70_clk_p2c),
    .A(clknet_5_8__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_71_clk_p2c (.X(clknet_leaf_71_clk_p2c),
    .A(clknet_5_8__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_72_clk_p2c (.X(clknet_leaf_72_clk_p2c),
    .A(clknet_5_8__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_73_clk_p2c (.X(clknet_leaf_73_clk_p2c),
    .A(clknet_5_8__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_74_clk_p2c (.X(clknet_leaf_74_clk_p2c),
    .A(clknet_5_8__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_75_clk_p2c (.X(clknet_leaf_75_clk_p2c),
    .A(clknet_5_10__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_76_clk_p2c (.X(clknet_leaf_76_clk_p2c),
    .A(clknet_5_10__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_77_clk_p2c (.X(clknet_leaf_77_clk_p2c),
    .A(clknet_5_10__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_78_clk_p2c (.X(clknet_leaf_78_clk_p2c),
    .A(clknet_5_11__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_79_clk_p2c (.X(clknet_leaf_79_clk_p2c),
    .A(clknet_5_11__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_80_clk_p2c (.X(clknet_leaf_80_clk_p2c),
    .A(clknet_5_11__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_81_clk_p2c (.X(clknet_leaf_81_clk_p2c),
    .A(clknet_5_11__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_82_clk_p2c (.X(clknet_leaf_82_clk_p2c),
    .A(clknet_5_11__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_83_clk_p2c (.X(clknet_leaf_83_clk_p2c),
    .A(clknet_5_10__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_84_clk_p2c (.X(clknet_leaf_84_clk_p2c),
    .A(clknet_5_10__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_85_clk_p2c (.X(clknet_leaf_85_clk_p2c),
    .A(clknet_5_10__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_86_clk_p2c (.X(clknet_leaf_86_clk_p2c),
    .A(clknet_5_10__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_87_clk_p2c (.X(clknet_leaf_87_clk_p2c),
    .A(clknet_5_10__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_88_clk_p2c (.X(clknet_leaf_88_clk_p2c),
    .A(clknet_5_14__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_89_clk_p2c (.X(clknet_leaf_89_clk_p2c),
    .A(clknet_5_11__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_90_clk_p2c (.X(clknet_leaf_90_clk_p2c),
    .A(clknet_5_14__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_91_clk_p2c (.X(clknet_leaf_91_clk_p2c),
    .A(clknet_5_14__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_92_clk_p2c (.X(clknet_leaf_92_clk_p2c),
    .A(clknet_5_14__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_93_clk_p2c (.X(clknet_leaf_93_clk_p2c),
    .A(clknet_5_14__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_94_clk_p2c (.X(clknet_leaf_94_clk_p2c),
    .A(clknet_5_15__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_95_clk_p2c (.X(clknet_leaf_95_clk_p2c),
    .A(clknet_5_14__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_96_clk_p2c (.X(clknet_leaf_96_clk_p2c),
    .A(clknet_5_14__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_97_clk_p2c (.X(clknet_leaf_97_clk_p2c),
    .A(clknet_5_15__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_98_clk_p2c (.X(clknet_leaf_98_clk_p2c),
    .A(clknet_5_15__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_99_clk_p2c (.X(clknet_leaf_99_clk_p2c),
    .A(clknet_5_15__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_100_clk_p2c (.X(clknet_leaf_100_clk_p2c),
    .A(clknet_5_26__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_101_clk_p2c (.X(clknet_leaf_101_clk_p2c),
    .A(clknet_5_26__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_102_clk_p2c (.X(clknet_leaf_102_clk_p2c),
    .A(clknet_5_26__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_103_clk_p2c (.X(clknet_leaf_103_clk_p2c),
    .A(clknet_5_26__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_104_clk_p2c (.X(clknet_leaf_104_clk_p2c),
    .A(clknet_5_15__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_105_clk_p2c (.X(clknet_leaf_105_clk_p2c),
    .A(clknet_5_26__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_106_clk_p2c (.X(clknet_leaf_106_clk_p2c),
    .A(clknet_5_26__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_107_clk_p2c (.X(clknet_leaf_107_clk_p2c),
    .A(clknet_5_24__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_108_clk_p2c (.X(clknet_leaf_108_clk_p2c),
    .A(clknet_5_15__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_109_clk_p2c (.X(clknet_leaf_109_clk_p2c),
    .A(clknet_5_15__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_110_clk_p2c (.X(clknet_leaf_110_clk_p2c),
    .A(clknet_5_15__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_111_clk_p2c (.X(clknet_leaf_111_clk_p2c),
    .A(clknet_5_15__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_112_clk_p2c (.X(clknet_leaf_112_clk_p2c),
    .A(clknet_5_14__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_113_clk_p2c (.X(clknet_leaf_113_clk_p2c),
    .A(clknet_5_14__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_114_clk_p2c (.X(clknet_leaf_114_clk_p2c),
    .A(clknet_5_15__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_115_clk_p2c (.X(clknet_leaf_115_clk_p2c),
    .A(clknet_5_12__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_116_clk_p2c (.X(clknet_leaf_116_clk_p2c),
    .A(clknet_5_13__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_117_clk_p2c (.X(clknet_leaf_117_clk_p2c),
    .A(clknet_5_13__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_118_clk_p2c (.X(clknet_leaf_118_clk_p2c),
    .A(clknet_5_24__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_119_clk_p2c (.X(clknet_leaf_119_clk_p2c),
    .A(clknet_5_24__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_120_clk_p2c (.X(clknet_leaf_120_clk_p2c),
    .A(clknet_5_24__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_121_clk_p2c (.X(clknet_leaf_121_clk_p2c),
    .A(clknet_5_24__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_122_clk_p2c (.X(clknet_leaf_122_clk_p2c),
    .A(clknet_5_24__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_123_clk_p2c (.X(clknet_leaf_123_clk_p2c),
    .A(clknet_5_24__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_124_clk_p2c (.X(clknet_leaf_124_clk_p2c),
    .A(clknet_5_18__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_125_clk_p2c (.X(clknet_leaf_125_clk_p2c),
    .A(clknet_5_18__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_126_clk_p2c (.X(clknet_leaf_126_clk_p2c),
    .A(clknet_5_24__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_127_clk_p2c (.X(clknet_leaf_127_clk_p2c),
    .A(clknet_5_25__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_128_clk_p2c (.X(clknet_leaf_128_clk_p2c),
    .A(clknet_5_25__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_129_clk_p2c (.X(clknet_leaf_129_clk_p2c),
    .A(clknet_5_24__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_130_clk_p2c (.X(clknet_leaf_130_clk_p2c),
    .A(clknet_5_24__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_131_clk_p2c (.X(clknet_leaf_131_clk_p2c),
    .A(clknet_5_25__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_132_clk_p2c (.X(clknet_leaf_132_clk_p2c),
    .A(clknet_5_25__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_133_clk_p2c (.X(clknet_leaf_133_clk_p2c),
    .A(clknet_5_25__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_134_clk_p2c (.X(clknet_leaf_134_clk_p2c),
    .A(clknet_5_25__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_135_clk_p2c (.X(clknet_leaf_135_clk_p2c),
    .A(clknet_5_28__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_136_clk_p2c (.X(clknet_leaf_136_clk_p2c),
    .A(clknet_5_28__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_137_clk_p2c (.X(clknet_leaf_137_clk_p2c),
    .A(clknet_5_25__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_138_clk_p2c (.X(clknet_leaf_138_clk_p2c),
    .A(clknet_5_28__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_139_clk_p2c (.X(clknet_leaf_139_clk_p2c),
    .A(clknet_5_27__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_140_clk_p2c (.X(clknet_leaf_140_clk_p2c),
    .A(clknet_5_25__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_141_clk_p2c (.X(clknet_leaf_141_clk_p2c),
    .A(clknet_5_25__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_142_clk_p2c (.X(clknet_leaf_142_clk_p2c),
    .A(clknet_5_26__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_143_clk_p2c (.X(clknet_leaf_143_clk_p2c),
    .A(clknet_5_27__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_144_clk_p2c (.X(clknet_leaf_144_clk_p2c),
    .A(clknet_5_27__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_145_clk_p2c (.X(clknet_leaf_145_clk_p2c),
    .A(clknet_5_27__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_146_clk_p2c (.X(clknet_leaf_146_clk_p2c),
    .A(clknet_5_27__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_147_clk_p2c (.X(clknet_leaf_147_clk_p2c),
    .A(clknet_5_26__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_148_clk_p2c (.X(clknet_leaf_148_clk_p2c),
    .A(clknet_5_27__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_149_clk_p2c (.X(clknet_leaf_149_clk_p2c),
    .A(clknet_5_27__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_150_clk_p2c (.X(clknet_leaf_150_clk_p2c),
    .A(clknet_5_27__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_151_clk_p2c (.X(clknet_leaf_151_clk_p2c),
    .A(clknet_5_30__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_152_clk_p2c (.X(clknet_leaf_152_clk_p2c),
    .A(clknet_5_30__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_153_clk_p2c (.X(clknet_leaf_153_clk_p2c),
    .A(clknet_5_30__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_154_clk_p2c (.X(clknet_leaf_154_clk_p2c),
    .A(clknet_5_30__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_155_clk_p2c (.X(clknet_leaf_155_clk_p2c),
    .A(clknet_5_30__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_156_clk_p2c (.X(clknet_leaf_156_clk_p2c),
    .A(clknet_5_30__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_157_clk_p2c (.X(clknet_leaf_157_clk_p2c),
    .A(clknet_5_30__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_158_clk_p2c (.X(clknet_leaf_158_clk_p2c),
    .A(clknet_5_30__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_159_clk_p2c (.X(clknet_leaf_159_clk_p2c),
    .A(clknet_5_28__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_160_clk_p2c (.X(clknet_leaf_160_clk_p2c),
    .A(clknet_5_28__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_161_clk_p2c (.X(clknet_leaf_161_clk_p2c),
    .A(clknet_5_31__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_162_clk_p2c (.X(clknet_leaf_162_clk_p2c),
    .A(clknet_5_31__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_163_clk_p2c (.X(clknet_leaf_163_clk_p2c),
    .A(clknet_5_31__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_164_clk_p2c (.X(clknet_leaf_164_clk_p2c),
    .A(clknet_5_30__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_165_clk_p2c (.X(clknet_leaf_165_clk_p2c),
    .A(clknet_5_31__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_166_clk_p2c (.X(clknet_leaf_166_clk_p2c),
    .A(clknet_5_30__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_167_clk_p2c (.X(clknet_leaf_167_clk_p2c),
    .A(clknet_5_31__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_168_clk_p2c (.X(clknet_leaf_168_clk_p2c),
    .A(clknet_5_31__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_169_clk_p2c (.X(clknet_leaf_169_clk_p2c),
    .A(clknet_5_31__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_170_clk_p2c (.X(clknet_leaf_170_clk_p2c),
    .A(clknet_5_29__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_171_clk_p2c (.X(clknet_leaf_171_clk_p2c),
    .A(clknet_5_29__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_172_clk_p2c (.X(clknet_leaf_172_clk_p2c),
    .A(clknet_5_31__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_173_clk_p2c (.X(clknet_leaf_173_clk_p2c),
    .A(clknet_5_29__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_174_clk_p2c (.X(clknet_leaf_174_clk_p2c),
    .A(clknet_5_23__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_175_clk_p2c (.X(clknet_leaf_175_clk_p2c),
    .A(clknet_5_23__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_176_clk_p2c (.X(clknet_leaf_176_clk_p2c),
    .A(clknet_5_23__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_177_clk_p2c (.X(clknet_leaf_177_clk_p2c),
    .A(clknet_5_23__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_178_clk_p2c (.X(clknet_leaf_178_clk_p2c),
    .A(clknet_5_22__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_179_clk_p2c (.X(clknet_leaf_179_clk_p2c),
    .A(clknet_5_22__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_180_clk_p2c (.X(clknet_leaf_180_clk_p2c),
    .A(clknet_5_22__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_181_clk_p2c (.X(clknet_leaf_181_clk_p2c),
    .A(clknet_5_29__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_182_clk_p2c (.X(clknet_leaf_182_clk_p2c),
    .A(clknet_5_29__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_183_clk_p2c (.X(clknet_leaf_183_clk_p2c),
    .A(clknet_5_28__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_184_clk_p2c (.X(clknet_leaf_184_clk_p2c),
    .A(clknet_5_28__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_185_clk_p2c (.X(clknet_leaf_185_clk_p2c),
    .A(clknet_5_19__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_186_clk_p2c (.X(clknet_leaf_186_clk_p2c),
    .A(clknet_5_22__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_187_clk_p2c (.X(clknet_leaf_187_clk_p2c),
    .A(clknet_5_22__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_188_clk_p2c (.X(clknet_leaf_188_clk_p2c),
    .A(clknet_5_19__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_189_clk_p2c (.X(clknet_leaf_189_clk_p2c),
    .A(clknet_5_19__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_190_clk_p2c (.X(clknet_leaf_190_clk_p2c),
    .A(clknet_5_25__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_191_clk_p2c (.X(clknet_leaf_191_clk_p2c),
    .A(clknet_5_19__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_192_clk_p2c (.X(clknet_leaf_192_clk_p2c),
    .A(clknet_5_18__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_193_clk_p2c (.X(clknet_leaf_193_clk_p2c),
    .A(clknet_5_18__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_194_clk_p2c (.X(clknet_leaf_194_clk_p2c),
    .A(clknet_5_18__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_195_clk_p2c (.X(clknet_leaf_195_clk_p2c),
    .A(clknet_5_19__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_196_clk_p2c (.X(clknet_leaf_196_clk_p2c),
    .A(clknet_5_19__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_197_clk_p2c (.X(clknet_leaf_197_clk_p2c),
    .A(clknet_5_19__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_198_clk_p2c (.X(clknet_leaf_198_clk_p2c),
    .A(clknet_5_22__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_199_clk_p2c (.X(clknet_leaf_199_clk_p2c),
    .A(clknet_5_20__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_200_clk_p2c (.X(clknet_leaf_200_clk_p2c),
    .A(clknet_5_19__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_201_clk_p2c (.X(clknet_leaf_201_clk_p2c),
    .A(clknet_5_17__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_202_clk_p2c (.X(clknet_leaf_202_clk_p2c),
    .A(clknet_5_17__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_203_clk_p2c (.X(clknet_leaf_203_clk_p2c),
    .A(clknet_5_17__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_204_clk_p2c (.X(clknet_leaf_204_clk_p2c),
    .A(clknet_5_17__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_205_clk_p2c (.X(clknet_leaf_205_clk_p2c),
    .A(clknet_5_20__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_206_clk_p2c (.X(clknet_leaf_206_clk_p2c),
    .A(clknet_5_20__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_207_clk_p2c (.X(clknet_leaf_207_clk_p2c),
    .A(clknet_5_21__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_208_clk_p2c (.X(clknet_leaf_208_clk_p2c),
    .A(clknet_5_21__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_209_clk_p2c (.X(clknet_leaf_209_clk_p2c),
    .A(clknet_5_21__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_210_clk_p2c (.X(clknet_leaf_210_clk_p2c),
    .A(clknet_5_20__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_211_clk_p2c (.X(clknet_leaf_211_clk_p2c),
    .A(clknet_5_22__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_212_clk_p2c (.X(clknet_leaf_212_clk_p2c),
    .A(clknet_5_23__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_213_clk_p2c (.X(clknet_leaf_213_clk_p2c),
    .A(clknet_5_21__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_214_clk_p2c (.X(clknet_leaf_214_clk_p2c),
    .A(clknet_5_23__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_215_clk_p2c (.X(clknet_leaf_215_clk_p2c),
    .A(clknet_5_21__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_216_clk_p2c (.X(clknet_leaf_216_clk_p2c),
    .A(clknet_5_21__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_217_clk_p2c (.X(clknet_leaf_217_clk_p2c),
    .A(clknet_5_21__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_218_clk_p2c (.X(clknet_leaf_218_clk_p2c),
    .A(clknet_5_20__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_219_clk_p2c (.X(clknet_leaf_219_clk_p2c),
    .A(clknet_5_20__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_220_clk_p2c (.X(clknet_leaf_220_clk_p2c),
    .A(clknet_5_20__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_221_clk_p2c (.X(clknet_leaf_221_clk_p2c),
    .A(clknet_5_17__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_222_clk_p2c (.X(clknet_leaf_222_clk_p2c),
    .A(clknet_5_17__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_223_clk_p2c (.X(clknet_leaf_223_clk_p2c),
    .A(clknet_5_17__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_224_clk_p2c (.X(clknet_leaf_224_clk_p2c),
    .A(clknet_5_16__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_225_clk_p2c (.X(clknet_leaf_225_clk_p2c),
    .A(clknet_5_5__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_226_clk_p2c (.X(clknet_leaf_226_clk_p2c),
    .A(clknet_5_5__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_227_clk_p2c (.X(clknet_leaf_227_clk_p2c),
    .A(clknet_5_5__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_228_clk_p2c (.X(clknet_leaf_228_clk_p2c),
    .A(clknet_5_16__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_229_clk_p2c (.X(clknet_leaf_229_clk_p2c),
    .A(clknet_5_16__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_230_clk_p2c (.X(clknet_leaf_230_clk_p2c),
    .A(clknet_5_16__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_231_clk_p2c (.X(clknet_leaf_231_clk_p2c),
    .A(clknet_5_16__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_232_clk_p2c (.X(clknet_leaf_232_clk_p2c),
    .A(clknet_5_17__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_233_clk_p2c (.X(clknet_leaf_233_clk_p2c),
    .A(clknet_5_17__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_234_clk_p2c (.X(clknet_leaf_234_clk_p2c),
    .A(clknet_5_17__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_235_clk_p2c (.X(clknet_leaf_235_clk_p2c),
    .A(clknet_5_17__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_236_clk_p2c (.X(clknet_leaf_236_clk_p2c),
    .A(clknet_5_16__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_237_clk_p2c (.X(clknet_leaf_237_clk_p2c),
    .A(clknet_5_16__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_238_clk_p2c (.X(clknet_leaf_238_clk_p2c),
    .A(clknet_5_16__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_239_clk_p2c (.X(clknet_leaf_239_clk_p2c),
    .A(clknet_5_7__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_240_clk_p2c (.X(clknet_leaf_240_clk_p2c),
    .A(clknet_5_7__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_241_clk_p2c (.X(clknet_leaf_241_clk_p2c),
    .A(clknet_5_18__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_242_clk_p2c (.X(clknet_leaf_242_clk_p2c),
    .A(clknet_5_18__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_243_clk_p2c (.X(clknet_leaf_243_clk_p2c),
    .A(clknet_5_18__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_244_clk_p2c (.X(clknet_leaf_244_clk_p2c),
    .A(clknet_5_7__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_245_clk_p2c (.X(clknet_leaf_245_clk_p2c),
    .A(clknet_5_18__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_246_clk_p2c (.X(clknet_leaf_246_clk_p2c),
    .A(clknet_5_7__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_247_clk_p2c (.X(clknet_leaf_247_clk_p2c),
    .A(clknet_5_7__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_248_clk_p2c (.X(clknet_leaf_248_clk_p2c),
    .A(clknet_5_7__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_249_clk_p2c (.X(clknet_leaf_249_clk_p2c),
    .A(clknet_5_7__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_250_clk_p2c (.X(clknet_leaf_250_clk_p2c),
    .A(clknet_5_7__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_251_clk_p2c (.X(clknet_leaf_251_clk_p2c),
    .A(clknet_5_7__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_252_clk_p2c (.X(clknet_leaf_252_clk_p2c),
    .A(clknet_5_7__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_253_clk_p2c (.X(clknet_leaf_253_clk_p2c),
    .A(clknet_5_6__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_254_clk_p2c (.X(clknet_leaf_254_clk_p2c),
    .A(clknet_5_6__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_255_clk_p2c (.X(clknet_leaf_255_clk_p2c),
    .A(clknet_5_6__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_256_clk_p2c (.X(clknet_leaf_256_clk_p2c),
    .A(clknet_5_6__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_257_clk_p2c (.X(clknet_leaf_257_clk_p2c),
    .A(clknet_5_6__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_258_clk_p2c (.X(clknet_leaf_258_clk_p2c),
    .A(clknet_5_4__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_259_clk_p2c (.X(clknet_leaf_259_clk_p2c),
    .A(clknet_5_4__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_260_clk_p2c (.X(clknet_leaf_260_clk_p2c),
    .A(clknet_5_4__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_261_clk_p2c (.X(clknet_leaf_261_clk_p2c),
    .A(clknet_5_4__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_262_clk_p2c (.X(clknet_leaf_262_clk_p2c),
    .A(clknet_5_4__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_263_clk_p2c (.X(clknet_leaf_263_clk_p2c),
    .A(clknet_5_5__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_264_clk_p2c (.X(clknet_leaf_264_clk_p2c),
    .A(clknet_5_5__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_265_clk_p2c (.X(clknet_leaf_265_clk_p2c),
    .A(clknet_5_5__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_266_clk_p2c (.X(clknet_leaf_266_clk_p2c),
    .A(clknet_5_5__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_267_clk_p2c (.X(clknet_leaf_267_clk_p2c),
    .A(clknet_5_5__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_268_clk_p2c (.X(clknet_leaf_268_clk_p2c),
    .A(clknet_5_5__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_269_clk_p2c (.X(clknet_leaf_269_clk_p2c),
    .A(clknet_5_4__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_270_clk_p2c (.X(clknet_leaf_270_clk_p2c),
    .A(clknet_5_4__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_271_clk_p2c (.X(clknet_leaf_271_clk_p2c),
    .A(clknet_5_4__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_272_clk_p2c (.X(clknet_leaf_272_clk_p2c),
    .A(clknet_5_4__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_273_clk_p2c (.X(clknet_leaf_273_clk_p2c),
    .A(clknet_5_4__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_274_clk_p2c (.X(clknet_leaf_274_clk_p2c),
    .A(clknet_5_1__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_275_clk_p2c (.X(clknet_leaf_275_clk_p2c),
    .A(clknet_5_1__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_276_clk_p2c (.X(clknet_leaf_276_clk_p2c),
    .A(clknet_5_1__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_277_clk_p2c (.X(clknet_leaf_277_clk_p2c),
    .A(clknet_5_4__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_278_clk_p2c (.X(clknet_leaf_278_clk_p2c),
    .A(clknet_5_4__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_279_clk_p2c (.X(clknet_leaf_279_clk_p2c),
    .A(clknet_5_1__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_280_clk_p2c (.X(clknet_leaf_280_clk_p2c),
    .A(clknet_5_1__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_281_clk_p2c (.X(clknet_leaf_281_clk_p2c),
    .A(clknet_5_1__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_282_clk_p2c (.X(clknet_leaf_282_clk_p2c),
    .A(clknet_5_1__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_283_clk_p2c (.X(clknet_leaf_283_clk_p2c),
    .A(clknet_5_1__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_284_clk_p2c (.X(clknet_leaf_284_clk_p2c),
    .A(clknet_5_1__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_285_clk_p2c (.X(clknet_leaf_285_clk_p2c),
    .A(clknet_5_1__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_286_clk_p2c (.X(clknet_leaf_286_clk_p2c),
    .A(clknet_5_1__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_287_clk_p2c (.X(clknet_leaf_287_clk_p2c),
    .A(clknet_5_1__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_288_clk_p2c (.X(clknet_leaf_288_clk_p2c),
    .A(clknet_5_1__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_289_clk_p2c (.X(clknet_leaf_289_clk_p2c),
    .A(clknet_5_1__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_290_clk_p2c (.X(clknet_leaf_290_clk_p2c),
    .A(clknet_5_0__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_291_clk_p2c (.X(clknet_leaf_291_clk_p2c),
    .A(clknet_5_0__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_292_clk_p2c (.X(clknet_leaf_292_clk_p2c),
    .A(clknet_5_0__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_293_clk_p2c (.X(clknet_leaf_293_clk_p2c),
    .A(clknet_5_0__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_294_clk_p2c (.X(clknet_leaf_294_clk_p2c),
    .A(clknet_5_0__leaf_clk_p2c));
 sg13g2_buf_2 clkbuf_0_clk_p2c (.A(clk_p2c),
    .X(clknet_0_clk_p2c));
 sg13g2_buf_4 clkbuf_4_0_0_clk_p2c (.X(clknet_4_0_0_clk_p2c),
    .A(clknet_0_clk_p2c));
 sg13g2_buf_4 clkbuf_4_1_0_clk_p2c (.X(clknet_4_1_0_clk_p2c),
    .A(clknet_0_clk_p2c));
 sg13g2_buf_4 clkbuf_4_2_0_clk_p2c (.X(clknet_4_2_0_clk_p2c),
    .A(clknet_0_clk_p2c));
 sg13g2_buf_4 clkbuf_4_3_0_clk_p2c (.X(clknet_4_3_0_clk_p2c),
    .A(clknet_0_clk_p2c));
 sg13g2_buf_4 clkbuf_4_4_0_clk_p2c (.X(clknet_4_4_0_clk_p2c),
    .A(clknet_0_clk_p2c));
 sg13g2_buf_4 clkbuf_4_5_0_clk_p2c (.X(clknet_4_5_0_clk_p2c),
    .A(clknet_0_clk_p2c));
 sg13g2_buf_4 clkbuf_4_6_0_clk_p2c (.X(clknet_4_6_0_clk_p2c),
    .A(clknet_0_clk_p2c));
 sg13g2_buf_4 clkbuf_4_7_0_clk_p2c (.X(clknet_4_7_0_clk_p2c),
    .A(clknet_0_clk_p2c));
 sg13g2_buf_4 clkbuf_4_8_0_clk_p2c (.X(clknet_4_8_0_clk_p2c),
    .A(clknet_0_clk_p2c));
 sg13g2_buf_4 clkbuf_4_9_0_clk_p2c (.X(clknet_4_9_0_clk_p2c),
    .A(clknet_0_clk_p2c));
 sg13g2_buf_4 clkbuf_4_10_0_clk_p2c (.X(clknet_4_10_0_clk_p2c),
    .A(clknet_0_clk_p2c));
 sg13g2_buf_4 clkbuf_4_11_0_clk_p2c (.X(clknet_4_11_0_clk_p2c),
    .A(clknet_0_clk_p2c));
 sg13g2_buf_4 clkbuf_4_12_0_clk_p2c (.X(clknet_4_12_0_clk_p2c),
    .A(clknet_0_clk_p2c));
 sg13g2_buf_4 clkbuf_4_13_0_clk_p2c (.X(clknet_4_13_0_clk_p2c),
    .A(clknet_0_clk_p2c));
 sg13g2_buf_4 clkbuf_4_14_0_clk_p2c (.X(clknet_4_14_0_clk_p2c),
    .A(clknet_0_clk_p2c));
 sg13g2_buf_4 clkbuf_4_15_0_clk_p2c (.X(clknet_4_15_0_clk_p2c),
    .A(clknet_0_clk_p2c));
 sg13g2_buf_2 clkbuf_5_0__f_clk_p2c (.A(clknet_4_0_0_clk_p2c),
    .X(clknet_5_0__leaf_clk_p2c));
 sg13g2_buf_2 clkbuf_5_1__f_clk_p2c (.A(clknet_4_0_0_clk_p2c),
    .X(clknet_5_1__leaf_clk_p2c));
 sg13g2_buf_2 clkbuf_5_2__f_clk_p2c (.A(clknet_4_1_0_clk_p2c),
    .X(clknet_5_2__leaf_clk_p2c));
 sg13g2_buf_2 clkbuf_5_3__f_clk_p2c (.A(clknet_4_1_0_clk_p2c),
    .X(clknet_5_3__leaf_clk_p2c));
 sg13g2_buf_2 clkbuf_5_4__f_clk_p2c (.A(clknet_4_2_0_clk_p2c),
    .X(clknet_5_4__leaf_clk_p2c));
 sg13g2_buf_2 clkbuf_5_5__f_clk_p2c (.A(clknet_4_2_0_clk_p2c),
    .X(clknet_5_5__leaf_clk_p2c));
 sg13g2_buf_2 clkbuf_5_6__f_clk_p2c (.A(clknet_4_3_0_clk_p2c),
    .X(clknet_5_6__leaf_clk_p2c));
 sg13g2_buf_2 clkbuf_5_7__f_clk_p2c (.A(clknet_4_3_0_clk_p2c),
    .X(clknet_5_7__leaf_clk_p2c));
 sg13g2_buf_2 clkbuf_5_8__f_clk_p2c (.A(clknet_4_4_0_clk_p2c),
    .X(clknet_5_8__leaf_clk_p2c));
 sg13g2_buf_2 clkbuf_5_9__f_clk_p2c (.A(clknet_4_4_0_clk_p2c),
    .X(clknet_5_9__leaf_clk_p2c));
 sg13g2_buf_2 clkbuf_5_10__f_clk_p2c (.A(clknet_4_5_0_clk_p2c),
    .X(clknet_5_10__leaf_clk_p2c));
 sg13g2_buf_2 clkbuf_5_11__f_clk_p2c (.A(clknet_4_5_0_clk_p2c),
    .X(clknet_5_11__leaf_clk_p2c));
 sg13g2_buf_2 clkbuf_5_12__f_clk_p2c (.A(clknet_4_6_0_clk_p2c),
    .X(clknet_5_12__leaf_clk_p2c));
 sg13g2_buf_2 clkbuf_5_13__f_clk_p2c (.A(clknet_4_6_0_clk_p2c),
    .X(clknet_5_13__leaf_clk_p2c));
 sg13g2_buf_2 clkbuf_5_14__f_clk_p2c (.A(clknet_4_7_0_clk_p2c),
    .X(clknet_5_14__leaf_clk_p2c));
 sg13g2_buf_2 clkbuf_5_15__f_clk_p2c (.A(clknet_4_7_0_clk_p2c),
    .X(clknet_5_15__leaf_clk_p2c));
 sg13g2_buf_2 clkbuf_5_16__f_clk_p2c (.A(clknet_4_8_0_clk_p2c),
    .X(clknet_5_16__leaf_clk_p2c));
 sg13g2_buf_2 clkbuf_5_17__f_clk_p2c (.A(clknet_4_8_0_clk_p2c),
    .X(clknet_5_17__leaf_clk_p2c));
 sg13g2_buf_2 clkbuf_5_18__f_clk_p2c (.A(clknet_4_9_0_clk_p2c),
    .X(clknet_5_18__leaf_clk_p2c));
 sg13g2_buf_2 clkbuf_5_19__f_clk_p2c (.A(clknet_4_9_0_clk_p2c),
    .X(clknet_5_19__leaf_clk_p2c));
 sg13g2_buf_2 clkbuf_5_20__f_clk_p2c (.A(clknet_4_10_0_clk_p2c),
    .X(clknet_5_20__leaf_clk_p2c));
 sg13g2_buf_2 clkbuf_5_21__f_clk_p2c (.A(clknet_4_10_0_clk_p2c),
    .X(clknet_5_21__leaf_clk_p2c));
 sg13g2_buf_2 clkbuf_5_22__f_clk_p2c (.A(clknet_4_11_0_clk_p2c),
    .X(clknet_5_22__leaf_clk_p2c));
 sg13g2_buf_2 clkbuf_5_23__f_clk_p2c (.A(clknet_4_11_0_clk_p2c),
    .X(clknet_5_23__leaf_clk_p2c));
 sg13g2_buf_2 clkbuf_5_24__f_clk_p2c (.A(clknet_4_12_0_clk_p2c),
    .X(clknet_5_24__leaf_clk_p2c));
 sg13g2_buf_2 clkbuf_5_25__f_clk_p2c (.A(clknet_4_12_0_clk_p2c),
    .X(clknet_5_25__leaf_clk_p2c));
 sg13g2_buf_2 clkbuf_5_26__f_clk_p2c (.A(clknet_4_13_0_clk_p2c),
    .X(clknet_5_26__leaf_clk_p2c));
 sg13g2_buf_2 clkbuf_5_27__f_clk_p2c (.A(clknet_4_13_0_clk_p2c),
    .X(clknet_5_27__leaf_clk_p2c));
 sg13g2_buf_2 clkbuf_5_28__f_clk_p2c (.A(clknet_4_14_0_clk_p2c),
    .X(clknet_5_28__leaf_clk_p2c));
 sg13g2_buf_2 clkbuf_5_29__f_clk_p2c (.A(clknet_4_14_0_clk_p2c),
    .X(clknet_5_29__leaf_clk_p2c));
 sg13g2_buf_2 clkbuf_5_30__f_clk_p2c (.A(clknet_4_15_0_clk_p2c),
    .X(clknet_5_30__leaf_clk_p2c));
 sg13g2_buf_2 clkbuf_5_31__f_clk_p2c (.A(clknet_4_15_0_clk_p2c),
    .X(clknet_5_31__leaf_clk_p2c));
 sg13g2_fill_8 FILLER_0_0_0 ();
 sg13g2_fill_8 FILLER_0_0_8 ();
 sg13g2_fill_8 FILLER_0_0_16 ();
 sg13g2_fill_8 FILLER_0_0_24 ();
 sg13g2_fill_8 FILLER_0_0_32 ();
 sg13g2_fill_8 FILLER_0_0_40 ();
 sg13g2_fill_8 FILLER_0_0_48 ();
 sg13g2_fill_8 FILLER_0_0_56 ();
 sg13g2_fill_8 FILLER_0_0_64 ();
 sg13g2_fill_8 FILLER_0_0_72 ();
 sg13g2_fill_8 FILLER_0_0_80 ();
 sg13g2_fill_8 FILLER_0_0_88 ();
 sg13g2_fill_8 FILLER_0_0_96 ();
 sg13g2_fill_8 FILLER_0_0_104 ();
 sg13g2_fill_8 FILLER_0_0_112 ();
 sg13g2_fill_8 FILLER_0_0_120 ();
 sg13g2_fill_8 FILLER_0_0_128 ();
 sg13g2_fill_8 FILLER_0_0_136 ();
 sg13g2_fill_8 FILLER_0_0_144 ();
 sg13g2_fill_8 FILLER_0_0_152 ();
 sg13g2_fill_8 FILLER_0_0_160 ();
 sg13g2_fill_8 FILLER_0_0_168 ();
 sg13g2_fill_8 FILLER_0_0_176 ();
 sg13g2_fill_8 FILLER_0_0_184 ();
 sg13g2_fill_8 FILLER_0_0_192 ();
 sg13g2_fill_8 FILLER_0_0_200 ();
 sg13g2_fill_8 FILLER_0_0_208 ();
 sg13g2_fill_8 FILLER_0_0_216 ();
 sg13g2_fill_8 FILLER_0_0_224 ();
 sg13g2_fill_8 FILLER_0_0_232 ();
 sg13g2_fill_8 FILLER_0_0_240 ();
 sg13g2_fill_8 FILLER_0_0_248 ();
 sg13g2_fill_8 FILLER_0_0_256 ();
 sg13g2_fill_8 FILLER_0_0_264 ();
 sg13g2_fill_8 FILLER_0_0_272 ();
 sg13g2_fill_8 FILLER_0_0_280 ();
 sg13g2_fill_8 FILLER_0_0_288 ();
 sg13g2_fill_8 FILLER_0_0_296 ();
 sg13g2_fill_8 FILLER_0_0_304 ();
 sg13g2_fill_8 FILLER_0_0_312 ();
 sg13g2_fill_8 FILLER_0_0_320 ();
 sg13g2_fill_8 FILLER_0_0_328 ();
 sg13g2_fill_8 FILLER_0_0_336 ();
 sg13g2_fill_8 FILLER_0_0_344 ();
 sg13g2_fill_8 FILLER_0_0_352 ();
 sg13g2_fill_8 FILLER_0_0_360 ();
 sg13g2_fill_8 FILLER_0_0_368 ();
 sg13g2_fill_8 FILLER_0_0_376 ();
 sg13g2_fill_8 FILLER_0_0_384 ();
 sg13g2_fill_8 FILLER_0_0_392 ();
 sg13g2_fill_8 FILLER_0_0_400 ();
 sg13g2_fill_8 FILLER_0_0_408 ();
 sg13g2_fill_8 FILLER_0_0_416 ();
 sg13g2_fill_8 FILLER_0_0_424 ();
 sg13g2_fill_8 FILLER_0_0_432 ();
 sg13g2_fill_8 FILLER_0_0_440 ();
 sg13g2_fill_8 FILLER_0_0_448 ();
 sg13g2_fill_8 FILLER_0_0_456 ();
 sg13g2_fill_8 FILLER_0_0_464 ();
 sg13g2_fill_8 FILLER_0_0_472 ();
 sg13g2_fill_8 FILLER_0_0_480 ();
 sg13g2_fill_8 FILLER_0_0_488 ();
 sg13g2_fill_8 FILLER_0_0_496 ();
 sg13g2_fill_8 FILLER_0_0_504 ();
 sg13g2_fill_8 FILLER_0_0_512 ();
 sg13g2_fill_8 FILLER_0_0_520 ();
 sg13g2_fill_8 FILLER_0_0_528 ();
 sg13g2_fill_8 FILLER_0_0_536 ();
 sg13g2_fill_8 FILLER_0_0_544 ();
 sg13g2_fill_8 FILLER_0_0_552 ();
 sg13g2_fill_8 FILLER_0_0_560 ();
 sg13g2_fill_8 FILLER_0_0_568 ();
 sg13g2_fill_8 FILLER_0_0_576 ();
 sg13g2_fill_8 FILLER_0_0_584 ();
 sg13g2_fill_8 FILLER_0_0_592 ();
 sg13g2_fill_8 FILLER_0_0_600 ();
 sg13g2_fill_8 FILLER_0_0_608 ();
 sg13g2_fill_8 FILLER_0_0_616 ();
 sg13g2_fill_8 FILLER_0_0_624 ();
 sg13g2_fill_8 FILLER_0_0_632 ();
 sg13g2_fill_8 FILLER_0_0_640 ();
 sg13g2_fill_8 FILLER_0_0_648 ();
 sg13g2_fill_8 FILLER_0_0_656 ();
 sg13g2_fill_8 FILLER_0_0_664 ();
 sg13g2_fill_8 FILLER_0_0_672 ();
 sg13g2_fill_8 FILLER_0_0_680 ();
 sg13g2_fill_8 FILLER_0_0_688 ();
 sg13g2_fill_8 FILLER_0_0_696 ();
 sg13g2_fill_8 FILLER_0_0_704 ();
 sg13g2_fill_8 FILLER_0_0_712 ();
 sg13g2_fill_8 FILLER_0_0_720 ();
 sg13g2_fill_8 FILLER_0_0_728 ();
 sg13g2_fill_8 FILLER_0_0_736 ();
 sg13g2_fill_8 FILLER_0_0_744 ();
 sg13g2_fill_8 FILLER_0_0_752 ();
 sg13g2_fill_8 FILLER_0_0_760 ();
 sg13g2_fill_8 FILLER_0_0_768 ();
 sg13g2_fill_8 FILLER_0_0_776 ();
 sg13g2_fill_8 FILLER_0_0_784 ();
 sg13g2_fill_8 FILLER_0_0_792 ();
 sg13g2_fill_8 FILLER_0_0_800 ();
 sg13g2_fill_8 FILLER_0_0_808 ();
 sg13g2_fill_8 FILLER_0_0_816 ();
 sg13g2_fill_8 FILLER_0_0_824 ();
 sg13g2_fill_8 FILLER_0_0_832 ();
 sg13g2_fill_8 FILLER_0_0_840 ();
 sg13g2_fill_8 FILLER_0_0_848 ();
 sg13g2_fill_8 FILLER_0_0_856 ();
 sg13g2_fill_8 FILLER_0_0_864 ();
 sg13g2_fill_8 FILLER_0_0_872 ();
 sg13g2_fill_8 FILLER_0_0_880 ();
 sg13g2_fill_8 FILLER_0_0_888 ();
 sg13g2_fill_8 FILLER_0_0_896 ();
 sg13g2_fill_8 FILLER_0_0_904 ();
 sg13g2_fill_8 FILLER_0_0_912 ();
 sg13g2_fill_8 FILLER_0_0_920 ();
 sg13g2_fill_8 FILLER_0_0_928 ();
 sg13g2_fill_8 FILLER_0_0_936 ();
 sg13g2_fill_8 FILLER_0_0_944 ();
 sg13g2_fill_8 FILLER_0_0_952 ();
 sg13g2_fill_8 FILLER_0_0_960 ();
 sg13g2_fill_8 FILLER_0_0_968 ();
 sg13g2_fill_8 FILLER_0_0_976 ();
 sg13g2_fill_8 FILLER_0_0_984 ();
 sg13g2_fill_8 FILLER_0_0_992 ();
 sg13g2_fill_8 FILLER_0_0_1000 ();
 sg13g2_fill_8 FILLER_0_0_1008 ();
 sg13g2_fill_8 FILLER_0_0_1016 ();
 sg13g2_fill_8 FILLER_0_0_1024 ();
 sg13g2_fill_8 FILLER_0_0_1032 ();
 sg13g2_fill_8 FILLER_0_0_1040 ();
 sg13g2_fill_8 FILLER_0_0_1048 ();
 sg13g2_fill_8 FILLER_0_0_1056 ();
 sg13g2_fill_8 FILLER_0_0_1064 ();
 sg13g2_fill_8 FILLER_0_0_1072 ();
 sg13g2_fill_8 FILLER_0_0_1080 ();
 sg13g2_fill_8 FILLER_0_0_1088 ();
 sg13g2_fill_8 FILLER_0_0_1096 ();
 sg13g2_fill_8 FILLER_0_0_1104 ();
 sg13g2_fill_8 FILLER_0_0_1112 ();
 sg13g2_fill_8 FILLER_0_0_1120 ();
 sg13g2_fill_8 FILLER_0_0_1128 ();
 sg13g2_fill_8 FILLER_0_0_1136 ();
 sg13g2_fill_8 FILLER_0_0_1144 ();
 sg13g2_fill_8 FILLER_0_0_1152 ();
 sg13g2_fill_8 FILLER_0_0_1160 ();
 sg13g2_fill_8 FILLER_0_0_1168 ();
 sg13g2_fill_8 FILLER_0_0_1176 ();
 sg13g2_fill_8 FILLER_0_0_1184 ();
 sg13g2_fill_8 FILLER_0_0_1192 ();
 sg13g2_fill_8 FILLER_0_0_1200 ();
 sg13g2_fill_8 FILLER_0_0_1208 ();
 sg13g2_fill_8 FILLER_0_0_1216 ();
 sg13g2_fill_4 FILLER_0_0_1224 ();
 sg13g2_fill_8 FILLER_0_1_0 ();
 sg13g2_fill_8 FILLER_0_1_8 ();
 sg13g2_fill_8 FILLER_0_1_16 ();
 sg13g2_fill_8 FILLER_0_1_24 ();
 sg13g2_fill_8 FILLER_0_1_32 ();
 sg13g2_fill_8 FILLER_0_1_40 ();
 sg13g2_fill_8 FILLER_0_1_48 ();
 sg13g2_fill_8 FILLER_0_1_56 ();
 sg13g2_fill_8 FILLER_0_1_64 ();
 sg13g2_fill_8 FILLER_0_1_72 ();
 sg13g2_fill_8 FILLER_0_1_80 ();
 sg13g2_fill_8 FILLER_0_1_88 ();
 sg13g2_fill_8 FILLER_0_1_96 ();
 sg13g2_fill_8 FILLER_0_1_104 ();
 sg13g2_fill_8 FILLER_0_1_112 ();
 sg13g2_fill_8 FILLER_0_1_120 ();
 sg13g2_fill_8 FILLER_0_1_128 ();
 sg13g2_fill_8 FILLER_0_1_136 ();
 sg13g2_fill_8 FILLER_0_1_144 ();
 sg13g2_fill_8 FILLER_0_1_152 ();
 sg13g2_fill_8 FILLER_0_1_160 ();
 sg13g2_fill_8 FILLER_0_1_168 ();
 sg13g2_fill_8 FILLER_0_1_176 ();
 sg13g2_fill_8 FILLER_0_1_184 ();
 sg13g2_fill_8 FILLER_0_1_192 ();
 sg13g2_fill_8 FILLER_0_1_200 ();
 sg13g2_fill_8 FILLER_0_1_208 ();
 sg13g2_fill_8 FILLER_0_1_216 ();
 sg13g2_fill_8 FILLER_0_1_224 ();
 sg13g2_fill_8 FILLER_0_1_232 ();
 sg13g2_fill_8 FILLER_0_1_240 ();
 sg13g2_fill_8 FILLER_0_1_248 ();
 sg13g2_fill_8 FILLER_0_1_256 ();
 sg13g2_fill_8 FILLER_0_1_264 ();
 sg13g2_fill_8 FILLER_0_1_272 ();
 sg13g2_fill_8 FILLER_0_1_280 ();
 sg13g2_fill_8 FILLER_0_1_288 ();
 sg13g2_fill_8 FILLER_0_1_296 ();
 sg13g2_fill_8 FILLER_0_1_304 ();
 sg13g2_fill_8 FILLER_0_1_312 ();
 sg13g2_fill_8 FILLER_0_1_320 ();
 sg13g2_fill_8 FILLER_0_1_328 ();
 sg13g2_fill_8 FILLER_0_1_336 ();
 sg13g2_fill_8 FILLER_0_1_344 ();
 sg13g2_fill_8 FILLER_0_1_352 ();
 sg13g2_fill_8 FILLER_0_1_360 ();
 sg13g2_fill_8 FILLER_0_1_368 ();
 sg13g2_fill_8 FILLER_0_1_376 ();
 sg13g2_fill_8 FILLER_0_1_384 ();
 sg13g2_fill_8 FILLER_0_1_392 ();
 sg13g2_fill_8 FILLER_0_1_400 ();
 sg13g2_fill_8 FILLER_0_1_408 ();
 sg13g2_fill_8 FILLER_0_1_416 ();
 sg13g2_fill_8 FILLER_0_1_424 ();
 sg13g2_fill_8 FILLER_0_1_432 ();
 sg13g2_fill_8 FILLER_0_1_440 ();
 sg13g2_fill_8 FILLER_0_1_448 ();
 sg13g2_fill_8 FILLER_0_1_456 ();
 sg13g2_fill_8 FILLER_0_1_464 ();
 sg13g2_fill_8 FILLER_0_1_472 ();
 sg13g2_fill_8 FILLER_0_1_480 ();
 sg13g2_fill_8 FILLER_0_1_488 ();
 sg13g2_fill_8 FILLER_0_1_496 ();
 sg13g2_fill_8 FILLER_0_1_504 ();
 sg13g2_fill_8 FILLER_0_1_512 ();
 sg13g2_fill_8 FILLER_0_1_520 ();
 sg13g2_fill_8 FILLER_0_1_528 ();
 sg13g2_fill_8 FILLER_0_1_536 ();
 sg13g2_fill_8 FILLER_0_1_544 ();
 sg13g2_fill_8 FILLER_0_1_552 ();
 sg13g2_fill_8 FILLER_0_1_560 ();
 sg13g2_fill_8 FILLER_0_1_568 ();
 sg13g2_fill_8 FILLER_0_1_576 ();
 sg13g2_fill_8 FILLER_0_1_584 ();
 sg13g2_fill_8 FILLER_0_1_592 ();
 sg13g2_fill_8 FILLER_0_1_600 ();
 sg13g2_fill_8 FILLER_0_1_608 ();
 sg13g2_fill_8 FILLER_0_1_616 ();
 sg13g2_fill_8 FILLER_0_1_624 ();
 sg13g2_fill_8 FILLER_0_1_632 ();
 sg13g2_fill_8 FILLER_0_1_640 ();
 sg13g2_fill_8 FILLER_0_1_648 ();
 sg13g2_fill_8 FILLER_0_1_656 ();
 sg13g2_fill_8 FILLER_0_1_664 ();
 sg13g2_fill_8 FILLER_0_1_672 ();
 sg13g2_fill_8 FILLER_0_1_680 ();
 sg13g2_fill_8 FILLER_0_1_688 ();
 sg13g2_fill_8 FILLER_0_1_696 ();
 sg13g2_fill_8 FILLER_0_1_704 ();
 sg13g2_fill_8 FILLER_0_1_712 ();
 sg13g2_fill_8 FILLER_0_1_720 ();
 sg13g2_fill_8 FILLER_0_1_728 ();
 sg13g2_fill_8 FILLER_0_1_736 ();
 sg13g2_fill_8 FILLER_0_1_744 ();
 sg13g2_fill_8 FILLER_0_1_752 ();
 sg13g2_fill_8 FILLER_0_1_760 ();
 sg13g2_fill_8 FILLER_0_1_768 ();
 sg13g2_fill_8 FILLER_0_1_776 ();
 sg13g2_fill_8 FILLER_0_1_784 ();
 sg13g2_fill_8 FILLER_0_1_792 ();
 sg13g2_fill_8 FILLER_0_1_800 ();
 sg13g2_fill_8 FILLER_0_1_808 ();
 sg13g2_fill_8 FILLER_0_1_816 ();
 sg13g2_fill_8 FILLER_0_1_824 ();
 sg13g2_fill_8 FILLER_0_1_832 ();
 sg13g2_fill_8 FILLER_0_1_840 ();
 sg13g2_fill_8 FILLER_0_1_848 ();
 sg13g2_fill_8 FILLER_0_1_856 ();
 sg13g2_fill_8 FILLER_0_1_864 ();
 sg13g2_fill_8 FILLER_0_1_872 ();
 sg13g2_fill_8 FILLER_0_1_880 ();
 sg13g2_fill_8 FILLER_0_1_888 ();
 sg13g2_fill_8 FILLER_0_1_896 ();
 sg13g2_fill_8 FILLER_0_1_904 ();
 sg13g2_fill_8 FILLER_0_1_912 ();
 sg13g2_fill_8 FILLER_0_1_920 ();
 sg13g2_fill_8 FILLER_0_1_928 ();
 sg13g2_fill_8 FILLER_0_1_936 ();
 sg13g2_fill_8 FILLER_0_1_944 ();
 sg13g2_fill_8 FILLER_0_1_952 ();
 sg13g2_fill_8 FILLER_0_1_960 ();
 sg13g2_fill_8 FILLER_0_1_968 ();
 sg13g2_fill_8 FILLER_0_1_976 ();
 sg13g2_fill_8 FILLER_0_1_984 ();
 sg13g2_fill_8 FILLER_0_1_992 ();
 sg13g2_fill_8 FILLER_0_1_1000 ();
 sg13g2_fill_8 FILLER_0_1_1008 ();
 sg13g2_fill_8 FILLER_0_1_1016 ();
 sg13g2_fill_8 FILLER_0_1_1024 ();
 sg13g2_fill_8 FILLER_0_1_1032 ();
 sg13g2_fill_8 FILLER_0_1_1040 ();
 sg13g2_fill_8 FILLER_0_1_1048 ();
 sg13g2_fill_8 FILLER_0_1_1056 ();
 sg13g2_fill_8 FILLER_0_1_1064 ();
 sg13g2_fill_8 FILLER_0_1_1072 ();
 sg13g2_fill_8 FILLER_0_1_1080 ();
 sg13g2_fill_8 FILLER_0_1_1088 ();
 sg13g2_fill_8 FILLER_0_1_1096 ();
 sg13g2_fill_8 FILLER_0_1_1104 ();
 sg13g2_fill_8 FILLER_0_1_1112 ();
 sg13g2_fill_8 FILLER_0_1_1120 ();
 sg13g2_fill_8 FILLER_0_1_1128 ();
 sg13g2_fill_8 FILLER_0_1_1136 ();
 sg13g2_fill_8 FILLER_0_1_1144 ();
 sg13g2_fill_8 FILLER_0_1_1152 ();
 sg13g2_fill_8 FILLER_0_1_1160 ();
 sg13g2_fill_8 FILLER_0_1_1168 ();
 sg13g2_fill_8 FILLER_0_1_1176 ();
 sg13g2_fill_8 FILLER_0_1_1184 ();
 sg13g2_fill_8 FILLER_0_1_1192 ();
 sg13g2_fill_8 FILLER_0_1_1200 ();
 sg13g2_fill_8 FILLER_0_1_1208 ();
 sg13g2_fill_8 FILLER_0_1_1216 ();
 sg13g2_fill_4 FILLER_0_1_1224 ();
 sg13g2_fill_8 FILLER_0_2_0 ();
 sg13g2_fill_8 FILLER_0_2_8 ();
 sg13g2_fill_8 FILLER_0_2_16 ();
 sg13g2_fill_8 FILLER_0_2_24 ();
 sg13g2_fill_8 FILLER_0_2_32 ();
 sg13g2_fill_8 FILLER_0_2_40 ();
 sg13g2_fill_8 FILLER_0_2_48 ();
 sg13g2_fill_8 FILLER_0_2_56 ();
 sg13g2_fill_8 FILLER_0_2_64 ();
 sg13g2_fill_8 FILLER_0_2_72 ();
 sg13g2_fill_8 FILLER_0_2_80 ();
 sg13g2_fill_8 FILLER_0_2_88 ();
 sg13g2_fill_8 FILLER_0_2_96 ();
 sg13g2_fill_8 FILLER_0_2_104 ();
 sg13g2_fill_8 FILLER_0_2_112 ();
 sg13g2_fill_8 FILLER_0_2_120 ();
 sg13g2_fill_8 FILLER_0_2_128 ();
 sg13g2_fill_8 FILLER_0_2_136 ();
 sg13g2_fill_8 FILLER_0_2_144 ();
 sg13g2_fill_8 FILLER_0_2_152 ();
 sg13g2_fill_8 FILLER_0_2_160 ();
 sg13g2_fill_8 FILLER_0_2_168 ();
 sg13g2_fill_8 FILLER_0_2_176 ();
 sg13g2_fill_8 FILLER_0_2_184 ();
 sg13g2_fill_8 FILLER_0_2_192 ();
 sg13g2_fill_8 FILLER_0_2_200 ();
 sg13g2_fill_8 FILLER_0_2_208 ();
 sg13g2_fill_8 FILLER_0_2_216 ();
 sg13g2_fill_8 FILLER_0_2_224 ();
 sg13g2_fill_8 FILLER_0_2_232 ();
 sg13g2_fill_8 FILLER_0_2_240 ();
 sg13g2_fill_8 FILLER_0_2_248 ();
 sg13g2_fill_8 FILLER_0_2_256 ();
 sg13g2_fill_8 FILLER_0_2_264 ();
 sg13g2_fill_8 FILLER_0_2_272 ();
 sg13g2_fill_8 FILLER_0_2_280 ();
 sg13g2_fill_8 FILLER_0_2_288 ();
 sg13g2_fill_8 FILLER_0_2_296 ();
 sg13g2_fill_8 FILLER_0_2_304 ();
 sg13g2_fill_8 FILLER_0_2_312 ();
 sg13g2_fill_8 FILLER_0_2_320 ();
 sg13g2_fill_8 FILLER_0_2_328 ();
 sg13g2_fill_8 FILLER_0_2_336 ();
 sg13g2_fill_8 FILLER_0_2_344 ();
 sg13g2_fill_8 FILLER_0_2_352 ();
 sg13g2_fill_8 FILLER_0_2_360 ();
 sg13g2_fill_8 FILLER_0_2_368 ();
 sg13g2_fill_8 FILLER_0_2_376 ();
 sg13g2_fill_8 FILLER_0_2_384 ();
 sg13g2_fill_8 FILLER_0_2_392 ();
 sg13g2_fill_8 FILLER_0_2_400 ();
 sg13g2_fill_8 FILLER_0_2_408 ();
 sg13g2_fill_8 FILLER_0_2_416 ();
 sg13g2_fill_8 FILLER_0_2_424 ();
 sg13g2_fill_8 FILLER_0_2_432 ();
 sg13g2_fill_8 FILLER_0_2_440 ();
 sg13g2_fill_8 FILLER_0_2_448 ();
 sg13g2_fill_8 FILLER_0_2_456 ();
 sg13g2_fill_8 FILLER_0_2_464 ();
 sg13g2_fill_8 FILLER_0_2_472 ();
 sg13g2_fill_8 FILLER_0_2_480 ();
 sg13g2_fill_8 FILLER_0_2_488 ();
 sg13g2_fill_8 FILLER_0_2_496 ();
 sg13g2_fill_8 FILLER_0_2_504 ();
 sg13g2_fill_8 FILLER_0_2_512 ();
 sg13g2_fill_8 FILLER_0_2_520 ();
 sg13g2_fill_8 FILLER_0_2_528 ();
 sg13g2_fill_8 FILLER_0_2_536 ();
 sg13g2_fill_8 FILLER_0_2_544 ();
 sg13g2_fill_8 FILLER_0_2_552 ();
 sg13g2_fill_8 FILLER_0_2_560 ();
 sg13g2_fill_8 FILLER_0_2_568 ();
 sg13g2_fill_8 FILLER_0_2_576 ();
 sg13g2_fill_8 FILLER_0_2_584 ();
 sg13g2_fill_8 FILLER_0_2_592 ();
 sg13g2_fill_8 FILLER_0_2_600 ();
 sg13g2_fill_8 FILLER_0_2_608 ();
 sg13g2_fill_8 FILLER_0_2_616 ();
 sg13g2_fill_8 FILLER_0_2_624 ();
 sg13g2_fill_8 FILLER_0_2_632 ();
 sg13g2_fill_8 FILLER_0_2_640 ();
 sg13g2_fill_8 FILLER_0_2_648 ();
 sg13g2_fill_8 FILLER_0_2_656 ();
 sg13g2_fill_8 FILLER_0_2_664 ();
 sg13g2_fill_8 FILLER_0_2_672 ();
 sg13g2_fill_8 FILLER_0_2_680 ();
 sg13g2_fill_8 FILLER_0_2_688 ();
 sg13g2_fill_8 FILLER_0_2_696 ();
 sg13g2_fill_8 FILLER_0_2_704 ();
 sg13g2_fill_8 FILLER_0_2_712 ();
 sg13g2_fill_8 FILLER_0_2_720 ();
 sg13g2_fill_8 FILLER_0_2_728 ();
 sg13g2_fill_8 FILLER_0_2_736 ();
 sg13g2_fill_8 FILLER_0_2_744 ();
 sg13g2_fill_8 FILLER_0_2_752 ();
 sg13g2_fill_8 FILLER_0_2_760 ();
 sg13g2_fill_8 FILLER_0_2_768 ();
 sg13g2_fill_8 FILLER_0_2_776 ();
 sg13g2_fill_8 FILLER_0_2_784 ();
 sg13g2_fill_8 FILLER_0_2_792 ();
 sg13g2_fill_8 FILLER_0_2_800 ();
 sg13g2_fill_8 FILLER_0_2_808 ();
 sg13g2_fill_8 FILLER_0_2_816 ();
 sg13g2_fill_8 FILLER_0_2_824 ();
 sg13g2_fill_8 FILLER_0_2_832 ();
 sg13g2_fill_8 FILLER_0_2_840 ();
 sg13g2_fill_8 FILLER_0_2_848 ();
 sg13g2_fill_8 FILLER_0_2_856 ();
 sg13g2_fill_8 FILLER_0_2_864 ();
 sg13g2_fill_8 FILLER_0_2_872 ();
 sg13g2_fill_8 FILLER_0_2_880 ();
 sg13g2_fill_8 FILLER_0_2_888 ();
 sg13g2_fill_8 FILLER_0_2_896 ();
 sg13g2_fill_8 FILLER_0_2_904 ();
 sg13g2_fill_8 FILLER_0_2_912 ();
 sg13g2_fill_8 FILLER_0_2_920 ();
 sg13g2_fill_8 FILLER_0_2_928 ();
 sg13g2_fill_8 FILLER_0_2_936 ();
 sg13g2_fill_8 FILLER_0_2_944 ();
 sg13g2_fill_8 FILLER_0_2_952 ();
 sg13g2_fill_8 FILLER_0_2_960 ();
 sg13g2_fill_8 FILLER_0_2_968 ();
 sg13g2_fill_8 FILLER_0_2_976 ();
 sg13g2_fill_8 FILLER_0_2_984 ();
 sg13g2_fill_8 FILLER_0_2_992 ();
 sg13g2_fill_8 FILLER_0_2_1000 ();
 sg13g2_fill_8 FILLER_0_2_1008 ();
 sg13g2_fill_8 FILLER_0_2_1016 ();
 sg13g2_fill_8 FILLER_0_2_1024 ();
 sg13g2_fill_8 FILLER_0_2_1032 ();
 sg13g2_fill_8 FILLER_0_2_1040 ();
 sg13g2_fill_8 FILLER_0_2_1048 ();
 sg13g2_fill_8 FILLER_0_2_1056 ();
 sg13g2_fill_8 FILLER_0_2_1064 ();
 sg13g2_fill_8 FILLER_0_2_1072 ();
 sg13g2_fill_8 FILLER_0_2_1080 ();
 sg13g2_fill_8 FILLER_0_2_1088 ();
 sg13g2_fill_8 FILLER_0_2_1096 ();
 sg13g2_fill_8 FILLER_0_2_1104 ();
 sg13g2_fill_8 FILLER_0_2_1112 ();
 sg13g2_fill_8 FILLER_0_2_1120 ();
 sg13g2_fill_8 FILLER_0_2_1128 ();
 sg13g2_fill_8 FILLER_0_2_1136 ();
 sg13g2_fill_8 FILLER_0_2_1144 ();
 sg13g2_fill_8 FILLER_0_2_1152 ();
 sg13g2_fill_8 FILLER_0_2_1160 ();
 sg13g2_fill_8 FILLER_0_2_1168 ();
 sg13g2_fill_8 FILLER_0_2_1176 ();
 sg13g2_fill_8 FILLER_0_2_1184 ();
 sg13g2_fill_8 FILLER_0_2_1192 ();
 sg13g2_fill_8 FILLER_0_2_1200 ();
 sg13g2_fill_8 FILLER_0_2_1208 ();
 sg13g2_fill_8 FILLER_0_2_1216 ();
 sg13g2_fill_4 FILLER_0_2_1224 ();
 sg13g2_fill_8 FILLER_0_3_0 ();
 sg13g2_fill_8 FILLER_0_3_8 ();
 sg13g2_fill_8 FILLER_0_3_16 ();
 sg13g2_fill_8 FILLER_0_3_24 ();
 sg13g2_fill_8 FILLER_0_3_32 ();
 sg13g2_fill_8 FILLER_0_3_40 ();
 sg13g2_fill_8 FILLER_0_3_48 ();
 sg13g2_fill_8 FILLER_0_3_56 ();
 sg13g2_fill_8 FILLER_0_3_64 ();
 sg13g2_fill_8 FILLER_0_3_72 ();
 sg13g2_fill_8 FILLER_0_3_80 ();
 sg13g2_fill_8 FILLER_0_3_88 ();
 sg13g2_fill_8 FILLER_0_3_96 ();
 sg13g2_fill_8 FILLER_0_3_104 ();
 sg13g2_fill_8 FILLER_0_3_112 ();
 sg13g2_fill_8 FILLER_0_3_120 ();
 sg13g2_fill_8 FILLER_0_3_128 ();
 sg13g2_fill_8 FILLER_0_3_136 ();
 sg13g2_fill_8 FILLER_0_3_144 ();
 sg13g2_fill_8 FILLER_0_3_152 ();
 sg13g2_fill_8 FILLER_0_3_160 ();
 sg13g2_fill_8 FILLER_0_3_168 ();
 sg13g2_fill_8 FILLER_0_3_176 ();
 sg13g2_fill_8 FILLER_0_3_184 ();
 sg13g2_fill_8 FILLER_0_3_192 ();
 sg13g2_fill_8 FILLER_0_3_200 ();
 sg13g2_fill_8 FILLER_0_3_208 ();
 sg13g2_fill_8 FILLER_0_3_216 ();
 sg13g2_fill_8 FILLER_0_3_224 ();
 sg13g2_fill_8 FILLER_0_3_232 ();
 sg13g2_fill_8 FILLER_0_3_240 ();
 sg13g2_fill_8 FILLER_0_3_248 ();
 sg13g2_fill_8 FILLER_0_3_256 ();
 sg13g2_fill_8 FILLER_0_3_264 ();
 sg13g2_fill_8 FILLER_0_3_272 ();
 sg13g2_fill_8 FILLER_0_3_280 ();
 sg13g2_fill_8 FILLER_0_3_288 ();
 sg13g2_fill_8 FILLER_0_3_296 ();
 sg13g2_fill_8 FILLER_0_3_304 ();
 sg13g2_fill_8 FILLER_0_3_312 ();
 sg13g2_fill_8 FILLER_0_3_320 ();
 sg13g2_fill_8 FILLER_0_3_328 ();
 sg13g2_fill_8 FILLER_0_3_336 ();
 sg13g2_fill_8 FILLER_0_3_344 ();
 sg13g2_fill_8 FILLER_0_3_352 ();
 sg13g2_fill_8 FILLER_0_3_360 ();
 sg13g2_fill_8 FILLER_0_3_368 ();
 sg13g2_fill_8 FILLER_0_3_376 ();
 sg13g2_fill_8 FILLER_0_3_384 ();
 sg13g2_fill_8 FILLER_0_3_392 ();
 sg13g2_fill_8 FILLER_0_3_400 ();
 sg13g2_fill_8 FILLER_0_3_408 ();
 sg13g2_fill_8 FILLER_0_3_416 ();
 sg13g2_fill_8 FILLER_0_3_424 ();
 sg13g2_fill_8 FILLER_0_3_432 ();
 sg13g2_fill_8 FILLER_0_3_440 ();
 sg13g2_fill_8 FILLER_0_3_448 ();
 sg13g2_fill_8 FILLER_0_3_456 ();
 sg13g2_fill_8 FILLER_0_3_464 ();
 sg13g2_fill_8 FILLER_0_3_472 ();
 sg13g2_fill_8 FILLER_0_3_480 ();
 sg13g2_fill_8 FILLER_0_3_488 ();
 sg13g2_fill_8 FILLER_0_3_496 ();
 sg13g2_fill_8 FILLER_0_3_504 ();
 sg13g2_fill_8 FILLER_0_3_512 ();
 sg13g2_fill_8 FILLER_0_3_520 ();
 sg13g2_fill_8 FILLER_0_3_528 ();
 sg13g2_fill_8 FILLER_0_3_536 ();
 sg13g2_fill_8 FILLER_0_3_544 ();
 sg13g2_fill_8 FILLER_0_3_552 ();
 sg13g2_fill_8 FILLER_0_3_560 ();
 sg13g2_fill_8 FILLER_0_3_568 ();
 sg13g2_fill_8 FILLER_0_3_576 ();
 sg13g2_fill_8 FILLER_0_3_584 ();
 sg13g2_fill_8 FILLER_0_3_592 ();
 sg13g2_fill_8 FILLER_0_3_600 ();
 sg13g2_fill_8 FILLER_0_3_608 ();
 sg13g2_fill_8 FILLER_0_3_616 ();
 sg13g2_fill_8 FILLER_0_3_624 ();
 sg13g2_fill_8 FILLER_0_3_632 ();
 sg13g2_fill_8 FILLER_0_3_640 ();
 sg13g2_fill_8 FILLER_0_3_648 ();
 sg13g2_fill_8 FILLER_0_3_656 ();
 sg13g2_fill_8 FILLER_0_3_664 ();
 sg13g2_fill_8 FILLER_0_3_672 ();
 sg13g2_fill_8 FILLER_0_3_680 ();
 sg13g2_fill_8 FILLER_0_3_688 ();
 sg13g2_fill_8 FILLER_0_3_696 ();
 sg13g2_fill_8 FILLER_0_3_704 ();
 sg13g2_fill_8 FILLER_0_3_712 ();
 sg13g2_fill_8 FILLER_0_3_720 ();
 sg13g2_fill_8 FILLER_0_3_728 ();
 sg13g2_fill_8 FILLER_0_3_736 ();
 sg13g2_fill_8 FILLER_0_3_744 ();
 sg13g2_fill_8 FILLER_0_3_752 ();
 sg13g2_fill_8 FILLER_0_3_760 ();
 sg13g2_fill_8 FILLER_0_3_768 ();
 sg13g2_fill_8 FILLER_0_3_776 ();
 sg13g2_fill_8 FILLER_0_3_784 ();
 sg13g2_fill_8 FILLER_0_3_792 ();
 sg13g2_fill_8 FILLER_0_3_800 ();
 sg13g2_fill_8 FILLER_0_3_808 ();
 sg13g2_fill_8 FILLER_0_3_816 ();
 sg13g2_fill_8 FILLER_0_3_824 ();
 sg13g2_fill_8 FILLER_0_3_832 ();
 sg13g2_fill_8 FILLER_0_3_840 ();
 sg13g2_fill_8 FILLER_0_3_848 ();
 sg13g2_fill_8 FILLER_0_3_856 ();
 sg13g2_fill_8 FILLER_0_3_864 ();
 sg13g2_fill_8 FILLER_0_3_872 ();
 sg13g2_fill_8 FILLER_0_3_880 ();
 sg13g2_fill_8 FILLER_0_3_888 ();
 sg13g2_fill_8 FILLER_0_3_896 ();
 sg13g2_fill_8 FILLER_0_3_904 ();
 sg13g2_fill_8 FILLER_0_3_912 ();
 sg13g2_fill_8 FILLER_0_3_920 ();
 sg13g2_fill_8 FILLER_0_3_928 ();
 sg13g2_fill_8 FILLER_0_3_936 ();
 sg13g2_fill_8 FILLER_0_3_944 ();
 sg13g2_fill_8 FILLER_0_3_952 ();
 sg13g2_fill_8 FILLER_0_3_960 ();
 sg13g2_fill_8 FILLER_0_3_968 ();
 sg13g2_fill_8 FILLER_0_3_976 ();
 sg13g2_fill_8 FILLER_0_3_984 ();
 sg13g2_fill_8 FILLER_0_3_992 ();
 sg13g2_fill_8 FILLER_0_3_1000 ();
 sg13g2_fill_8 FILLER_0_3_1008 ();
 sg13g2_fill_8 FILLER_0_3_1016 ();
 sg13g2_fill_8 FILLER_0_3_1024 ();
 sg13g2_fill_8 FILLER_0_3_1032 ();
 sg13g2_fill_8 FILLER_0_3_1040 ();
 sg13g2_fill_8 FILLER_0_3_1048 ();
 sg13g2_fill_8 FILLER_0_3_1056 ();
 sg13g2_fill_8 FILLER_0_3_1064 ();
 sg13g2_fill_8 FILLER_0_3_1072 ();
 sg13g2_fill_8 FILLER_0_3_1080 ();
 sg13g2_fill_8 FILLER_0_3_1088 ();
 sg13g2_fill_8 FILLER_0_3_1096 ();
 sg13g2_fill_8 FILLER_0_3_1104 ();
 sg13g2_fill_8 FILLER_0_3_1112 ();
 sg13g2_fill_8 FILLER_0_3_1120 ();
 sg13g2_fill_8 FILLER_0_3_1128 ();
 sg13g2_fill_8 FILLER_0_3_1136 ();
 sg13g2_fill_8 FILLER_0_3_1144 ();
 sg13g2_fill_8 FILLER_0_3_1152 ();
 sg13g2_fill_8 FILLER_0_3_1160 ();
 sg13g2_fill_8 FILLER_0_3_1168 ();
 sg13g2_fill_8 FILLER_0_3_1176 ();
 sg13g2_fill_8 FILLER_0_3_1184 ();
 sg13g2_fill_8 FILLER_0_3_1192 ();
 sg13g2_fill_8 FILLER_0_3_1200 ();
 sg13g2_fill_8 FILLER_0_3_1208 ();
 sg13g2_fill_8 FILLER_0_3_1216 ();
 sg13g2_fill_4 FILLER_0_3_1224 ();
 sg13g2_fill_8 FILLER_0_4_0 ();
 sg13g2_fill_8 FILLER_0_4_8 ();
 sg13g2_fill_8 FILLER_0_4_16 ();
 sg13g2_fill_8 FILLER_0_4_24 ();
 sg13g2_fill_8 FILLER_0_4_32 ();
 sg13g2_fill_8 FILLER_0_4_40 ();
 sg13g2_fill_8 FILLER_0_4_48 ();
 sg13g2_fill_8 FILLER_0_4_56 ();
 sg13g2_fill_8 FILLER_0_4_64 ();
 sg13g2_fill_8 FILLER_0_4_72 ();
 sg13g2_fill_8 FILLER_0_4_80 ();
 sg13g2_fill_8 FILLER_0_4_88 ();
 sg13g2_fill_8 FILLER_0_4_96 ();
 sg13g2_fill_8 FILLER_0_4_104 ();
 sg13g2_fill_8 FILLER_0_4_112 ();
 sg13g2_fill_8 FILLER_0_4_120 ();
 sg13g2_fill_8 FILLER_0_4_128 ();
 sg13g2_fill_8 FILLER_0_4_136 ();
 sg13g2_fill_8 FILLER_0_4_144 ();
 sg13g2_fill_8 FILLER_0_4_152 ();
 sg13g2_fill_8 FILLER_0_4_160 ();
 sg13g2_fill_8 FILLER_0_4_168 ();
 sg13g2_fill_8 FILLER_0_4_176 ();
 sg13g2_fill_8 FILLER_0_4_184 ();
 sg13g2_fill_8 FILLER_0_4_192 ();
 sg13g2_fill_8 FILLER_0_4_200 ();
 sg13g2_fill_8 FILLER_0_4_208 ();
 sg13g2_fill_8 FILLER_0_4_216 ();
 sg13g2_fill_8 FILLER_0_4_224 ();
 sg13g2_fill_8 FILLER_0_4_232 ();
 sg13g2_fill_8 FILLER_0_4_240 ();
 sg13g2_fill_8 FILLER_0_4_248 ();
 sg13g2_fill_8 FILLER_0_4_256 ();
 sg13g2_fill_8 FILLER_0_4_264 ();
 sg13g2_fill_8 FILLER_0_4_272 ();
 sg13g2_fill_8 FILLER_0_4_280 ();
 sg13g2_fill_8 FILLER_0_4_288 ();
 sg13g2_fill_8 FILLER_0_4_296 ();
 sg13g2_fill_8 FILLER_0_4_304 ();
 sg13g2_fill_8 FILLER_0_4_312 ();
 sg13g2_fill_8 FILLER_0_4_320 ();
 sg13g2_fill_8 FILLER_0_4_328 ();
 sg13g2_fill_8 FILLER_0_4_336 ();
 sg13g2_fill_8 FILLER_0_4_344 ();
 sg13g2_fill_8 FILLER_0_4_352 ();
 sg13g2_fill_8 FILLER_0_4_360 ();
 sg13g2_fill_8 FILLER_0_4_368 ();
 sg13g2_fill_8 FILLER_0_4_376 ();
 sg13g2_fill_8 FILLER_0_4_384 ();
 sg13g2_fill_8 FILLER_0_4_392 ();
 sg13g2_fill_8 FILLER_0_4_400 ();
 sg13g2_fill_8 FILLER_0_4_408 ();
 sg13g2_fill_8 FILLER_0_4_416 ();
 sg13g2_fill_8 FILLER_0_4_424 ();
 sg13g2_fill_8 FILLER_0_4_432 ();
 sg13g2_fill_8 FILLER_0_4_440 ();
 sg13g2_fill_8 FILLER_0_4_448 ();
 sg13g2_fill_8 FILLER_0_4_456 ();
 sg13g2_fill_8 FILLER_0_4_464 ();
 sg13g2_fill_8 FILLER_0_4_472 ();
 sg13g2_fill_8 FILLER_0_4_480 ();
 sg13g2_fill_8 FILLER_0_4_488 ();
 sg13g2_fill_8 FILLER_0_4_496 ();
 sg13g2_fill_8 FILLER_0_4_504 ();
 sg13g2_fill_8 FILLER_0_4_512 ();
 sg13g2_fill_8 FILLER_0_4_520 ();
 sg13g2_fill_8 FILLER_0_4_528 ();
 sg13g2_fill_8 FILLER_0_4_536 ();
 sg13g2_fill_8 FILLER_0_4_544 ();
 sg13g2_fill_8 FILLER_0_4_552 ();
 sg13g2_fill_8 FILLER_0_4_560 ();
 sg13g2_fill_8 FILLER_0_4_568 ();
 sg13g2_fill_8 FILLER_0_4_576 ();
 sg13g2_fill_8 FILLER_0_4_584 ();
 sg13g2_fill_8 FILLER_0_4_592 ();
 sg13g2_fill_8 FILLER_0_4_600 ();
 sg13g2_fill_8 FILLER_0_4_608 ();
 sg13g2_fill_8 FILLER_0_4_616 ();
 sg13g2_fill_8 FILLER_0_4_624 ();
 sg13g2_fill_8 FILLER_0_4_632 ();
 sg13g2_fill_8 FILLER_0_4_640 ();
 sg13g2_fill_8 FILLER_0_4_648 ();
 sg13g2_fill_8 FILLER_0_4_656 ();
 sg13g2_fill_8 FILLER_0_4_664 ();
 sg13g2_fill_8 FILLER_0_4_672 ();
 sg13g2_fill_8 FILLER_0_4_680 ();
 sg13g2_fill_8 FILLER_0_4_688 ();
 sg13g2_fill_8 FILLER_0_4_696 ();
 sg13g2_fill_8 FILLER_0_4_704 ();
 sg13g2_fill_8 FILLER_0_4_712 ();
 sg13g2_fill_8 FILLER_0_4_720 ();
 sg13g2_fill_8 FILLER_0_4_728 ();
 sg13g2_fill_8 FILLER_0_4_736 ();
 sg13g2_fill_8 FILLER_0_4_744 ();
 sg13g2_fill_8 FILLER_0_4_752 ();
 sg13g2_fill_8 FILLER_0_4_760 ();
 sg13g2_fill_8 FILLER_0_4_768 ();
 sg13g2_fill_8 FILLER_0_4_776 ();
 sg13g2_fill_8 FILLER_0_4_784 ();
 sg13g2_fill_8 FILLER_0_4_792 ();
 sg13g2_fill_8 FILLER_0_4_800 ();
 sg13g2_fill_8 FILLER_0_4_808 ();
 sg13g2_fill_8 FILLER_0_4_816 ();
 sg13g2_fill_8 FILLER_0_4_824 ();
 sg13g2_fill_8 FILLER_0_4_832 ();
 sg13g2_fill_8 FILLER_0_4_840 ();
 sg13g2_fill_8 FILLER_0_4_848 ();
 sg13g2_fill_8 FILLER_0_4_856 ();
 sg13g2_fill_8 FILLER_0_4_864 ();
 sg13g2_fill_8 FILLER_0_4_872 ();
 sg13g2_fill_8 FILLER_0_4_880 ();
 sg13g2_fill_8 FILLER_0_4_888 ();
 sg13g2_fill_8 FILLER_0_4_896 ();
 sg13g2_fill_8 FILLER_0_4_904 ();
 sg13g2_fill_8 FILLER_0_4_912 ();
 sg13g2_fill_8 FILLER_0_4_920 ();
 sg13g2_fill_8 FILLER_0_4_928 ();
 sg13g2_fill_8 FILLER_0_4_936 ();
 sg13g2_fill_8 FILLER_0_4_944 ();
 sg13g2_fill_8 FILLER_0_4_952 ();
 sg13g2_fill_8 FILLER_0_4_960 ();
 sg13g2_fill_8 FILLER_0_4_968 ();
 sg13g2_fill_8 FILLER_0_4_976 ();
 sg13g2_fill_8 FILLER_0_4_984 ();
 sg13g2_fill_8 FILLER_0_4_992 ();
 sg13g2_fill_8 FILLER_0_4_1000 ();
 sg13g2_fill_8 FILLER_0_4_1008 ();
 sg13g2_fill_8 FILLER_0_4_1016 ();
 sg13g2_fill_8 FILLER_0_4_1024 ();
 sg13g2_fill_8 FILLER_0_4_1032 ();
 sg13g2_fill_8 FILLER_0_4_1040 ();
 sg13g2_fill_8 FILLER_0_4_1048 ();
 sg13g2_fill_8 FILLER_0_4_1056 ();
 sg13g2_fill_8 FILLER_0_4_1064 ();
 sg13g2_fill_8 FILLER_0_4_1072 ();
 sg13g2_fill_8 FILLER_0_4_1080 ();
 sg13g2_fill_8 FILLER_0_4_1088 ();
 sg13g2_fill_8 FILLER_0_4_1096 ();
 sg13g2_fill_8 FILLER_0_4_1104 ();
 sg13g2_fill_8 FILLER_0_4_1112 ();
 sg13g2_fill_8 FILLER_0_4_1120 ();
 sg13g2_fill_8 FILLER_0_4_1128 ();
 sg13g2_fill_8 FILLER_0_4_1136 ();
 sg13g2_fill_8 FILLER_0_4_1144 ();
 sg13g2_fill_8 FILLER_0_4_1152 ();
 sg13g2_fill_8 FILLER_0_4_1160 ();
 sg13g2_fill_8 FILLER_0_4_1168 ();
 sg13g2_fill_8 FILLER_0_4_1176 ();
 sg13g2_fill_8 FILLER_0_4_1184 ();
 sg13g2_fill_8 FILLER_0_4_1192 ();
 sg13g2_fill_8 FILLER_0_4_1200 ();
 sg13g2_fill_8 FILLER_0_4_1208 ();
 sg13g2_fill_8 FILLER_0_4_1216 ();
 sg13g2_fill_4 FILLER_0_4_1224 ();
 sg13g2_fill_8 FILLER_0_5_0 ();
 sg13g2_fill_8 FILLER_0_5_8 ();
 sg13g2_fill_8 FILLER_0_5_16 ();
 sg13g2_fill_8 FILLER_0_5_24 ();
 sg13g2_fill_8 FILLER_0_5_32 ();
 sg13g2_fill_8 FILLER_0_5_40 ();
 sg13g2_fill_8 FILLER_0_5_48 ();
 sg13g2_fill_8 FILLER_0_5_56 ();
 sg13g2_fill_8 FILLER_0_5_64 ();
 sg13g2_fill_8 FILLER_0_5_72 ();
 sg13g2_fill_8 FILLER_0_5_80 ();
 sg13g2_fill_8 FILLER_0_5_88 ();
 sg13g2_fill_8 FILLER_0_5_96 ();
 sg13g2_fill_8 FILLER_0_5_104 ();
 sg13g2_fill_8 FILLER_0_5_112 ();
 sg13g2_fill_8 FILLER_0_5_120 ();
 sg13g2_fill_8 FILLER_0_5_128 ();
 sg13g2_fill_8 FILLER_0_5_136 ();
 sg13g2_fill_8 FILLER_0_5_144 ();
 sg13g2_fill_8 FILLER_0_5_152 ();
 sg13g2_fill_8 FILLER_0_5_160 ();
 sg13g2_fill_8 FILLER_0_5_168 ();
 sg13g2_fill_8 FILLER_0_5_176 ();
 sg13g2_fill_8 FILLER_0_5_184 ();
 sg13g2_fill_8 FILLER_0_5_192 ();
 sg13g2_fill_8 FILLER_0_5_200 ();
 sg13g2_fill_8 FILLER_0_5_208 ();
 sg13g2_fill_8 FILLER_0_5_216 ();
 sg13g2_fill_8 FILLER_0_5_224 ();
 sg13g2_fill_8 FILLER_0_5_232 ();
 sg13g2_fill_8 FILLER_0_5_240 ();
 sg13g2_fill_8 FILLER_0_5_248 ();
 sg13g2_fill_8 FILLER_0_5_256 ();
 sg13g2_fill_8 FILLER_0_5_264 ();
 sg13g2_fill_8 FILLER_0_5_272 ();
 sg13g2_fill_8 FILLER_0_5_280 ();
 sg13g2_fill_8 FILLER_0_5_288 ();
 sg13g2_fill_8 FILLER_0_5_296 ();
 sg13g2_fill_8 FILLER_0_5_304 ();
 sg13g2_fill_8 FILLER_0_5_312 ();
 sg13g2_fill_8 FILLER_0_5_320 ();
 sg13g2_fill_8 FILLER_0_5_328 ();
 sg13g2_fill_8 FILLER_0_5_336 ();
 sg13g2_fill_8 FILLER_0_5_344 ();
 sg13g2_fill_8 FILLER_0_5_352 ();
 sg13g2_fill_8 FILLER_0_5_360 ();
 sg13g2_fill_8 FILLER_0_5_368 ();
 sg13g2_fill_8 FILLER_0_5_376 ();
 sg13g2_fill_8 FILLER_0_5_384 ();
 sg13g2_fill_8 FILLER_0_5_392 ();
 sg13g2_fill_8 FILLER_0_5_400 ();
 sg13g2_fill_8 FILLER_0_5_408 ();
 sg13g2_fill_8 FILLER_0_5_416 ();
 sg13g2_fill_8 FILLER_0_5_424 ();
 sg13g2_fill_8 FILLER_0_5_432 ();
 sg13g2_fill_8 FILLER_0_5_440 ();
 sg13g2_fill_8 FILLER_0_5_448 ();
 sg13g2_fill_8 FILLER_0_5_456 ();
 sg13g2_fill_8 FILLER_0_5_464 ();
 sg13g2_fill_8 FILLER_0_5_472 ();
 sg13g2_fill_8 FILLER_0_5_480 ();
 sg13g2_fill_8 FILLER_0_5_488 ();
 sg13g2_fill_8 FILLER_0_5_496 ();
 sg13g2_fill_8 FILLER_0_5_504 ();
 sg13g2_fill_8 FILLER_0_5_512 ();
 sg13g2_fill_8 FILLER_0_5_520 ();
 sg13g2_fill_8 FILLER_0_5_528 ();
 sg13g2_fill_8 FILLER_0_5_536 ();
 sg13g2_fill_8 FILLER_0_5_544 ();
 sg13g2_fill_8 FILLER_0_5_552 ();
 sg13g2_fill_8 FILLER_0_5_560 ();
 sg13g2_fill_8 FILLER_0_5_568 ();
 sg13g2_fill_8 FILLER_0_5_576 ();
 sg13g2_fill_8 FILLER_0_5_584 ();
 sg13g2_fill_8 FILLER_0_5_592 ();
 sg13g2_fill_8 FILLER_0_5_600 ();
 sg13g2_fill_8 FILLER_0_5_608 ();
 sg13g2_fill_8 FILLER_0_5_616 ();
 sg13g2_fill_8 FILLER_0_5_624 ();
 sg13g2_fill_8 FILLER_0_5_632 ();
 sg13g2_fill_8 FILLER_0_5_640 ();
 sg13g2_fill_8 FILLER_0_5_648 ();
 sg13g2_fill_8 FILLER_0_5_656 ();
 sg13g2_fill_8 FILLER_0_5_664 ();
 sg13g2_fill_8 FILLER_0_5_672 ();
 sg13g2_fill_8 FILLER_0_5_680 ();
 sg13g2_fill_8 FILLER_0_5_688 ();
 sg13g2_fill_8 FILLER_0_5_696 ();
 sg13g2_fill_8 FILLER_0_5_704 ();
 sg13g2_fill_8 FILLER_0_5_712 ();
 sg13g2_fill_8 FILLER_0_5_720 ();
 sg13g2_fill_8 FILLER_0_5_728 ();
 sg13g2_fill_8 FILLER_0_5_736 ();
 sg13g2_fill_8 FILLER_0_5_744 ();
 sg13g2_fill_8 FILLER_0_5_752 ();
 sg13g2_fill_8 FILLER_0_5_760 ();
 sg13g2_fill_8 FILLER_0_5_768 ();
 sg13g2_fill_8 FILLER_0_5_776 ();
 sg13g2_fill_8 FILLER_0_5_784 ();
 sg13g2_fill_8 FILLER_0_5_792 ();
 sg13g2_fill_8 FILLER_0_5_800 ();
 sg13g2_fill_8 FILLER_0_5_808 ();
 sg13g2_fill_8 FILLER_0_5_816 ();
 sg13g2_fill_8 FILLER_0_5_824 ();
 sg13g2_fill_8 FILLER_0_5_832 ();
 sg13g2_fill_8 FILLER_0_5_840 ();
 sg13g2_fill_8 FILLER_0_5_848 ();
 sg13g2_fill_8 FILLER_0_5_856 ();
 sg13g2_fill_8 FILLER_0_5_864 ();
 sg13g2_fill_8 FILLER_0_5_872 ();
 sg13g2_fill_8 FILLER_0_5_880 ();
 sg13g2_fill_8 FILLER_0_5_888 ();
 sg13g2_fill_8 FILLER_0_5_896 ();
 sg13g2_fill_8 FILLER_0_5_904 ();
 sg13g2_fill_8 FILLER_0_5_912 ();
 sg13g2_fill_8 FILLER_0_5_920 ();
 sg13g2_fill_8 FILLER_0_5_928 ();
 sg13g2_fill_8 FILLER_0_5_936 ();
 sg13g2_fill_8 FILLER_0_5_944 ();
 sg13g2_fill_8 FILLER_0_5_952 ();
 sg13g2_fill_8 FILLER_0_5_960 ();
 sg13g2_fill_8 FILLER_0_5_968 ();
 sg13g2_fill_8 FILLER_0_5_976 ();
 sg13g2_fill_8 FILLER_0_5_984 ();
 sg13g2_fill_8 FILLER_0_5_992 ();
 sg13g2_fill_8 FILLER_0_5_1000 ();
 sg13g2_fill_8 FILLER_0_5_1008 ();
 sg13g2_fill_8 FILLER_0_5_1016 ();
 sg13g2_fill_8 FILLER_0_5_1024 ();
 sg13g2_fill_8 FILLER_0_5_1032 ();
 sg13g2_fill_8 FILLER_0_5_1040 ();
 sg13g2_fill_8 FILLER_0_5_1048 ();
 sg13g2_fill_8 FILLER_0_5_1056 ();
 sg13g2_fill_8 FILLER_0_5_1064 ();
 sg13g2_fill_8 FILLER_0_5_1072 ();
 sg13g2_fill_8 FILLER_0_5_1080 ();
 sg13g2_fill_8 FILLER_0_5_1088 ();
 sg13g2_fill_8 FILLER_0_5_1096 ();
 sg13g2_fill_8 FILLER_0_5_1104 ();
 sg13g2_fill_8 FILLER_0_5_1112 ();
 sg13g2_fill_8 FILLER_0_5_1120 ();
 sg13g2_fill_8 FILLER_0_5_1128 ();
 sg13g2_fill_8 FILLER_0_5_1136 ();
 sg13g2_fill_8 FILLER_0_5_1144 ();
 sg13g2_fill_8 FILLER_0_5_1152 ();
 sg13g2_fill_8 FILLER_0_5_1160 ();
 sg13g2_fill_8 FILLER_0_5_1168 ();
 sg13g2_fill_8 FILLER_0_5_1176 ();
 sg13g2_fill_8 FILLER_0_5_1184 ();
 sg13g2_fill_8 FILLER_0_5_1192 ();
 sg13g2_fill_8 FILLER_0_5_1200 ();
 sg13g2_fill_8 FILLER_0_5_1208 ();
 sg13g2_fill_8 FILLER_0_5_1216 ();
 sg13g2_fill_4 FILLER_0_5_1224 ();
 sg13g2_fill_8 FILLER_0_6_0 ();
 sg13g2_fill_8 FILLER_0_6_8 ();
 sg13g2_fill_8 FILLER_0_6_16 ();
 sg13g2_fill_8 FILLER_0_6_24 ();
 sg13g2_fill_8 FILLER_0_6_32 ();
 sg13g2_fill_8 FILLER_0_6_40 ();
 sg13g2_fill_8 FILLER_0_6_48 ();
 sg13g2_fill_8 FILLER_0_6_56 ();
 sg13g2_fill_8 FILLER_0_6_64 ();
 sg13g2_fill_8 FILLER_0_6_72 ();
 sg13g2_fill_8 FILLER_0_6_80 ();
 sg13g2_fill_8 FILLER_0_6_88 ();
 sg13g2_fill_8 FILLER_0_6_96 ();
 sg13g2_fill_8 FILLER_0_6_104 ();
 sg13g2_fill_8 FILLER_0_6_112 ();
 sg13g2_fill_8 FILLER_0_6_120 ();
 sg13g2_fill_8 FILLER_0_6_128 ();
 sg13g2_fill_8 FILLER_0_6_136 ();
 sg13g2_fill_8 FILLER_0_6_144 ();
 sg13g2_fill_8 FILLER_0_6_152 ();
 sg13g2_fill_8 FILLER_0_6_160 ();
 sg13g2_fill_8 FILLER_0_6_168 ();
 sg13g2_fill_8 FILLER_0_6_176 ();
 sg13g2_fill_8 FILLER_0_6_184 ();
 sg13g2_fill_8 FILLER_0_6_192 ();
 sg13g2_fill_8 FILLER_0_6_200 ();
 sg13g2_fill_8 FILLER_0_6_208 ();
 sg13g2_fill_8 FILLER_0_6_216 ();
 sg13g2_fill_8 FILLER_0_6_224 ();
 sg13g2_fill_8 FILLER_0_6_232 ();
 sg13g2_fill_8 FILLER_0_6_240 ();
 sg13g2_fill_8 FILLER_0_6_248 ();
 sg13g2_fill_8 FILLER_0_6_256 ();
 sg13g2_fill_8 FILLER_0_6_264 ();
 sg13g2_fill_8 FILLER_0_6_272 ();
 sg13g2_fill_8 FILLER_0_6_280 ();
 sg13g2_fill_8 FILLER_0_6_288 ();
 sg13g2_fill_8 FILLER_0_6_296 ();
 sg13g2_fill_8 FILLER_0_6_304 ();
 sg13g2_fill_8 FILLER_0_6_312 ();
 sg13g2_fill_8 FILLER_0_6_320 ();
 sg13g2_fill_8 FILLER_0_6_328 ();
 sg13g2_fill_8 FILLER_0_6_336 ();
 sg13g2_fill_8 FILLER_0_6_344 ();
 sg13g2_fill_8 FILLER_0_6_352 ();
 sg13g2_fill_8 FILLER_0_6_360 ();
 sg13g2_fill_8 FILLER_0_6_368 ();
 sg13g2_fill_8 FILLER_0_6_376 ();
 sg13g2_fill_8 FILLER_0_6_384 ();
 sg13g2_fill_8 FILLER_0_6_392 ();
 sg13g2_fill_8 FILLER_0_6_400 ();
 sg13g2_fill_8 FILLER_0_6_408 ();
 sg13g2_fill_8 FILLER_0_6_416 ();
 sg13g2_fill_8 FILLER_0_6_424 ();
 sg13g2_fill_8 FILLER_0_6_432 ();
 sg13g2_fill_8 FILLER_0_6_440 ();
 sg13g2_fill_8 FILLER_0_6_448 ();
 sg13g2_fill_8 FILLER_0_6_456 ();
 sg13g2_fill_8 FILLER_0_6_464 ();
 sg13g2_fill_8 FILLER_0_6_472 ();
 sg13g2_fill_8 FILLER_0_6_480 ();
 sg13g2_fill_8 FILLER_0_6_488 ();
 sg13g2_fill_8 FILLER_0_6_496 ();
 sg13g2_fill_8 FILLER_0_6_504 ();
 sg13g2_fill_8 FILLER_0_6_512 ();
 sg13g2_fill_8 FILLER_0_6_520 ();
 sg13g2_fill_8 FILLER_0_6_528 ();
 sg13g2_fill_8 FILLER_0_6_536 ();
 sg13g2_fill_8 FILLER_0_6_544 ();
 sg13g2_fill_8 FILLER_0_6_552 ();
 sg13g2_fill_8 FILLER_0_6_560 ();
 sg13g2_fill_8 FILLER_0_6_568 ();
 sg13g2_fill_8 FILLER_0_6_576 ();
 sg13g2_fill_8 FILLER_0_6_584 ();
 sg13g2_fill_8 FILLER_0_6_592 ();
 sg13g2_fill_8 FILLER_0_6_600 ();
 sg13g2_fill_8 FILLER_0_6_608 ();
 sg13g2_fill_8 FILLER_0_6_616 ();
 sg13g2_fill_8 FILLER_0_6_624 ();
 sg13g2_fill_8 FILLER_0_6_632 ();
 sg13g2_fill_8 FILLER_0_6_640 ();
 sg13g2_fill_8 FILLER_0_6_648 ();
 sg13g2_fill_8 FILLER_0_6_656 ();
 sg13g2_fill_8 FILLER_0_6_664 ();
 sg13g2_fill_8 FILLER_0_6_672 ();
 sg13g2_fill_8 FILLER_0_6_680 ();
 sg13g2_fill_8 FILLER_0_6_688 ();
 sg13g2_fill_8 FILLER_0_6_696 ();
 sg13g2_fill_8 FILLER_0_6_704 ();
 sg13g2_fill_8 FILLER_0_6_712 ();
 sg13g2_fill_8 FILLER_0_6_720 ();
 sg13g2_fill_8 FILLER_0_6_728 ();
 sg13g2_fill_8 FILLER_0_6_736 ();
 sg13g2_fill_8 FILLER_0_6_744 ();
 sg13g2_fill_8 FILLER_0_6_752 ();
 sg13g2_fill_8 FILLER_0_6_760 ();
 sg13g2_fill_8 FILLER_0_6_768 ();
 sg13g2_fill_8 FILLER_0_6_776 ();
 sg13g2_fill_8 FILLER_0_6_784 ();
 sg13g2_fill_8 FILLER_0_6_792 ();
 sg13g2_fill_8 FILLER_0_6_800 ();
 sg13g2_fill_8 FILLER_0_6_808 ();
 sg13g2_fill_8 FILLER_0_6_816 ();
 sg13g2_fill_8 FILLER_0_6_824 ();
 sg13g2_fill_8 FILLER_0_6_832 ();
 sg13g2_fill_8 FILLER_0_6_840 ();
 sg13g2_fill_8 FILLER_0_6_848 ();
 sg13g2_fill_8 FILLER_0_6_856 ();
 sg13g2_fill_8 FILLER_0_6_864 ();
 sg13g2_fill_8 FILLER_0_6_872 ();
 sg13g2_fill_8 FILLER_0_6_880 ();
 sg13g2_fill_8 FILLER_0_6_888 ();
 sg13g2_fill_8 FILLER_0_6_896 ();
 sg13g2_fill_8 FILLER_0_6_904 ();
 sg13g2_fill_8 FILLER_0_6_912 ();
 sg13g2_fill_8 FILLER_0_6_920 ();
 sg13g2_fill_8 FILLER_0_6_928 ();
 sg13g2_fill_8 FILLER_0_6_936 ();
 sg13g2_fill_8 FILLER_0_6_944 ();
 sg13g2_fill_8 FILLER_0_6_952 ();
 sg13g2_fill_8 FILLER_0_6_960 ();
 sg13g2_fill_8 FILLER_0_6_968 ();
 sg13g2_fill_8 FILLER_0_6_976 ();
 sg13g2_fill_8 FILLER_0_6_984 ();
 sg13g2_fill_8 FILLER_0_6_992 ();
 sg13g2_fill_8 FILLER_0_6_1000 ();
 sg13g2_fill_8 FILLER_0_6_1008 ();
 sg13g2_fill_8 FILLER_0_6_1016 ();
 sg13g2_fill_8 FILLER_0_6_1024 ();
 sg13g2_fill_8 FILLER_0_6_1032 ();
 sg13g2_fill_8 FILLER_0_6_1040 ();
 sg13g2_fill_8 FILLER_0_6_1048 ();
 sg13g2_fill_8 FILLER_0_6_1056 ();
 sg13g2_fill_8 FILLER_0_6_1064 ();
 sg13g2_fill_8 FILLER_0_6_1072 ();
 sg13g2_fill_8 FILLER_0_6_1080 ();
 sg13g2_fill_8 FILLER_0_6_1088 ();
 sg13g2_fill_8 FILLER_0_6_1096 ();
 sg13g2_fill_8 FILLER_0_6_1104 ();
 sg13g2_fill_8 FILLER_0_6_1112 ();
 sg13g2_fill_8 FILLER_0_6_1120 ();
 sg13g2_fill_8 FILLER_0_6_1128 ();
 sg13g2_fill_8 FILLER_0_6_1136 ();
 sg13g2_fill_8 FILLER_0_6_1144 ();
 sg13g2_fill_8 FILLER_0_6_1152 ();
 sg13g2_fill_8 FILLER_0_6_1160 ();
 sg13g2_fill_8 FILLER_0_6_1168 ();
 sg13g2_fill_8 FILLER_0_6_1176 ();
 sg13g2_fill_8 FILLER_0_6_1184 ();
 sg13g2_fill_8 FILLER_0_6_1192 ();
 sg13g2_fill_8 FILLER_0_6_1200 ();
 sg13g2_fill_8 FILLER_0_6_1208 ();
 sg13g2_fill_8 FILLER_0_6_1216 ();
 sg13g2_fill_4 FILLER_0_6_1224 ();
 sg13g2_fill_8 FILLER_0_7_0 ();
 sg13g2_fill_8 FILLER_0_7_8 ();
 sg13g2_fill_8 FILLER_0_7_16 ();
 sg13g2_fill_8 FILLER_0_7_24 ();
 sg13g2_fill_8 FILLER_0_7_32 ();
 sg13g2_fill_8 FILLER_0_7_40 ();
 sg13g2_fill_8 FILLER_0_7_48 ();
 sg13g2_fill_8 FILLER_0_7_56 ();
 sg13g2_fill_8 FILLER_0_7_64 ();
 sg13g2_fill_8 FILLER_0_7_72 ();
 sg13g2_fill_8 FILLER_0_7_80 ();
 sg13g2_fill_8 FILLER_0_7_88 ();
 sg13g2_fill_8 FILLER_0_7_96 ();
 sg13g2_fill_8 FILLER_0_7_104 ();
 sg13g2_fill_8 FILLER_0_7_112 ();
 sg13g2_fill_8 FILLER_0_7_120 ();
 sg13g2_fill_8 FILLER_0_7_128 ();
 sg13g2_fill_8 FILLER_0_7_136 ();
 sg13g2_fill_8 FILLER_0_7_144 ();
 sg13g2_fill_8 FILLER_0_7_152 ();
 sg13g2_fill_8 FILLER_0_7_160 ();
 sg13g2_fill_8 FILLER_0_7_168 ();
 sg13g2_fill_8 FILLER_0_7_176 ();
 sg13g2_fill_8 FILLER_0_7_184 ();
 sg13g2_fill_8 FILLER_0_7_192 ();
 sg13g2_fill_8 FILLER_0_7_200 ();
 sg13g2_fill_8 FILLER_0_7_208 ();
 sg13g2_fill_8 FILLER_0_7_216 ();
 sg13g2_fill_8 FILLER_0_7_224 ();
 sg13g2_fill_8 FILLER_0_7_232 ();
 sg13g2_fill_8 FILLER_0_7_240 ();
 sg13g2_fill_8 FILLER_0_7_248 ();
 sg13g2_fill_8 FILLER_0_7_256 ();
 sg13g2_fill_8 FILLER_0_7_264 ();
 sg13g2_fill_8 FILLER_0_7_272 ();
 sg13g2_fill_8 FILLER_0_7_280 ();
 sg13g2_fill_8 FILLER_0_7_288 ();
 sg13g2_fill_8 FILLER_0_7_296 ();
 sg13g2_fill_8 FILLER_0_7_304 ();
 sg13g2_fill_8 FILLER_0_7_312 ();
 sg13g2_fill_8 FILLER_0_7_320 ();
 sg13g2_fill_8 FILLER_0_7_328 ();
 sg13g2_fill_8 FILLER_0_7_336 ();
 sg13g2_fill_8 FILLER_0_7_344 ();
 sg13g2_fill_8 FILLER_0_7_352 ();
 sg13g2_fill_8 FILLER_0_7_360 ();
 sg13g2_fill_8 FILLER_0_7_368 ();
 sg13g2_fill_8 FILLER_0_7_376 ();
 sg13g2_fill_8 FILLER_0_7_384 ();
 sg13g2_fill_8 FILLER_0_7_392 ();
 sg13g2_fill_8 FILLER_0_7_400 ();
 sg13g2_fill_8 FILLER_0_7_408 ();
 sg13g2_fill_8 FILLER_0_7_416 ();
 sg13g2_fill_8 FILLER_0_7_424 ();
 sg13g2_fill_8 FILLER_0_7_432 ();
 sg13g2_fill_8 FILLER_0_7_440 ();
 sg13g2_fill_8 FILLER_0_7_448 ();
 sg13g2_fill_8 FILLER_0_7_456 ();
 sg13g2_fill_8 FILLER_0_7_464 ();
 sg13g2_fill_8 FILLER_0_7_472 ();
 sg13g2_fill_8 FILLER_0_7_480 ();
 sg13g2_fill_8 FILLER_0_7_488 ();
 sg13g2_fill_8 FILLER_0_7_496 ();
 sg13g2_fill_8 FILLER_0_7_504 ();
 sg13g2_fill_8 FILLER_0_7_512 ();
 sg13g2_fill_8 FILLER_0_7_520 ();
 sg13g2_fill_8 FILLER_0_7_528 ();
 sg13g2_fill_8 FILLER_0_7_536 ();
 sg13g2_fill_8 FILLER_0_7_544 ();
 sg13g2_fill_8 FILLER_0_7_552 ();
 sg13g2_fill_8 FILLER_0_7_560 ();
 sg13g2_fill_8 FILLER_0_7_568 ();
 sg13g2_fill_8 FILLER_0_7_576 ();
 sg13g2_fill_8 FILLER_0_7_584 ();
 sg13g2_fill_8 FILLER_0_7_592 ();
 sg13g2_fill_8 FILLER_0_7_600 ();
 sg13g2_fill_8 FILLER_0_7_608 ();
 sg13g2_fill_8 FILLER_0_7_616 ();
 sg13g2_fill_8 FILLER_0_7_624 ();
 sg13g2_fill_8 FILLER_0_7_632 ();
 sg13g2_fill_8 FILLER_0_7_640 ();
 sg13g2_fill_8 FILLER_0_7_648 ();
 sg13g2_fill_8 FILLER_0_7_656 ();
 sg13g2_fill_8 FILLER_0_7_664 ();
 sg13g2_fill_8 FILLER_0_7_672 ();
 sg13g2_fill_8 FILLER_0_7_680 ();
 sg13g2_fill_8 FILLER_0_7_688 ();
 sg13g2_fill_8 FILLER_0_7_696 ();
 sg13g2_fill_8 FILLER_0_7_704 ();
 sg13g2_fill_8 FILLER_0_7_712 ();
 sg13g2_fill_8 FILLER_0_7_720 ();
 sg13g2_fill_8 FILLER_0_7_728 ();
 sg13g2_fill_8 FILLER_0_7_736 ();
 sg13g2_fill_8 FILLER_0_7_744 ();
 sg13g2_fill_8 FILLER_0_7_752 ();
 sg13g2_fill_8 FILLER_0_7_760 ();
 sg13g2_fill_8 FILLER_0_7_768 ();
 sg13g2_fill_8 FILLER_0_7_776 ();
 sg13g2_fill_8 FILLER_0_7_784 ();
 sg13g2_fill_8 FILLER_0_7_792 ();
 sg13g2_fill_8 FILLER_0_7_800 ();
 sg13g2_fill_8 FILLER_0_7_808 ();
 sg13g2_fill_8 FILLER_0_7_816 ();
 sg13g2_fill_8 FILLER_0_7_824 ();
 sg13g2_fill_8 FILLER_0_7_832 ();
 sg13g2_fill_8 FILLER_0_7_840 ();
 sg13g2_fill_8 FILLER_0_7_848 ();
 sg13g2_fill_8 FILLER_0_7_856 ();
 sg13g2_fill_8 FILLER_0_7_864 ();
 sg13g2_fill_8 FILLER_0_7_872 ();
 sg13g2_fill_8 FILLER_0_7_880 ();
 sg13g2_fill_8 FILLER_0_7_888 ();
 sg13g2_fill_8 FILLER_0_7_896 ();
 sg13g2_fill_8 FILLER_0_7_904 ();
 sg13g2_fill_8 FILLER_0_7_912 ();
 sg13g2_fill_8 FILLER_0_7_920 ();
 sg13g2_fill_8 FILLER_0_7_928 ();
 sg13g2_fill_8 FILLER_0_7_936 ();
 sg13g2_fill_8 FILLER_0_7_944 ();
 sg13g2_fill_8 FILLER_0_7_952 ();
 sg13g2_fill_8 FILLER_0_7_960 ();
 sg13g2_fill_8 FILLER_0_7_968 ();
 sg13g2_fill_8 FILLER_0_7_976 ();
 sg13g2_fill_8 FILLER_0_7_984 ();
 sg13g2_fill_8 FILLER_0_7_992 ();
 sg13g2_fill_8 FILLER_0_7_1000 ();
 sg13g2_fill_8 FILLER_0_7_1008 ();
 sg13g2_fill_8 FILLER_0_7_1016 ();
 sg13g2_fill_8 FILLER_0_7_1024 ();
 sg13g2_fill_8 FILLER_0_7_1032 ();
 sg13g2_fill_8 FILLER_0_7_1040 ();
 sg13g2_fill_8 FILLER_0_7_1048 ();
 sg13g2_fill_8 FILLER_0_7_1056 ();
 sg13g2_fill_8 FILLER_0_7_1064 ();
 sg13g2_fill_8 FILLER_0_7_1072 ();
 sg13g2_fill_8 FILLER_0_7_1080 ();
 sg13g2_fill_8 FILLER_0_7_1088 ();
 sg13g2_fill_8 FILLER_0_7_1096 ();
 sg13g2_fill_8 FILLER_0_7_1104 ();
 sg13g2_fill_8 FILLER_0_7_1112 ();
 sg13g2_fill_8 FILLER_0_7_1120 ();
 sg13g2_fill_8 FILLER_0_7_1128 ();
 sg13g2_fill_8 FILLER_0_7_1136 ();
 sg13g2_fill_8 FILLER_0_7_1144 ();
 sg13g2_fill_8 FILLER_0_7_1152 ();
 sg13g2_fill_8 FILLER_0_7_1160 ();
 sg13g2_fill_8 FILLER_0_7_1168 ();
 sg13g2_fill_8 FILLER_0_7_1176 ();
 sg13g2_fill_8 FILLER_0_7_1184 ();
 sg13g2_fill_8 FILLER_0_7_1192 ();
 sg13g2_fill_8 FILLER_0_7_1200 ();
 sg13g2_fill_8 FILLER_0_7_1208 ();
 sg13g2_fill_8 FILLER_0_7_1216 ();
 sg13g2_fill_4 FILLER_0_7_1224 ();
 sg13g2_fill_8 FILLER_0_8_0 ();
 sg13g2_fill_8 FILLER_0_8_8 ();
 sg13g2_fill_8 FILLER_0_8_16 ();
 sg13g2_fill_8 FILLER_0_8_24 ();
 sg13g2_fill_8 FILLER_0_8_32 ();
 sg13g2_fill_8 FILLER_0_8_40 ();
 sg13g2_fill_8 FILLER_0_8_48 ();
 sg13g2_fill_8 FILLER_0_8_56 ();
 sg13g2_fill_8 FILLER_0_8_64 ();
 sg13g2_fill_8 FILLER_0_8_72 ();
 sg13g2_fill_8 FILLER_0_8_80 ();
 sg13g2_fill_8 FILLER_0_8_88 ();
 sg13g2_fill_8 FILLER_0_8_96 ();
 sg13g2_fill_8 FILLER_0_8_104 ();
 sg13g2_fill_8 FILLER_0_8_112 ();
 sg13g2_fill_8 FILLER_0_8_120 ();
 sg13g2_fill_8 FILLER_0_8_128 ();
 sg13g2_fill_8 FILLER_0_8_136 ();
 sg13g2_fill_8 FILLER_0_8_144 ();
 sg13g2_fill_8 FILLER_0_8_152 ();
 sg13g2_fill_8 FILLER_0_8_160 ();
 sg13g2_fill_8 FILLER_0_8_168 ();
 sg13g2_fill_8 FILLER_0_8_176 ();
 sg13g2_fill_8 FILLER_0_8_184 ();
 sg13g2_fill_8 FILLER_0_8_192 ();
 sg13g2_fill_8 FILLER_0_8_200 ();
 sg13g2_fill_8 FILLER_0_8_208 ();
 sg13g2_fill_8 FILLER_0_8_216 ();
 sg13g2_fill_8 FILLER_0_8_224 ();
 sg13g2_fill_8 FILLER_0_8_232 ();
 sg13g2_fill_8 FILLER_0_8_240 ();
 sg13g2_fill_8 FILLER_0_8_248 ();
 sg13g2_fill_8 FILLER_0_8_256 ();
 sg13g2_fill_8 FILLER_0_8_264 ();
 sg13g2_fill_8 FILLER_0_8_272 ();
 sg13g2_fill_8 FILLER_0_8_280 ();
 sg13g2_fill_8 FILLER_0_8_288 ();
 sg13g2_fill_8 FILLER_0_8_296 ();
 sg13g2_fill_8 FILLER_0_8_304 ();
 sg13g2_fill_8 FILLER_0_8_312 ();
 sg13g2_fill_8 FILLER_0_8_320 ();
 sg13g2_fill_8 FILLER_0_8_328 ();
 sg13g2_fill_8 FILLER_0_8_336 ();
 sg13g2_fill_8 FILLER_0_8_344 ();
 sg13g2_fill_8 FILLER_0_8_352 ();
 sg13g2_fill_8 FILLER_0_8_360 ();
 sg13g2_fill_8 FILLER_0_8_368 ();
 sg13g2_fill_8 FILLER_0_8_376 ();
 sg13g2_fill_8 FILLER_0_8_384 ();
 sg13g2_fill_8 FILLER_0_8_392 ();
 sg13g2_fill_8 FILLER_0_8_400 ();
 sg13g2_fill_8 FILLER_0_8_408 ();
 sg13g2_fill_8 FILLER_0_8_416 ();
 sg13g2_fill_8 FILLER_0_8_424 ();
 sg13g2_fill_8 FILLER_0_8_432 ();
 sg13g2_fill_8 FILLER_0_8_440 ();
 sg13g2_fill_8 FILLER_0_8_448 ();
 sg13g2_fill_8 FILLER_0_8_456 ();
 sg13g2_fill_8 FILLER_0_8_464 ();
 sg13g2_fill_8 FILLER_0_8_472 ();
 sg13g2_fill_8 FILLER_0_8_480 ();
 sg13g2_fill_8 FILLER_0_8_488 ();
 sg13g2_fill_8 FILLER_0_8_496 ();
 sg13g2_fill_8 FILLER_0_8_504 ();
 sg13g2_fill_8 FILLER_0_8_512 ();
 sg13g2_fill_8 FILLER_0_8_520 ();
 sg13g2_fill_8 FILLER_0_8_528 ();
 sg13g2_fill_8 FILLER_0_8_536 ();
 sg13g2_fill_8 FILLER_0_8_544 ();
 sg13g2_fill_8 FILLER_0_8_552 ();
 sg13g2_fill_8 FILLER_0_8_560 ();
 sg13g2_fill_8 FILLER_0_8_568 ();
 sg13g2_fill_8 FILLER_0_8_576 ();
 sg13g2_fill_8 FILLER_0_8_584 ();
 sg13g2_fill_8 FILLER_0_8_592 ();
 sg13g2_fill_8 FILLER_0_8_600 ();
 sg13g2_fill_8 FILLER_0_8_608 ();
 sg13g2_fill_8 FILLER_0_8_616 ();
 sg13g2_fill_8 FILLER_0_8_624 ();
 sg13g2_fill_8 FILLER_0_8_632 ();
 sg13g2_fill_8 FILLER_0_8_640 ();
 sg13g2_fill_8 FILLER_0_8_648 ();
 sg13g2_fill_8 FILLER_0_8_656 ();
 sg13g2_fill_8 FILLER_0_8_664 ();
 sg13g2_fill_8 FILLER_0_8_672 ();
 sg13g2_fill_8 FILLER_0_8_680 ();
 sg13g2_fill_8 FILLER_0_8_688 ();
 sg13g2_fill_8 FILLER_0_8_696 ();
 sg13g2_fill_8 FILLER_0_8_704 ();
 sg13g2_fill_8 FILLER_0_8_712 ();
 sg13g2_fill_8 FILLER_0_8_720 ();
 sg13g2_fill_8 FILLER_0_8_728 ();
 sg13g2_fill_8 FILLER_0_8_736 ();
 sg13g2_fill_8 FILLER_0_8_744 ();
 sg13g2_fill_8 FILLER_0_8_752 ();
 sg13g2_fill_8 FILLER_0_8_760 ();
 sg13g2_fill_8 FILLER_0_8_768 ();
 sg13g2_fill_8 FILLER_0_8_776 ();
 sg13g2_fill_8 FILLER_0_8_784 ();
 sg13g2_fill_8 FILLER_0_8_792 ();
 sg13g2_fill_8 FILLER_0_8_800 ();
 sg13g2_fill_8 FILLER_0_8_808 ();
 sg13g2_fill_8 FILLER_0_8_816 ();
 sg13g2_fill_8 FILLER_0_8_824 ();
 sg13g2_fill_8 FILLER_0_8_832 ();
 sg13g2_fill_8 FILLER_0_8_840 ();
 sg13g2_fill_8 FILLER_0_8_848 ();
 sg13g2_fill_8 FILLER_0_8_856 ();
 sg13g2_fill_8 FILLER_0_8_864 ();
 sg13g2_fill_8 FILLER_0_8_872 ();
 sg13g2_fill_8 FILLER_0_8_880 ();
 sg13g2_fill_8 FILLER_0_8_888 ();
 sg13g2_fill_8 FILLER_0_8_896 ();
 sg13g2_fill_8 FILLER_0_8_904 ();
 sg13g2_fill_8 FILLER_0_8_912 ();
 sg13g2_fill_8 FILLER_0_8_920 ();
 sg13g2_fill_8 FILLER_0_8_928 ();
 sg13g2_fill_8 FILLER_0_8_936 ();
 sg13g2_fill_8 FILLER_0_8_944 ();
 sg13g2_fill_8 FILLER_0_8_952 ();
 sg13g2_fill_8 FILLER_0_8_960 ();
 sg13g2_fill_8 FILLER_0_8_968 ();
 sg13g2_fill_8 FILLER_0_8_976 ();
 sg13g2_fill_8 FILLER_0_8_984 ();
 sg13g2_fill_8 FILLER_0_8_992 ();
 sg13g2_fill_8 FILLER_0_8_1000 ();
 sg13g2_fill_8 FILLER_0_8_1008 ();
 sg13g2_fill_8 FILLER_0_8_1016 ();
 sg13g2_fill_8 FILLER_0_8_1024 ();
 sg13g2_fill_8 FILLER_0_8_1032 ();
 sg13g2_fill_8 FILLER_0_8_1040 ();
 sg13g2_fill_8 FILLER_0_8_1048 ();
 sg13g2_fill_8 FILLER_0_8_1056 ();
 sg13g2_fill_8 FILLER_0_8_1064 ();
 sg13g2_fill_8 FILLER_0_8_1072 ();
 sg13g2_fill_8 FILLER_0_8_1080 ();
 sg13g2_fill_8 FILLER_0_8_1088 ();
 sg13g2_fill_8 FILLER_0_8_1096 ();
 sg13g2_fill_8 FILLER_0_8_1104 ();
 sg13g2_fill_8 FILLER_0_8_1112 ();
 sg13g2_fill_8 FILLER_0_8_1120 ();
 sg13g2_fill_8 FILLER_0_8_1128 ();
 sg13g2_fill_8 FILLER_0_8_1136 ();
 sg13g2_fill_8 FILLER_0_8_1144 ();
 sg13g2_fill_8 FILLER_0_8_1152 ();
 sg13g2_fill_8 FILLER_0_8_1160 ();
 sg13g2_fill_8 FILLER_0_8_1168 ();
 sg13g2_fill_8 FILLER_0_8_1176 ();
 sg13g2_fill_8 FILLER_0_8_1184 ();
 sg13g2_fill_8 FILLER_0_8_1192 ();
 sg13g2_fill_8 FILLER_0_8_1200 ();
 sg13g2_fill_8 FILLER_0_8_1208 ();
 sg13g2_fill_8 FILLER_0_8_1216 ();
 sg13g2_fill_4 FILLER_0_8_1224 ();
 sg13g2_fill_8 FILLER_0_9_0 ();
 sg13g2_fill_8 FILLER_0_9_8 ();
 sg13g2_fill_8 FILLER_0_9_16 ();
 sg13g2_fill_8 FILLER_0_9_24 ();
 sg13g2_fill_8 FILLER_0_9_32 ();
 sg13g2_fill_8 FILLER_0_9_40 ();
 sg13g2_fill_8 FILLER_0_9_48 ();
 sg13g2_fill_8 FILLER_0_9_56 ();
 sg13g2_fill_8 FILLER_0_9_64 ();
 sg13g2_fill_8 FILLER_0_9_72 ();
 sg13g2_fill_8 FILLER_0_9_80 ();
 sg13g2_fill_8 FILLER_0_9_88 ();
 sg13g2_fill_8 FILLER_0_9_96 ();
 sg13g2_fill_8 FILLER_0_9_104 ();
 sg13g2_fill_8 FILLER_0_9_112 ();
 sg13g2_fill_8 FILLER_0_9_120 ();
 sg13g2_fill_8 FILLER_0_9_128 ();
 sg13g2_fill_8 FILLER_0_9_136 ();
 sg13g2_fill_8 FILLER_0_9_144 ();
 sg13g2_fill_8 FILLER_0_9_152 ();
 sg13g2_fill_8 FILLER_0_9_160 ();
 sg13g2_fill_8 FILLER_0_9_168 ();
 sg13g2_fill_8 FILLER_0_9_176 ();
 sg13g2_fill_8 FILLER_0_9_184 ();
 sg13g2_fill_8 FILLER_0_9_192 ();
 sg13g2_fill_8 FILLER_0_9_200 ();
 sg13g2_fill_8 FILLER_0_9_208 ();
 sg13g2_fill_8 FILLER_0_9_216 ();
 sg13g2_fill_8 FILLER_0_9_224 ();
 sg13g2_fill_8 FILLER_0_9_232 ();
 sg13g2_fill_8 FILLER_0_9_240 ();
 sg13g2_fill_8 FILLER_0_9_248 ();
 sg13g2_fill_8 FILLER_0_9_256 ();
 sg13g2_fill_8 FILLER_0_9_264 ();
 sg13g2_fill_8 FILLER_0_9_272 ();
 sg13g2_fill_8 FILLER_0_9_280 ();
 sg13g2_fill_8 FILLER_0_9_288 ();
 sg13g2_fill_8 FILLER_0_9_296 ();
 sg13g2_fill_8 FILLER_0_9_304 ();
 sg13g2_fill_8 FILLER_0_9_312 ();
 sg13g2_fill_8 FILLER_0_9_320 ();
 sg13g2_fill_8 FILLER_0_9_328 ();
 sg13g2_fill_8 FILLER_0_9_336 ();
 sg13g2_fill_8 FILLER_0_9_344 ();
 sg13g2_fill_8 FILLER_0_9_352 ();
 sg13g2_fill_8 FILLER_0_9_360 ();
 sg13g2_fill_8 FILLER_0_9_368 ();
 sg13g2_fill_8 FILLER_0_9_376 ();
 sg13g2_fill_8 FILLER_0_9_384 ();
 sg13g2_fill_8 FILLER_0_9_392 ();
 sg13g2_fill_8 FILLER_0_9_400 ();
 sg13g2_fill_8 FILLER_0_9_408 ();
 sg13g2_fill_8 FILLER_0_9_416 ();
 sg13g2_fill_8 FILLER_0_9_424 ();
 sg13g2_fill_8 FILLER_0_9_432 ();
 sg13g2_fill_8 FILLER_0_9_440 ();
 sg13g2_fill_8 FILLER_0_9_448 ();
 sg13g2_fill_8 FILLER_0_9_456 ();
 sg13g2_fill_8 FILLER_0_9_464 ();
 sg13g2_fill_8 FILLER_0_9_472 ();
 sg13g2_fill_8 FILLER_0_9_480 ();
 sg13g2_fill_8 FILLER_0_9_488 ();
 sg13g2_fill_8 FILLER_0_9_496 ();
 sg13g2_fill_8 FILLER_0_9_504 ();
 sg13g2_fill_8 FILLER_0_9_512 ();
 sg13g2_fill_8 FILLER_0_9_520 ();
 sg13g2_fill_8 FILLER_0_9_528 ();
 sg13g2_fill_8 FILLER_0_9_536 ();
 sg13g2_fill_8 FILLER_0_9_544 ();
 sg13g2_fill_8 FILLER_0_9_552 ();
 sg13g2_fill_8 FILLER_0_9_560 ();
 sg13g2_fill_8 FILLER_0_9_568 ();
 sg13g2_fill_8 FILLER_0_9_576 ();
 sg13g2_fill_8 FILLER_0_9_584 ();
 sg13g2_fill_8 FILLER_0_9_592 ();
 sg13g2_fill_8 FILLER_0_9_600 ();
 sg13g2_fill_8 FILLER_0_9_608 ();
 sg13g2_fill_8 FILLER_0_9_616 ();
 sg13g2_fill_8 FILLER_0_9_624 ();
 sg13g2_fill_8 FILLER_0_9_632 ();
 sg13g2_fill_8 FILLER_0_9_640 ();
 sg13g2_fill_8 FILLER_0_9_648 ();
 sg13g2_fill_8 FILLER_0_9_656 ();
 sg13g2_fill_8 FILLER_0_9_664 ();
 sg13g2_fill_8 FILLER_0_9_672 ();
 sg13g2_fill_8 FILLER_0_9_680 ();
 sg13g2_fill_8 FILLER_0_9_688 ();
 sg13g2_fill_8 FILLER_0_9_696 ();
 sg13g2_fill_8 FILLER_0_9_704 ();
 sg13g2_fill_8 FILLER_0_9_712 ();
 sg13g2_fill_8 FILLER_0_9_720 ();
 sg13g2_fill_8 FILLER_0_9_728 ();
 sg13g2_fill_8 FILLER_0_9_736 ();
 sg13g2_fill_8 FILLER_0_9_744 ();
 sg13g2_fill_8 FILLER_0_9_752 ();
 sg13g2_fill_8 FILLER_0_9_760 ();
 sg13g2_fill_8 FILLER_0_9_768 ();
 sg13g2_fill_8 FILLER_0_9_776 ();
 sg13g2_fill_8 FILLER_0_9_784 ();
 sg13g2_fill_8 FILLER_0_9_792 ();
 sg13g2_fill_8 FILLER_0_9_800 ();
 sg13g2_fill_8 FILLER_0_9_808 ();
 sg13g2_fill_8 FILLER_0_9_816 ();
 sg13g2_fill_8 FILLER_0_9_824 ();
 sg13g2_fill_8 FILLER_0_9_832 ();
 sg13g2_fill_8 FILLER_0_9_840 ();
 sg13g2_fill_8 FILLER_0_9_848 ();
 sg13g2_fill_8 FILLER_0_9_856 ();
 sg13g2_fill_8 FILLER_0_9_864 ();
 sg13g2_fill_8 FILLER_0_9_872 ();
 sg13g2_fill_8 FILLER_0_9_880 ();
 sg13g2_fill_8 FILLER_0_9_888 ();
 sg13g2_fill_8 FILLER_0_9_896 ();
 sg13g2_fill_8 FILLER_0_9_904 ();
 sg13g2_fill_8 FILLER_0_9_912 ();
 sg13g2_fill_8 FILLER_0_9_920 ();
 sg13g2_fill_8 FILLER_0_9_928 ();
 sg13g2_fill_8 FILLER_0_9_936 ();
 sg13g2_fill_8 FILLER_0_9_944 ();
 sg13g2_fill_8 FILLER_0_9_952 ();
 sg13g2_fill_8 FILLER_0_9_960 ();
 sg13g2_fill_8 FILLER_0_9_968 ();
 sg13g2_fill_8 FILLER_0_9_976 ();
 sg13g2_fill_8 FILLER_0_9_984 ();
 sg13g2_fill_8 FILLER_0_9_992 ();
 sg13g2_fill_8 FILLER_0_9_1000 ();
 sg13g2_fill_8 FILLER_0_9_1008 ();
 sg13g2_fill_8 FILLER_0_9_1016 ();
 sg13g2_fill_8 FILLER_0_9_1024 ();
 sg13g2_fill_8 FILLER_0_9_1032 ();
 sg13g2_fill_8 FILLER_0_9_1040 ();
 sg13g2_fill_8 FILLER_0_9_1048 ();
 sg13g2_fill_8 FILLER_0_9_1056 ();
 sg13g2_fill_8 FILLER_0_9_1064 ();
 sg13g2_fill_8 FILLER_0_9_1072 ();
 sg13g2_fill_8 FILLER_0_9_1080 ();
 sg13g2_fill_8 FILLER_0_9_1088 ();
 sg13g2_fill_8 FILLER_0_9_1096 ();
 sg13g2_fill_8 FILLER_0_9_1104 ();
 sg13g2_fill_8 FILLER_0_9_1112 ();
 sg13g2_fill_8 FILLER_0_9_1120 ();
 sg13g2_fill_8 FILLER_0_9_1128 ();
 sg13g2_fill_8 FILLER_0_9_1136 ();
 sg13g2_fill_8 FILLER_0_9_1144 ();
 sg13g2_fill_8 FILLER_0_9_1152 ();
 sg13g2_fill_8 FILLER_0_9_1160 ();
 sg13g2_fill_8 FILLER_0_9_1168 ();
 sg13g2_fill_8 FILLER_0_9_1176 ();
 sg13g2_fill_8 FILLER_0_9_1184 ();
 sg13g2_fill_8 FILLER_0_9_1192 ();
 sg13g2_fill_8 FILLER_0_9_1200 ();
 sg13g2_fill_8 FILLER_0_9_1208 ();
 sg13g2_fill_8 FILLER_0_9_1216 ();
 sg13g2_fill_4 FILLER_0_9_1224 ();
 sg13g2_fill_8 FILLER_0_10_0 ();
 sg13g2_fill_8 FILLER_0_10_8 ();
 sg13g2_fill_8 FILLER_0_10_16 ();
 sg13g2_fill_8 FILLER_0_10_24 ();
 sg13g2_fill_8 FILLER_0_10_32 ();
 sg13g2_fill_8 FILLER_0_10_40 ();
 sg13g2_fill_8 FILLER_0_10_48 ();
 sg13g2_fill_8 FILLER_0_10_56 ();
 sg13g2_fill_8 FILLER_0_10_64 ();
 sg13g2_fill_8 FILLER_0_10_72 ();
 sg13g2_fill_8 FILLER_0_10_80 ();
 sg13g2_fill_8 FILLER_0_10_88 ();
 sg13g2_fill_8 FILLER_0_10_96 ();
 sg13g2_fill_8 FILLER_0_10_104 ();
 sg13g2_fill_8 FILLER_0_10_112 ();
 sg13g2_fill_8 FILLER_0_10_120 ();
 sg13g2_fill_8 FILLER_0_10_128 ();
 sg13g2_fill_8 FILLER_0_10_136 ();
 sg13g2_fill_8 FILLER_0_10_144 ();
 sg13g2_fill_8 FILLER_0_10_152 ();
 sg13g2_fill_8 FILLER_0_10_160 ();
 sg13g2_fill_8 FILLER_0_10_168 ();
 sg13g2_fill_8 FILLER_0_10_176 ();
 sg13g2_fill_8 FILLER_0_10_184 ();
 sg13g2_fill_8 FILLER_0_10_192 ();
 sg13g2_fill_8 FILLER_0_10_200 ();
 sg13g2_fill_8 FILLER_0_10_208 ();
 sg13g2_fill_8 FILLER_0_10_216 ();
 sg13g2_fill_8 FILLER_0_10_224 ();
 sg13g2_fill_8 FILLER_0_10_232 ();
 sg13g2_fill_8 FILLER_0_10_240 ();
 sg13g2_fill_8 FILLER_0_10_248 ();
 sg13g2_fill_8 FILLER_0_10_256 ();
 sg13g2_fill_8 FILLER_0_10_264 ();
 sg13g2_fill_8 FILLER_0_10_272 ();
 sg13g2_fill_8 FILLER_0_10_280 ();
 sg13g2_fill_8 FILLER_0_10_288 ();
 sg13g2_fill_8 FILLER_0_10_296 ();
 sg13g2_fill_8 FILLER_0_10_304 ();
 sg13g2_fill_8 FILLER_0_10_312 ();
 sg13g2_fill_8 FILLER_0_10_320 ();
 sg13g2_fill_8 FILLER_0_10_328 ();
 sg13g2_fill_8 FILLER_0_10_336 ();
 sg13g2_fill_8 FILLER_0_10_344 ();
 sg13g2_fill_8 FILLER_0_10_352 ();
 sg13g2_fill_8 FILLER_0_10_360 ();
 sg13g2_fill_8 FILLER_0_10_368 ();
 sg13g2_fill_8 FILLER_0_10_376 ();
 sg13g2_fill_8 FILLER_0_10_384 ();
 sg13g2_fill_8 FILLER_0_10_392 ();
 sg13g2_fill_8 FILLER_0_10_400 ();
 sg13g2_fill_8 FILLER_0_10_408 ();
 sg13g2_fill_8 FILLER_0_10_416 ();
 sg13g2_fill_8 FILLER_0_10_424 ();
 sg13g2_fill_8 FILLER_0_10_432 ();
 sg13g2_fill_8 FILLER_0_10_440 ();
 sg13g2_fill_8 FILLER_0_10_448 ();
 sg13g2_fill_8 FILLER_0_10_456 ();
 sg13g2_fill_8 FILLER_0_10_464 ();
 sg13g2_fill_8 FILLER_0_10_472 ();
 sg13g2_fill_8 FILLER_0_10_480 ();
 sg13g2_fill_8 FILLER_0_10_488 ();
 sg13g2_fill_8 FILLER_0_10_496 ();
 sg13g2_fill_8 FILLER_0_10_504 ();
 sg13g2_fill_8 FILLER_0_10_512 ();
 sg13g2_fill_8 FILLER_0_10_520 ();
 sg13g2_fill_8 FILLER_0_10_528 ();
 sg13g2_fill_8 FILLER_0_10_536 ();
 sg13g2_fill_8 FILLER_0_10_544 ();
 sg13g2_fill_8 FILLER_0_10_552 ();
 sg13g2_fill_8 FILLER_0_10_560 ();
 sg13g2_fill_8 FILLER_0_10_568 ();
 sg13g2_fill_8 FILLER_0_10_576 ();
 sg13g2_fill_8 FILLER_0_10_584 ();
 sg13g2_fill_8 FILLER_0_10_592 ();
 sg13g2_fill_8 FILLER_0_10_600 ();
 sg13g2_fill_8 FILLER_0_10_608 ();
 sg13g2_fill_8 FILLER_0_10_616 ();
 sg13g2_fill_8 FILLER_0_10_624 ();
 sg13g2_fill_8 FILLER_0_10_632 ();
 sg13g2_fill_8 FILLER_0_10_640 ();
 sg13g2_fill_8 FILLER_0_10_648 ();
 sg13g2_fill_8 FILLER_0_10_656 ();
 sg13g2_fill_8 FILLER_0_10_664 ();
 sg13g2_fill_8 FILLER_0_10_672 ();
 sg13g2_fill_8 FILLER_0_10_680 ();
 sg13g2_fill_8 FILLER_0_10_688 ();
 sg13g2_fill_8 FILLER_0_10_696 ();
 sg13g2_fill_8 FILLER_0_10_704 ();
 sg13g2_fill_8 FILLER_0_10_712 ();
 sg13g2_fill_8 FILLER_0_10_720 ();
 sg13g2_fill_8 FILLER_0_10_728 ();
 sg13g2_fill_8 FILLER_0_10_736 ();
 sg13g2_fill_8 FILLER_0_10_744 ();
 sg13g2_fill_8 FILLER_0_10_752 ();
 sg13g2_fill_8 FILLER_0_10_760 ();
 sg13g2_fill_8 FILLER_0_10_768 ();
 sg13g2_fill_8 FILLER_0_10_776 ();
 sg13g2_fill_8 FILLER_0_10_784 ();
 sg13g2_fill_8 FILLER_0_10_792 ();
 sg13g2_fill_8 FILLER_0_10_800 ();
 sg13g2_fill_8 FILLER_0_10_808 ();
 sg13g2_fill_8 FILLER_0_10_816 ();
 sg13g2_fill_8 FILLER_0_10_824 ();
 sg13g2_fill_8 FILLER_0_10_832 ();
 sg13g2_fill_8 FILLER_0_10_840 ();
 sg13g2_fill_8 FILLER_0_10_848 ();
 sg13g2_fill_8 FILLER_0_10_856 ();
 sg13g2_fill_8 FILLER_0_10_864 ();
 sg13g2_fill_8 FILLER_0_10_872 ();
 sg13g2_fill_8 FILLER_0_10_880 ();
 sg13g2_fill_8 FILLER_0_10_888 ();
 sg13g2_fill_8 FILLER_0_10_896 ();
 sg13g2_fill_8 FILLER_0_10_904 ();
 sg13g2_fill_8 FILLER_0_10_912 ();
 sg13g2_fill_8 FILLER_0_10_920 ();
 sg13g2_fill_8 FILLER_0_10_928 ();
 sg13g2_fill_8 FILLER_0_10_936 ();
 sg13g2_fill_8 FILLER_0_10_944 ();
 sg13g2_fill_8 FILLER_0_10_952 ();
 sg13g2_fill_8 FILLER_0_10_960 ();
 sg13g2_fill_8 FILLER_0_10_968 ();
 sg13g2_fill_8 FILLER_0_10_976 ();
 sg13g2_fill_8 FILLER_0_10_984 ();
 sg13g2_fill_8 FILLER_0_10_992 ();
 sg13g2_fill_8 FILLER_0_10_1000 ();
 sg13g2_fill_8 FILLER_0_10_1008 ();
 sg13g2_fill_8 FILLER_0_10_1016 ();
 sg13g2_fill_8 FILLER_0_10_1024 ();
 sg13g2_fill_8 FILLER_0_10_1032 ();
 sg13g2_fill_8 FILLER_0_10_1040 ();
 sg13g2_fill_8 FILLER_0_10_1048 ();
 sg13g2_fill_8 FILLER_0_10_1056 ();
 sg13g2_fill_8 FILLER_0_10_1064 ();
 sg13g2_fill_8 FILLER_0_10_1072 ();
 sg13g2_fill_8 FILLER_0_10_1080 ();
 sg13g2_fill_8 FILLER_0_10_1088 ();
 sg13g2_fill_8 FILLER_0_10_1096 ();
 sg13g2_fill_8 FILLER_0_10_1104 ();
 sg13g2_fill_8 FILLER_0_10_1112 ();
 sg13g2_fill_8 FILLER_0_10_1120 ();
 sg13g2_fill_8 FILLER_0_10_1128 ();
 sg13g2_fill_8 FILLER_0_10_1136 ();
 sg13g2_fill_8 FILLER_0_10_1144 ();
 sg13g2_fill_8 FILLER_0_10_1152 ();
 sg13g2_fill_8 FILLER_0_10_1160 ();
 sg13g2_fill_8 FILLER_0_10_1168 ();
 sg13g2_fill_8 FILLER_0_10_1176 ();
 sg13g2_fill_8 FILLER_0_10_1184 ();
 sg13g2_fill_8 FILLER_0_10_1192 ();
 sg13g2_fill_8 FILLER_0_10_1200 ();
 sg13g2_fill_8 FILLER_0_10_1208 ();
 sg13g2_fill_8 FILLER_0_10_1216 ();
 sg13g2_fill_4 FILLER_0_10_1224 ();
 sg13g2_fill_8 FILLER_0_11_0 ();
 sg13g2_fill_8 FILLER_0_11_8 ();
 sg13g2_fill_8 FILLER_0_11_16 ();
 sg13g2_fill_8 FILLER_0_11_24 ();
 sg13g2_fill_8 FILLER_0_11_32 ();
 sg13g2_fill_8 FILLER_0_11_40 ();
 sg13g2_fill_8 FILLER_0_11_48 ();
 sg13g2_fill_8 FILLER_0_11_56 ();
 sg13g2_fill_8 FILLER_0_11_64 ();
 sg13g2_fill_8 FILLER_0_11_72 ();
 sg13g2_fill_8 FILLER_0_11_80 ();
 sg13g2_fill_8 FILLER_0_11_88 ();
 sg13g2_fill_8 FILLER_0_11_96 ();
 sg13g2_fill_8 FILLER_0_11_104 ();
 sg13g2_fill_8 FILLER_0_11_112 ();
 sg13g2_fill_8 FILLER_0_11_120 ();
 sg13g2_fill_8 FILLER_0_11_128 ();
 sg13g2_fill_8 FILLER_0_11_136 ();
 sg13g2_fill_8 FILLER_0_11_144 ();
 sg13g2_fill_8 FILLER_0_11_152 ();
 sg13g2_fill_8 FILLER_0_11_160 ();
 sg13g2_fill_8 FILLER_0_11_168 ();
 sg13g2_fill_8 FILLER_0_11_176 ();
 sg13g2_fill_8 FILLER_0_11_184 ();
 sg13g2_fill_8 FILLER_0_11_192 ();
 sg13g2_fill_8 FILLER_0_11_200 ();
 sg13g2_fill_8 FILLER_0_11_208 ();
 sg13g2_fill_8 FILLER_0_11_216 ();
 sg13g2_fill_8 FILLER_0_11_224 ();
 sg13g2_fill_8 FILLER_0_11_232 ();
 sg13g2_fill_8 FILLER_0_11_240 ();
 sg13g2_fill_8 FILLER_0_11_248 ();
 sg13g2_fill_8 FILLER_0_11_256 ();
 sg13g2_fill_8 FILLER_0_11_264 ();
 sg13g2_fill_8 FILLER_0_11_272 ();
 sg13g2_fill_8 FILLER_0_11_280 ();
 sg13g2_fill_8 FILLER_0_11_288 ();
 sg13g2_fill_8 FILLER_0_11_296 ();
 sg13g2_fill_8 FILLER_0_11_304 ();
 sg13g2_fill_8 FILLER_0_11_312 ();
 sg13g2_fill_8 FILLER_0_11_320 ();
 sg13g2_fill_8 FILLER_0_11_328 ();
 sg13g2_fill_8 FILLER_0_11_336 ();
 sg13g2_fill_8 FILLER_0_11_344 ();
 sg13g2_fill_8 FILLER_0_11_352 ();
 sg13g2_fill_8 FILLER_0_11_360 ();
 sg13g2_fill_8 FILLER_0_11_368 ();
 sg13g2_fill_8 FILLER_0_11_376 ();
 sg13g2_fill_8 FILLER_0_11_384 ();
 sg13g2_fill_8 FILLER_0_11_392 ();
 sg13g2_fill_8 FILLER_0_11_400 ();
 sg13g2_fill_8 FILLER_0_11_408 ();
 sg13g2_fill_8 FILLER_0_11_416 ();
 sg13g2_fill_8 FILLER_0_11_424 ();
 sg13g2_fill_8 FILLER_0_11_432 ();
 sg13g2_fill_8 FILLER_0_11_440 ();
 sg13g2_fill_8 FILLER_0_11_448 ();
 sg13g2_fill_8 FILLER_0_11_456 ();
 sg13g2_fill_8 FILLER_0_11_464 ();
 sg13g2_fill_8 FILLER_0_11_472 ();
 sg13g2_fill_8 FILLER_0_11_480 ();
 sg13g2_fill_8 FILLER_0_11_488 ();
 sg13g2_fill_8 FILLER_0_11_496 ();
 sg13g2_fill_8 FILLER_0_11_504 ();
 sg13g2_fill_8 FILLER_0_11_512 ();
 sg13g2_fill_8 FILLER_0_11_520 ();
 sg13g2_fill_8 FILLER_0_11_528 ();
 sg13g2_fill_8 FILLER_0_11_536 ();
 sg13g2_fill_8 FILLER_0_11_544 ();
 sg13g2_fill_8 FILLER_0_11_552 ();
 sg13g2_fill_8 FILLER_0_11_560 ();
 sg13g2_fill_8 FILLER_0_11_568 ();
 sg13g2_fill_8 FILLER_0_11_576 ();
 sg13g2_fill_8 FILLER_0_11_584 ();
 sg13g2_fill_8 FILLER_0_11_592 ();
 sg13g2_fill_8 FILLER_0_11_600 ();
 sg13g2_fill_8 FILLER_0_11_608 ();
 sg13g2_fill_8 FILLER_0_11_616 ();
 sg13g2_fill_8 FILLER_0_11_624 ();
 sg13g2_fill_8 FILLER_0_11_632 ();
 sg13g2_fill_8 FILLER_0_11_640 ();
 sg13g2_fill_8 FILLER_0_11_648 ();
 sg13g2_fill_8 FILLER_0_11_656 ();
 sg13g2_fill_8 FILLER_0_11_664 ();
 sg13g2_fill_8 FILLER_0_11_672 ();
 sg13g2_fill_8 FILLER_0_11_680 ();
 sg13g2_fill_8 FILLER_0_11_688 ();
 sg13g2_fill_8 FILLER_0_11_696 ();
 sg13g2_fill_8 FILLER_0_11_704 ();
 sg13g2_fill_8 FILLER_0_11_712 ();
 sg13g2_fill_8 FILLER_0_11_720 ();
 sg13g2_fill_8 FILLER_0_11_728 ();
 sg13g2_fill_8 FILLER_0_11_736 ();
 sg13g2_fill_8 FILLER_0_11_744 ();
 sg13g2_fill_8 FILLER_0_11_752 ();
 sg13g2_fill_8 FILLER_0_11_760 ();
 sg13g2_fill_8 FILLER_0_11_768 ();
 sg13g2_fill_8 FILLER_0_11_776 ();
 sg13g2_fill_8 FILLER_0_11_784 ();
 sg13g2_fill_8 FILLER_0_11_792 ();
 sg13g2_fill_8 FILLER_0_11_800 ();
 sg13g2_fill_8 FILLER_0_11_808 ();
 sg13g2_fill_8 FILLER_0_11_816 ();
 sg13g2_fill_8 FILLER_0_11_824 ();
 sg13g2_fill_8 FILLER_0_11_832 ();
 sg13g2_fill_8 FILLER_0_11_840 ();
 sg13g2_fill_8 FILLER_0_11_848 ();
 sg13g2_fill_8 FILLER_0_11_856 ();
 sg13g2_fill_8 FILLER_0_11_864 ();
 sg13g2_fill_8 FILLER_0_11_872 ();
 sg13g2_fill_8 FILLER_0_11_880 ();
 sg13g2_fill_8 FILLER_0_11_888 ();
 sg13g2_fill_8 FILLER_0_11_896 ();
 sg13g2_fill_8 FILLER_0_11_904 ();
 sg13g2_fill_8 FILLER_0_11_912 ();
 sg13g2_fill_8 FILLER_0_11_920 ();
 sg13g2_fill_8 FILLER_0_11_928 ();
 sg13g2_fill_8 FILLER_0_11_936 ();
 sg13g2_fill_8 FILLER_0_11_944 ();
 sg13g2_fill_8 FILLER_0_11_952 ();
 sg13g2_fill_8 FILLER_0_11_960 ();
 sg13g2_fill_8 FILLER_0_11_968 ();
 sg13g2_fill_8 FILLER_0_11_976 ();
 sg13g2_fill_8 FILLER_0_11_984 ();
 sg13g2_fill_8 FILLER_0_11_992 ();
 sg13g2_fill_8 FILLER_0_11_1000 ();
 sg13g2_fill_8 FILLER_0_11_1008 ();
 sg13g2_fill_8 FILLER_0_11_1016 ();
 sg13g2_fill_8 FILLER_0_11_1024 ();
 sg13g2_fill_8 FILLER_0_11_1032 ();
 sg13g2_fill_8 FILLER_0_11_1040 ();
 sg13g2_fill_8 FILLER_0_11_1048 ();
 sg13g2_fill_8 FILLER_0_11_1056 ();
 sg13g2_fill_8 FILLER_0_11_1064 ();
 sg13g2_fill_8 FILLER_0_11_1072 ();
 sg13g2_fill_8 FILLER_0_11_1080 ();
 sg13g2_fill_8 FILLER_0_11_1088 ();
 sg13g2_fill_8 FILLER_0_11_1096 ();
 sg13g2_fill_8 FILLER_0_11_1104 ();
 sg13g2_fill_8 FILLER_0_11_1112 ();
 sg13g2_fill_8 FILLER_0_11_1120 ();
 sg13g2_fill_8 FILLER_0_11_1128 ();
 sg13g2_fill_8 FILLER_0_11_1136 ();
 sg13g2_fill_8 FILLER_0_11_1144 ();
 sg13g2_fill_8 FILLER_0_11_1152 ();
 sg13g2_fill_8 FILLER_0_11_1160 ();
 sg13g2_fill_8 FILLER_0_11_1168 ();
 sg13g2_fill_8 FILLER_0_11_1176 ();
 sg13g2_fill_8 FILLER_0_11_1184 ();
 sg13g2_fill_8 FILLER_0_11_1192 ();
 sg13g2_fill_8 FILLER_0_11_1200 ();
 sg13g2_fill_8 FILLER_0_11_1208 ();
 sg13g2_fill_8 FILLER_0_11_1216 ();
 sg13g2_fill_4 FILLER_0_11_1224 ();
 sg13g2_fill_8 FILLER_0_12_0 ();
 sg13g2_fill_8 FILLER_0_12_8 ();
 sg13g2_fill_8 FILLER_0_12_16 ();
 sg13g2_fill_8 FILLER_0_12_24 ();
 sg13g2_fill_8 FILLER_0_12_32 ();
 sg13g2_fill_8 FILLER_0_12_40 ();
 sg13g2_fill_8 FILLER_0_12_48 ();
 sg13g2_fill_8 FILLER_0_12_56 ();
 sg13g2_fill_8 FILLER_0_12_64 ();
 sg13g2_fill_8 FILLER_0_12_72 ();
 sg13g2_fill_8 FILLER_0_12_80 ();
 sg13g2_fill_8 FILLER_0_12_88 ();
 sg13g2_fill_8 FILLER_0_12_96 ();
 sg13g2_fill_8 FILLER_0_12_104 ();
 sg13g2_fill_8 FILLER_0_12_112 ();
 sg13g2_fill_8 FILLER_0_12_120 ();
 sg13g2_fill_8 FILLER_0_12_128 ();
 sg13g2_fill_8 FILLER_0_12_136 ();
 sg13g2_fill_8 FILLER_0_12_144 ();
 sg13g2_fill_8 FILLER_0_12_152 ();
 sg13g2_fill_8 FILLER_0_12_160 ();
 sg13g2_fill_8 FILLER_0_12_168 ();
 sg13g2_fill_8 FILLER_0_12_176 ();
 sg13g2_fill_8 FILLER_0_12_184 ();
 sg13g2_fill_8 FILLER_0_12_192 ();
 sg13g2_fill_8 FILLER_0_12_200 ();
 sg13g2_fill_8 FILLER_0_12_208 ();
 sg13g2_fill_8 FILLER_0_12_216 ();
 sg13g2_fill_8 FILLER_0_12_224 ();
 sg13g2_fill_8 FILLER_0_12_232 ();
 sg13g2_fill_8 FILLER_0_12_240 ();
 sg13g2_fill_8 FILLER_0_12_248 ();
 sg13g2_fill_8 FILLER_0_12_256 ();
 sg13g2_fill_8 FILLER_0_12_264 ();
 sg13g2_fill_8 FILLER_0_12_272 ();
 sg13g2_fill_8 FILLER_0_12_280 ();
 sg13g2_fill_8 FILLER_0_12_288 ();
 sg13g2_fill_8 FILLER_0_12_296 ();
 sg13g2_fill_8 FILLER_0_12_304 ();
 sg13g2_fill_8 FILLER_0_12_312 ();
 sg13g2_fill_8 FILLER_0_12_320 ();
 sg13g2_fill_8 FILLER_0_12_328 ();
 sg13g2_fill_8 FILLER_0_12_336 ();
 sg13g2_fill_8 FILLER_0_12_344 ();
 sg13g2_fill_8 FILLER_0_12_352 ();
 sg13g2_fill_8 FILLER_0_12_360 ();
 sg13g2_fill_8 FILLER_0_12_368 ();
 sg13g2_fill_8 FILLER_0_12_376 ();
 sg13g2_fill_8 FILLER_0_12_384 ();
 sg13g2_fill_8 FILLER_0_12_392 ();
 sg13g2_fill_8 FILLER_0_12_400 ();
 sg13g2_fill_8 FILLER_0_12_408 ();
 sg13g2_fill_8 FILLER_0_12_416 ();
 sg13g2_fill_8 FILLER_0_12_424 ();
 sg13g2_fill_8 FILLER_0_12_432 ();
 sg13g2_fill_8 FILLER_0_12_440 ();
 sg13g2_fill_8 FILLER_0_12_448 ();
 sg13g2_fill_8 FILLER_0_12_456 ();
 sg13g2_fill_8 FILLER_0_12_464 ();
 sg13g2_fill_8 FILLER_0_12_472 ();
 sg13g2_fill_8 FILLER_0_12_480 ();
 sg13g2_fill_8 FILLER_0_12_488 ();
 sg13g2_fill_8 FILLER_0_12_496 ();
 sg13g2_fill_8 FILLER_0_12_504 ();
 sg13g2_fill_8 FILLER_0_12_512 ();
 sg13g2_fill_8 FILLER_0_12_520 ();
 sg13g2_fill_8 FILLER_0_12_528 ();
 sg13g2_fill_8 FILLER_0_12_536 ();
 sg13g2_fill_8 FILLER_0_12_544 ();
 sg13g2_fill_8 FILLER_0_12_552 ();
 sg13g2_fill_8 FILLER_0_12_560 ();
 sg13g2_fill_8 FILLER_0_12_568 ();
 sg13g2_fill_8 FILLER_0_12_576 ();
 sg13g2_fill_8 FILLER_0_12_584 ();
 sg13g2_fill_8 FILLER_0_12_592 ();
 sg13g2_fill_8 FILLER_0_12_600 ();
 sg13g2_fill_8 FILLER_0_12_608 ();
 sg13g2_fill_8 FILLER_0_12_616 ();
 sg13g2_fill_8 FILLER_0_12_624 ();
 sg13g2_fill_8 FILLER_0_12_632 ();
 sg13g2_fill_8 FILLER_0_12_640 ();
 sg13g2_fill_8 FILLER_0_12_648 ();
 sg13g2_fill_8 FILLER_0_12_656 ();
 sg13g2_fill_8 FILLER_0_12_664 ();
 sg13g2_fill_8 FILLER_0_12_672 ();
 sg13g2_fill_8 FILLER_0_12_680 ();
 sg13g2_fill_8 FILLER_0_12_688 ();
 sg13g2_fill_8 FILLER_0_12_696 ();
 sg13g2_fill_8 FILLER_0_12_704 ();
 sg13g2_fill_8 FILLER_0_12_712 ();
 sg13g2_fill_8 FILLER_0_12_720 ();
 sg13g2_fill_8 FILLER_0_12_728 ();
 sg13g2_fill_8 FILLER_0_12_736 ();
 sg13g2_fill_8 FILLER_0_12_744 ();
 sg13g2_fill_8 FILLER_0_12_752 ();
 sg13g2_fill_8 FILLER_0_12_760 ();
 sg13g2_fill_8 FILLER_0_12_768 ();
 sg13g2_fill_8 FILLER_0_12_776 ();
 sg13g2_fill_8 FILLER_0_12_784 ();
 sg13g2_fill_8 FILLER_0_12_792 ();
 sg13g2_fill_8 FILLER_0_12_800 ();
 sg13g2_fill_8 FILLER_0_12_808 ();
 sg13g2_fill_8 FILLER_0_12_816 ();
 sg13g2_fill_8 FILLER_0_12_824 ();
 sg13g2_fill_8 FILLER_0_12_832 ();
 sg13g2_fill_8 FILLER_0_12_840 ();
 sg13g2_fill_8 FILLER_0_12_848 ();
 sg13g2_fill_8 FILLER_0_12_856 ();
 sg13g2_fill_8 FILLER_0_12_864 ();
 sg13g2_fill_8 FILLER_0_12_872 ();
 sg13g2_fill_8 FILLER_0_12_880 ();
 sg13g2_fill_8 FILLER_0_12_888 ();
 sg13g2_fill_8 FILLER_0_12_896 ();
 sg13g2_fill_8 FILLER_0_12_904 ();
 sg13g2_fill_8 FILLER_0_12_912 ();
 sg13g2_fill_8 FILLER_0_12_920 ();
 sg13g2_fill_8 FILLER_0_12_928 ();
 sg13g2_fill_8 FILLER_0_12_936 ();
 sg13g2_fill_8 FILLER_0_12_944 ();
 sg13g2_fill_8 FILLER_0_12_952 ();
 sg13g2_fill_8 FILLER_0_12_960 ();
 sg13g2_fill_8 FILLER_0_12_968 ();
 sg13g2_fill_8 FILLER_0_12_976 ();
 sg13g2_fill_8 FILLER_0_12_984 ();
 sg13g2_fill_8 FILLER_0_12_992 ();
 sg13g2_fill_8 FILLER_0_12_1000 ();
 sg13g2_fill_8 FILLER_0_12_1008 ();
 sg13g2_fill_8 FILLER_0_12_1016 ();
 sg13g2_fill_8 FILLER_0_12_1024 ();
 sg13g2_fill_8 FILLER_0_12_1032 ();
 sg13g2_fill_8 FILLER_0_12_1040 ();
 sg13g2_fill_8 FILLER_0_12_1048 ();
 sg13g2_fill_8 FILLER_0_12_1056 ();
 sg13g2_fill_8 FILLER_0_12_1064 ();
 sg13g2_fill_8 FILLER_0_12_1072 ();
 sg13g2_fill_8 FILLER_0_12_1080 ();
 sg13g2_fill_8 FILLER_0_12_1088 ();
 sg13g2_fill_8 FILLER_0_12_1096 ();
 sg13g2_fill_8 FILLER_0_12_1104 ();
 sg13g2_fill_8 FILLER_0_12_1112 ();
 sg13g2_fill_8 FILLER_0_12_1120 ();
 sg13g2_fill_8 FILLER_0_12_1128 ();
 sg13g2_fill_8 FILLER_0_12_1136 ();
 sg13g2_fill_8 FILLER_0_12_1144 ();
 sg13g2_fill_8 FILLER_0_12_1152 ();
 sg13g2_fill_8 FILLER_0_12_1160 ();
 sg13g2_fill_8 FILLER_0_12_1168 ();
 sg13g2_fill_8 FILLER_0_12_1176 ();
 sg13g2_fill_8 FILLER_0_12_1184 ();
 sg13g2_fill_8 FILLER_0_12_1192 ();
 sg13g2_fill_8 FILLER_0_12_1200 ();
 sg13g2_fill_8 FILLER_0_12_1208 ();
 sg13g2_fill_8 FILLER_0_12_1216 ();
 sg13g2_fill_4 FILLER_0_12_1224 ();
 sg13g2_fill_8 FILLER_0_13_0 ();
 sg13g2_fill_8 FILLER_0_13_8 ();
 sg13g2_fill_8 FILLER_0_13_16 ();
 sg13g2_fill_8 FILLER_0_13_24 ();
 sg13g2_fill_8 FILLER_0_13_32 ();
 sg13g2_fill_8 FILLER_0_13_40 ();
 sg13g2_fill_8 FILLER_0_13_48 ();
 sg13g2_fill_8 FILLER_0_13_56 ();
 sg13g2_fill_8 FILLER_0_13_64 ();
 sg13g2_fill_8 FILLER_0_13_72 ();
 sg13g2_fill_8 FILLER_0_13_80 ();
 sg13g2_fill_8 FILLER_0_13_88 ();
 sg13g2_fill_8 FILLER_0_13_96 ();
 sg13g2_fill_8 FILLER_0_13_104 ();
 sg13g2_fill_8 FILLER_0_13_112 ();
 sg13g2_fill_8 FILLER_0_13_120 ();
 sg13g2_fill_8 FILLER_0_13_128 ();
 sg13g2_fill_8 FILLER_0_13_136 ();
 sg13g2_fill_8 FILLER_0_13_144 ();
 sg13g2_fill_8 FILLER_0_13_152 ();
 sg13g2_fill_8 FILLER_0_13_160 ();
 sg13g2_fill_8 FILLER_0_13_168 ();
 sg13g2_fill_8 FILLER_0_13_176 ();
 sg13g2_fill_8 FILLER_0_13_184 ();
 sg13g2_fill_8 FILLER_0_13_192 ();
 sg13g2_fill_8 FILLER_0_13_200 ();
 sg13g2_fill_8 FILLER_0_13_208 ();
 sg13g2_fill_8 FILLER_0_13_216 ();
 sg13g2_fill_8 FILLER_0_13_224 ();
 sg13g2_fill_8 FILLER_0_13_232 ();
 sg13g2_fill_8 FILLER_0_13_240 ();
 sg13g2_fill_8 FILLER_0_13_248 ();
 sg13g2_fill_8 FILLER_0_13_256 ();
 sg13g2_fill_8 FILLER_0_13_264 ();
 sg13g2_fill_8 FILLER_0_13_272 ();
 sg13g2_fill_8 FILLER_0_13_280 ();
 sg13g2_fill_8 FILLER_0_13_288 ();
 sg13g2_fill_8 FILLER_0_13_296 ();
 sg13g2_fill_8 FILLER_0_13_304 ();
 sg13g2_fill_8 FILLER_0_13_312 ();
 sg13g2_fill_8 FILLER_0_13_320 ();
 sg13g2_fill_8 FILLER_0_13_328 ();
 sg13g2_fill_8 FILLER_0_13_336 ();
 sg13g2_fill_8 FILLER_0_13_344 ();
 sg13g2_fill_8 FILLER_0_13_352 ();
 sg13g2_fill_8 FILLER_0_13_360 ();
 sg13g2_fill_8 FILLER_0_13_368 ();
 sg13g2_fill_8 FILLER_0_13_376 ();
 sg13g2_fill_8 FILLER_0_13_384 ();
 sg13g2_fill_8 FILLER_0_13_392 ();
 sg13g2_fill_8 FILLER_0_13_400 ();
 sg13g2_fill_8 FILLER_0_13_408 ();
 sg13g2_fill_8 FILLER_0_13_416 ();
 sg13g2_fill_8 FILLER_0_13_424 ();
 sg13g2_fill_8 FILLER_0_13_432 ();
 sg13g2_fill_8 FILLER_0_13_440 ();
 sg13g2_fill_8 FILLER_0_13_448 ();
 sg13g2_fill_8 FILLER_0_13_456 ();
 sg13g2_fill_8 FILLER_0_13_464 ();
 sg13g2_fill_8 FILLER_0_13_472 ();
 sg13g2_fill_8 FILLER_0_13_480 ();
 sg13g2_fill_8 FILLER_0_13_488 ();
 sg13g2_fill_8 FILLER_0_13_496 ();
 sg13g2_fill_8 FILLER_0_13_504 ();
 sg13g2_fill_8 FILLER_0_13_512 ();
 sg13g2_fill_8 FILLER_0_13_520 ();
 sg13g2_fill_8 FILLER_0_13_528 ();
 sg13g2_fill_8 FILLER_0_13_536 ();
 sg13g2_fill_8 FILLER_0_13_544 ();
 sg13g2_fill_8 FILLER_0_13_552 ();
 sg13g2_fill_8 FILLER_0_13_560 ();
 sg13g2_fill_8 FILLER_0_13_568 ();
 sg13g2_fill_8 FILLER_0_13_576 ();
 sg13g2_fill_8 FILLER_0_13_584 ();
 sg13g2_fill_8 FILLER_0_13_592 ();
 sg13g2_fill_8 FILLER_0_13_600 ();
 sg13g2_fill_8 FILLER_0_13_608 ();
 sg13g2_fill_8 FILLER_0_13_616 ();
 sg13g2_fill_8 FILLER_0_13_624 ();
 sg13g2_fill_8 FILLER_0_13_632 ();
 sg13g2_fill_8 FILLER_0_13_640 ();
 sg13g2_fill_8 FILLER_0_13_648 ();
 sg13g2_fill_8 FILLER_0_13_656 ();
 sg13g2_fill_8 FILLER_0_13_664 ();
 sg13g2_fill_8 FILLER_0_13_672 ();
 sg13g2_fill_8 FILLER_0_13_680 ();
 sg13g2_fill_8 FILLER_0_13_688 ();
 sg13g2_fill_8 FILLER_0_13_696 ();
 sg13g2_fill_8 FILLER_0_13_704 ();
 sg13g2_fill_8 FILLER_0_13_712 ();
 sg13g2_fill_8 FILLER_0_13_720 ();
 sg13g2_fill_8 FILLER_0_13_728 ();
 sg13g2_fill_8 FILLER_0_13_736 ();
 sg13g2_fill_8 FILLER_0_13_744 ();
 sg13g2_fill_8 FILLER_0_13_752 ();
 sg13g2_fill_8 FILLER_0_13_760 ();
 sg13g2_fill_8 FILLER_0_13_768 ();
 sg13g2_fill_8 FILLER_0_13_776 ();
 sg13g2_fill_8 FILLER_0_13_784 ();
 sg13g2_fill_8 FILLER_0_13_792 ();
 sg13g2_fill_8 FILLER_0_13_800 ();
 sg13g2_fill_8 FILLER_0_13_808 ();
 sg13g2_fill_8 FILLER_0_13_816 ();
 sg13g2_fill_8 FILLER_0_13_824 ();
 sg13g2_fill_8 FILLER_0_13_832 ();
 sg13g2_fill_8 FILLER_0_13_840 ();
 sg13g2_fill_8 FILLER_0_13_848 ();
 sg13g2_fill_8 FILLER_0_13_856 ();
 sg13g2_fill_8 FILLER_0_13_864 ();
 sg13g2_fill_8 FILLER_0_13_872 ();
 sg13g2_fill_8 FILLER_0_13_880 ();
 sg13g2_fill_8 FILLER_0_13_888 ();
 sg13g2_fill_8 FILLER_0_13_896 ();
 sg13g2_fill_8 FILLER_0_13_904 ();
 sg13g2_fill_8 FILLER_0_13_912 ();
 sg13g2_fill_8 FILLER_0_13_920 ();
 sg13g2_fill_8 FILLER_0_13_928 ();
 sg13g2_fill_8 FILLER_0_13_936 ();
 sg13g2_fill_8 FILLER_0_13_944 ();
 sg13g2_fill_8 FILLER_0_13_952 ();
 sg13g2_fill_8 FILLER_0_13_960 ();
 sg13g2_fill_8 FILLER_0_13_968 ();
 sg13g2_fill_8 FILLER_0_13_976 ();
 sg13g2_fill_8 FILLER_0_13_984 ();
 sg13g2_fill_8 FILLER_0_13_992 ();
 sg13g2_fill_8 FILLER_0_13_1000 ();
 sg13g2_fill_8 FILLER_0_13_1008 ();
 sg13g2_fill_8 FILLER_0_13_1016 ();
 sg13g2_fill_8 FILLER_0_13_1024 ();
 sg13g2_fill_8 FILLER_0_13_1032 ();
 sg13g2_fill_8 FILLER_0_13_1040 ();
 sg13g2_fill_8 FILLER_0_13_1048 ();
 sg13g2_fill_8 FILLER_0_13_1056 ();
 sg13g2_fill_8 FILLER_0_13_1064 ();
 sg13g2_fill_8 FILLER_0_13_1072 ();
 sg13g2_fill_8 FILLER_0_13_1080 ();
 sg13g2_fill_8 FILLER_0_13_1088 ();
 sg13g2_fill_8 FILLER_0_13_1096 ();
 sg13g2_fill_8 FILLER_0_13_1104 ();
 sg13g2_fill_8 FILLER_0_13_1112 ();
 sg13g2_fill_8 FILLER_0_13_1120 ();
 sg13g2_fill_8 FILLER_0_13_1128 ();
 sg13g2_fill_8 FILLER_0_13_1136 ();
 sg13g2_fill_8 FILLER_0_13_1144 ();
 sg13g2_fill_8 FILLER_0_13_1152 ();
 sg13g2_fill_8 FILLER_0_13_1160 ();
 sg13g2_fill_8 FILLER_0_13_1168 ();
 sg13g2_fill_8 FILLER_0_13_1176 ();
 sg13g2_fill_8 FILLER_0_13_1184 ();
 sg13g2_fill_8 FILLER_0_13_1192 ();
 sg13g2_fill_8 FILLER_0_13_1200 ();
 sg13g2_fill_8 FILLER_0_13_1208 ();
 sg13g2_fill_8 FILLER_0_13_1216 ();
 sg13g2_fill_4 FILLER_0_13_1224 ();
 sg13g2_fill_8 FILLER_0_14_0 ();
 sg13g2_fill_8 FILLER_0_14_8 ();
 sg13g2_fill_8 FILLER_0_14_16 ();
 sg13g2_fill_8 FILLER_0_14_24 ();
 sg13g2_fill_8 FILLER_0_14_32 ();
 sg13g2_fill_8 FILLER_0_14_40 ();
 sg13g2_fill_8 FILLER_0_14_48 ();
 sg13g2_fill_8 FILLER_0_14_56 ();
 sg13g2_fill_8 FILLER_0_14_64 ();
 sg13g2_fill_8 FILLER_0_14_72 ();
 sg13g2_fill_8 FILLER_0_14_80 ();
 sg13g2_fill_8 FILLER_0_14_88 ();
 sg13g2_fill_8 FILLER_0_14_96 ();
 sg13g2_fill_8 FILLER_0_14_104 ();
 sg13g2_fill_8 FILLER_0_14_112 ();
 sg13g2_fill_8 FILLER_0_14_120 ();
 sg13g2_fill_8 FILLER_0_14_128 ();
 sg13g2_fill_8 FILLER_0_14_136 ();
 sg13g2_fill_8 FILLER_0_14_144 ();
 sg13g2_fill_8 FILLER_0_14_152 ();
 sg13g2_fill_8 FILLER_0_14_160 ();
 sg13g2_fill_8 FILLER_0_14_168 ();
 sg13g2_fill_8 FILLER_0_14_176 ();
 sg13g2_fill_8 FILLER_0_14_184 ();
 sg13g2_fill_8 FILLER_0_14_192 ();
 sg13g2_fill_8 FILLER_0_14_200 ();
 sg13g2_fill_8 FILLER_0_14_208 ();
 sg13g2_fill_8 FILLER_0_14_216 ();
 sg13g2_fill_8 FILLER_0_14_224 ();
 sg13g2_fill_8 FILLER_0_14_232 ();
 sg13g2_fill_8 FILLER_0_14_240 ();
 sg13g2_fill_8 FILLER_0_14_248 ();
 sg13g2_fill_8 FILLER_0_14_256 ();
 sg13g2_fill_8 FILLER_0_14_264 ();
 sg13g2_fill_8 FILLER_0_14_272 ();
 sg13g2_fill_8 FILLER_0_14_280 ();
 sg13g2_fill_8 FILLER_0_14_288 ();
 sg13g2_fill_8 FILLER_0_14_296 ();
 sg13g2_fill_8 FILLER_0_14_304 ();
 sg13g2_fill_8 FILLER_0_14_312 ();
 sg13g2_fill_8 FILLER_0_14_320 ();
 sg13g2_fill_8 FILLER_0_14_328 ();
 sg13g2_fill_8 FILLER_0_14_336 ();
 sg13g2_fill_8 FILLER_0_14_344 ();
 sg13g2_fill_8 FILLER_0_14_352 ();
 sg13g2_fill_8 FILLER_0_14_360 ();
 sg13g2_fill_8 FILLER_0_14_368 ();
 sg13g2_fill_8 FILLER_0_14_376 ();
 sg13g2_fill_8 FILLER_0_14_384 ();
 sg13g2_fill_8 FILLER_0_14_392 ();
 sg13g2_fill_8 FILLER_0_14_400 ();
 sg13g2_fill_8 FILLER_0_14_408 ();
 sg13g2_fill_8 FILLER_0_14_416 ();
 sg13g2_fill_8 FILLER_0_14_424 ();
 sg13g2_fill_8 FILLER_0_14_432 ();
 sg13g2_fill_8 FILLER_0_14_440 ();
 sg13g2_fill_8 FILLER_0_14_448 ();
 sg13g2_fill_8 FILLER_0_14_456 ();
 sg13g2_fill_8 FILLER_0_14_464 ();
 sg13g2_fill_8 FILLER_0_14_472 ();
 sg13g2_fill_8 FILLER_0_14_480 ();
 sg13g2_fill_8 FILLER_0_14_488 ();
 sg13g2_fill_8 FILLER_0_14_496 ();
 sg13g2_fill_8 FILLER_0_14_504 ();
 sg13g2_fill_8 FILLER_0_14_512 ();
 sg13g2_fill_8 FILLER_0_14_520 ();
 sg13g2_fill_8 FILLER_0_14_528 ();
 sg13g2_fill_8 FILLER_0_14_536 ();
 sg13g2_fill_8 FILLER_0_14_544 ();
 sg13g2_fill_8 FILLER_0_14_552 ();
 sg13g2_fill_8 FILLER_0_14_560 ();
 sg13g2_fill_8 FILLER_0_14_568 ();
 sg13g2_fill_8 FILLER_0_14_576 ();
 sg13g2_fill_8 FILLER_0_14_584 ();
 sg13g2_fill_8 FILLER_0_14_592 ();
 sg13g2_fill_8 FILLER_0_14_600 ();
 sg13g2_fill_8 FILLER_0_14_608 ();
 sg13g2_fill_8 FILLER_0_14_616 ();
 sg13g2_fill_8 FILLER_0_14_624 ();
 sg13g2_fill_8 FILLER_0_14_632 ();
 sg13g2_fill_8 FILLER_0_14_640 ();
 sg13g2_fill_8 FILLER_0_14_648 ();
 sg13g2_fill_8 FILLER_0_14_656 ();
 sg13g2_fill_8 FILLER_0_14_664 ();
 sg13g2_fill_8 FILLER_0_14_672 ();
 sg13g2_fill_8 FILLER_0_14_680 ();
 sg13g2_fill_8 FILLER_0_14_688 ();
 sg13g2_fill_8 FILLER_0_14_696 ();
 sg13g2_fill_8 FILLER_0_14_704 ();
 sg13g2_fill_8 FILLER_0_14_712 ();
 sg13g2_fill_8 FILLER_0_14_720 ();
 sg13g2_fill_8 FILLER_0_14_728 ();
 sg13g2_fill_8 FILLER_0_14_736 ();
 sg13g2_fill_8 FILLER_0_14_744 ();
 sg13g2_fill_8 FILLER_0_14_752 ();
 sg13g2_fill_8 FILLER_0_14_760 ();
 sg13g2_fill_8 FILLER_0_14_768 ();
 sg13g2_fill_8 FILLER_0_14_776 ();
 sg13g2_fill_8 FILLER_0_14_784 ();
 sg13g2_fill_8 FILLER_0_14_792 ();
 sg13g2_fill_8 FILLER_0_14_800 ();
 sg13g2_fill_8 FILLER_0_14_808 ();
 sg13g2_fill_8 FILLER_0_14_816 ();
 sg13g2_fill_8 FILLER_0_14_824 ();
 sg13g2_fill_8 FILLER_0_14_832 ();
 sg13g2_fill_8 FILLER_0_14_840 ();
 sg13g2_fill_8 FILLER_0_14_848 ();
 sg13g2_fill_8 FILLER_0_14_856 ();
 sg13g2_fill_8 FILLER_0_14_864 ();
 sg13g2_fill_8 FILLER_0_14_872 ();
 sg13g2_fill_8 FILLER_0_14_880 ();
 sg13g2_fill_8 FILLER_0_14_888 ();
 sg13g2_fill_8 FILLER_0_14_896 ();
 sg13g2_fill_8 FILLER_0_14_904 ();
 sg13g2_fill_8 FILLER_0_14_912 ();
 sg13g2_fill_8 FILLER_0_14_920 ();
 sg13g2_fill_8 FILLER_0_14_928 ();
 sg13g2_fill_8 FILLER_0_14_936 ();
 sg13g2_fill_8 FILLER_0_14_944 ();
 sg13g2_fill_8 FILLER_0_14_952 ();
 sg13g2_fill_8 FILLER_0_14_960 ();
 sg13g2_fill_8 FILLER_0_14_968 ();
 sg13g2_fill_8 FILLER_0_14_976 ();
 sg13g2_fill_8 FILLER_0_14_984 ();
 sg13g2_fill_8 FILLER_0_14_992 ();
 sg13g2_fill_8 FILLER_0_14_1000 ();
 sg13g2_fill_8 FILLER_0_14_1008 ();
 sg13g2_fill_8 FILLER_0_14_1016 ();
 sg13g2_fill_8 FILLER_0_14_1024 ();
 sg13g2_fill_8 FILLER_0_14_1032 ();
 sg13g2_fill_8 FILLER_0_14_1040 ();
 sg13g2_fill_8 FILLER_0_14_1048 ();
 sg13g2_fill_8 FILLER_0_14_1056 ();
 sg13g2_fill_8 FILLER_0_14_1064 ();
 sg13g2_fill_8 FILLER_0_14_1072 ();
 sg13g2_fill_8 FILLER_0_14_1080 ();
 sg13g2_fill_8 FILLER_0_14_1088 ();
 sg13g2_fill_8 FILLER_0_14_1096 ();
 sg13g2_fill_8 FILLER_0_14_1104 ();
 sg13g2_fill_8 FILLER_0_14_1112 ();
 sg13g2_fill_8 FILLER_0_14_1120 ();
 sg13g2_fill_8 FILLER_0_14_1128 ();
 sg13g2_fill_8 FILLER_0_14_1136 ();
 sg13g2_fill_8 FILLER_0_14_1144 ();
 sg13g2_fill_8 FILLER_0_14_1152 ();
 sg13g2_fill_8 FILLER_0_14_1160 ();
 sg13g2_fill_8 FILLER_0_14_1168 ();
 sg13g2_fill_8 FILLER_0_14_1176 ();
 sg13g2_fill_8 FILLER_0_14_1184 ();
 sg13g2_fill_8 FILLER_0_14_1192 ();
 sg13g2_fill_8 FILLER_0_14_1200 ();
 sg13g2_fill_8 FILLER_0_14_1208 ();
 sg13g2_fill_8 FILLER_0_14_1216 ();
 sg13g2_fill_4 FILLER_0_14_1224 ();
 sg13g2_fill_8 FILLER_0_15_0 ();
 sg13g2_fill_8 FILLER_0_15_8 ();
 sg13g2_fill_8 FILLER_0_15_16 ();
 sg13g2_fill_8 FILLER_0_15_24 ();
 sg13g2_fill_8 FILLER_0_15_32 ();
 sg13g2_fill_8 FILLER_0_15_40 ();
 sg13g2_fill_8 FILLER_0_15_48 ();
 sg13g2_fill_8 FILLER_0_15_56 ();
 sg13g2_fill_8 FILLER_0_15_64 ();
 sg13g2_fill_8 FILLER_0_15_72 ();
 sg13g2_fill_8 FILLER_0_15_80 ();
 sg13g2_fill_8 FILLER_0_15_88 ();
 sg13g2_fill_8 FILLER_0_15_96 ();
 sg13g2_fill_8 FILLER_0_15_104 ();
 sg13g2_fill_8 FILLER_0_15_112 ();
 sg13g2_fill_8 FILLER_0_15_120 ();
 sg13g2_fill_8 FILLER_0_15_128 ();
 sg13g2_fill_8 FILLER_0_15_136 ();
 sg13g2_fill_8 FILLER_0_15_144 ();
 sg13g2_fill_8 FILLER_0_15_152 ();
 sg13g2_fill_8 FILLER_0_15_160 ();
 sg13g2_fill_8 FILLER_0_15_168 ();
 sg13g2_fill_8 FILLER_0_15_176 ();
 sg13g2_fill_8 FILLER_0_15_184 ();
 sg13g2_fill_8 FILLER_0_15_192 ();
 sg13g2_fill_8 FILLER_0_15_200 ();
 sg13g2_fill_8 FILLER_0_15_208 ();
 sg13g2_fill_8 FILLER_0_15_216 ();
 sg13g2_fill_8 FILLER_0_15_224 ();
 sg13g2_fill_8 FILLER_0_15_232 ();
 sg13g2_fill_8 FILLER_0_15_240 ();
 sg13g2_fill_8 FILLER_0_15_248 ();
 sg13g2_fill_8 FILLER_0_15_256 ();
 sg13g2_fill_8 FILLER_0_15_264 ();
 sg13g2_fill_8 FILLER_0_15_272 ();
 sg13g2_fill_8 FILLER_0_15_280 ();
 sg13g2_fill_8 FILLER_0_15_288 ();
 sg13g2_fill_8 FILLER_0_15_296 ();
 sg13g2_fill_8 FILLER_0_15_304 ();
 sg13g2_fill_8 FILLER_0_15_312 ();
 sg13g2_fill_8 FILLER_0_15_320 ();
 sg13g2_fill_8 FILLER_0_15_328 ();
 sg13g2_fill_8 FILLER_0_15_336 ();
 sg13g2_fill_8 FILLER_0_15_344 ();
 sg13g2_fill_8 FILLER_0_15_352 ();
 sg13g2_fill_8 FILLER_0_15_360 ();
 sg13g2_fill_8 FILLER_0_15_368 ();
 sg13g2_fill_8 FILLER_0_15_376 ();
 sg13g2_fill_8 FILLER_0_15_384 ();
 sg13g2_fill_8 FILLER_0_15_392 ();
 sg13g2_fill_8 FILLER_0_15_400 ();
 sg13g2_fill_8 FILLER_0_15_408 ();
 sg13g2_fill_8 FILLER_0_15_416 ();
 sg13g2_fill_8 FILLER_0_15_424 ();
 sg13g2_fill_8 FILLER_0_15_432 ();
 sg13g2_fill_8 FILLER_0_15_440 ();
 sg13g2_fill_8 FILLER_0_15_448 ();
 sg13g2_fill_8 FILLER_0_15_456 ();
 sg13g2_fill_8 FILLER_0_15_464 ();
 sg13g2_fill_8 FILLER_0_15_472 ();
 sg13g2_fill_8 FILLER_0_15_480 ();
 sg13g2_fill_8 FILLER_0_15_488 ();
 sg13g2_fill_8 FILLER_0_15_496 ();
 sg13g2_fill_8 FILLER_0_15_504 ();
 sg13g2_fill_8 FILLER_0_15_512 ();
 sg13g2_fill_8 FILLER_0_15_520 ();
 sg13g2_fill_8 FILLER_0_15_528 ();
 sg13g2_fill_8 FILLER_0_15_536 ();
 sg13g2_fill_8 FILLER_0_15_544 ();
 sg13g2_fill_8 FILLER_0_15_552 ();
 sg13g2_fill_8 FILLER_0_15_560 ();
 sg13g2_fill_8 FILLER_0_15_568 ();
 sg13g2_fill_8 FILLER_0_15_576 ();
 sg13g2_fill_8 FILLER_0_15_584 ();
 sg13g2_fill_8 FILLER_0_15_592 ();
 sg13g2_fill_8 FILLER_0_15_600 ();
 sg13g2_fill_8 FILLER_0_15_608 ();
 sg13g2_fill_8 FILLER_0_15_616 ();
 sg13g2_fill_8 FILLER_0_15_624 ();
 sg13g2_fill_8 FILLER_0_15_632 ();
 sg13g2_fill_8 FILLER_0_15_640 ();
 sg13g2_fill_8 FILLER_0_15_648 ();
 sg13g2_fill_8 FILLER_0_15_656 ();
 sg13g2_fill_8 FILLER_0_15_664 ();
 sg13g2_fill_8 FILLER_0_15_672 ();
 sg13g2_fill_8 FILLER_0_15_680 ();
 sg13g2_fill_8 FILLER_0_15_688 ();
 sg13g2_fill_8 FILLER_0_15_696 ();
 sg13g2_fill_8 FILLER_0_15_704 ();
 sg13g2_fill_8 FILLER_0_15_712 ();
 sg13g2_fill_8 FILLER_0_15_720 ();
 sg13g2_fill_8 FILLER_0_15_728 ();
 sg13g2_fill_8 FILLER_0_15_736 ();
 sg13g2_fill_8 FILLER_0_15_744 ();
 sg13g2_fill_8 FILLER_0_15_752 ();
 sg13g2_fill_8 FILLER_0_15_760 ();
 sg13g2_fill_8 FILLER_0_15_768 ();
 sg13g2_fill_8 FILLER_0_15_776 ();
 sg13g2_fill_8 FILLER_0_15_784 ();
 sg13g2_fill_8 FILLER_0_15_792 ();
 sg13g2_fill_8 FILLER_0_15_800 ();
 sg13g2_fill_8 FILLER_0_15_808 ();
 sg13g2_fill_8 FILLER_0_15_816 ();
 sg13g2_fill_8 FILLER_0_15_824 ();
 sg13g2_fill_8 FILLER_0_15_832 ();
 sg13g2_fill_8 FILLER_0_15_840 ();
 sg13g2_fill_8 FILLER_0_15_848 ();
 sg13g2_fill_8 FILLER_0_15_856 ();
 sg13g2_fill_8 FILLER_0_15_864 ();
 sg13g2_fill_8 FILLER_0_15_872 ();
 sg13g2_fill_8 FILLER_0_15_880 ();
 sg13g2_fill_8 FILLER_0_15_888 ();
 sg13g2_fill_8 FILLER_0_15_896 ();
 sg13g2_fill_8 FILLER_0_15_904 ();
 sg13g2_fill_8 FILLER_0_15_912 ();
 sg13g2_fill_8 FILLER_0_15_920 ();
 sg13g2_fill_8 FILLER_0_15_928 ();
 sg13g2_fill_8 FILLER_0_15_936 ();
 sg13g2_fill_8 FILLER_0_15_944 ();
 sg13g2_fill_8 FILLER_0_15_952 ();
 sg13g2_fill_8 FILLER_0_15_960 ();
 sg13g2_fill_8 FILLER_0_15_968 ();
 sg13g2_fill_8 FILLER_0_15_976 ();
 sg13g2_fill_8 FILLER_0_15_984 ();
 sg13g2_fill_8 FILLER_0_15_992 ();
 sg13g2_fill_8 FILLER_0_15_1000 ();
 sg13g2_fill_8 FILLER_0_15_1008 ();
 sg13g2_fill_8 FILLER_0_15_1016 ();
 sg13g2_fill_8 FILLER_0_15_1024 ();
 sg13g2_fill_8 FILLER_0_15_1032 ();
 sg13g2_fill_8 FILLER_0_15_1040 ();
 sg13g2_fill_8 FILLER_0_15_1048 ();
 sg13g2_fill_8 FILLER_0_15_1056 ();
 sg13g2_fill_8 FILLER_0_15_1064 ();
 sg13g2_fill_8 FILLER_0_15_1072 ();
 sg13g2_fill_8 FILLER_0_15_1080 ();
 sg13g2_fill_8 FILLER_0_15_1088 ();
 sg13g2_fill_8 FILLER_0_15_1096 ();
 sg13g2_fill_8 FILLER_0_15_1104 ();
 sg13g2_fill_8 FILLER_0_15_1112 ();
 sg13g2_fill_8 FILLER_0_15_1120 ();
 sg13g2_fill_8 FILLER_0_15_1128 ();
 sg13g2_fill_8 FILLER_0_15_1136 ();
 sg13g2_fill_8 FILLER_0_15_1144 ();
 sg13g2_fill_8 FILLER_0_15_1152 ();
 sg13g2_fill_8 FILLER_0_15_1160 ();
 sg13g2_fill_8 FILLER_0_15_1168 ();
 sg13g2_fill_8 FILLER_0_15_1176 ();
 sg13g2_fill_8 FILLER_0_15_1184 ();
 sg13g2_fill_8 FILLER_0_15_1192 ();
 sg13g2_fill_8 FILLER_0_15_1200 ();
 sg13g2_fill_8 FILLER_0_15_1208 ();
 sg13g2_fill_8 FILLER_0_15_1216 ();
 sg13g2_fill_4 FILLER_0_15_1224 ();
 sg13g2_fill_8 FILLER_0_16_0 ();
 sg13g2_fill_8 FILLER_0_16_8 ();
 sg13g2_fill_8 FILLER_0_16_16 ();
 sg13g2_fill_8 FILLER_0_16_24 ();
 sg13g2_fill_8 FILLER_0_16_32 ();
 sg13g2_fill_8 FILLER_0_16_40 ();
 sg13g2_fill_8 FILLER_0_16_48 ();
 sg13g2_fill_8 FILLER_0_16_56 ();
 sg13g2_fill_8 FILLER_0_16_64 ();
 sg13g2_fill_8 FILLER_0_16_72 ();
 sg13g2_fill_8 FILLER_0_16_80 ();
 sg13g2_fill_8 FILLER_0_16_88 ();
 sg13g2_fill_8 FILLER_0_16_96 ();
 sg13g2_fill_8 FILLER_0_16_104 ();
 sg13g2_fill_8 FILLER_0_16_112 ();
 sg13g2_fill_8 FILLER_0_16_120 ();
 sg13g2_fill_8 FILLER_0_16_128 ();
 sg13g2_fill_8 FILLER_0_16_136 ();
 sg13g2_fill_8 FILLER_0_16_144 ();
 sg13g2_fill_8 FILLER_0_16_152 ();
 sg13g2_fill_8 FILLER_0_16_160 ();
 sg13g2_fill_8 FILLER_0_16_168 ();
 sg13g2_fill_8 FILLER_0_16_176 ();
 sg13g2_fill_8 FILLER_0_16_184 ();
 sg13g2_fill_8 FILLER_0_16_192 ();
 sg13g2_fill_8 FILLER_0_16_200 ();
 sg13g2_fill_8 FILLER_0_16_208 ();
 sg13g2_fill_8 FILLER_0_16_216 ();
 sg13g2_fill_8 FILLER_0_16_224 ();
 sg13g2_fill_8 FILLER_0_16_232 ();
 sg13g2_fill_8 FILLER_0_16_240 ();
 sg13g2_fill_8 FILLER_0_16_248 ();
 sg13g2_fill_8 FILLER_0_16_256 ();
 sg13g2_fill_8 FILLER_0_16_264 ();
 sg13g2_fill_8 FILLER_0_16_272 ();
 sg13g2_fill_8 FILLER_0_16_280 ();
 sg13g2_fill_8 FILLER_0_16_288 ();
 sg13g2_fill_8 FILLER_0_16_296 ();
 sg13g2_fill_8 FILLER_0_16_304 ();
 sg13g2_fill_8 FILLER_0_16_312 ();
 sg13g2_fill_8 FILLER_0_16_320 ();
 sg13g2_fill_8 FILLER_0_16_328 ();
 sg13g2_fill_8 FILLER_0_16_336 ();
 sg13g2_fill_8 FILLER_0_16_344 ();
 sg13g2_fill_8 FILLER_0_16_352 ();
 sg13g2_fill_8 FILLER_0_16_360 ();
 sg13g2_fill_8 FILLER_0_16_368 ();
 sg13g2_fill_8 FILLER_0_16_376 ();
 sg13g2_fill_8 FILLER_0_16_384 ();
 sg13g2_fill_8 FILLER_0_16_392 ();
 sg13g2_fill_8 FILLER_0_16_400 ();
 sg13g2_fill_8 FILLER_0_16_408 ();
 sg13g2_fill_8 FILLER_0_16_416 ();
 sg13g2_fill_8 FILLER_0_16_424 ();
 sg13g2_fill_8 FILLER_0_16_432 ();
 sg13g2_fill_8 FILLER_0_16_440 ();
 sg13g2_fill_8 FILLER_0_16_448 ();
 sg13g2_fill_8 FILLER_0_16_456 ();
 sg13g2_fill_8 FILLER_0_16_464 ();
 sg13g2_fill_8 FILLER_0_16_472 ();
 sg13g2_fill_8 FILLER_0_16_480 ();
 sg13g2_fill_8 FILLER_0_16_488 ();
 sg13g2_fill_8 FILLER_0_16_496 ();
 sg13g2_fill_8 FILLER_0_16_504 ();
 sg13g2_fill_8 FILLER_0_16_512 ();
 sg13g2_fill_8 FILLER_0_16_520 ();
 sg13g2_fill_8 FILLER_0_16_528 ();
 sg13g2_fill_8 FILLER_0_16_536 ();
 sg13g2_fill_8 FILLER_0_16_544 ();
 sg13g2_fill_8 FILLER_0_16_552 ();
 sg13g2_fill_8 FILLER_0_16_560 ();
 sg13g2_fill_8 FILLER_0_16_568 ();
 sg13g2_fill_8 FILLER_0_16_576 ();
 sg13g2_fill_8 FILLER_0_16_584 ();
 sg13g2_fill_8 FILLER_0_16_592 ();
 sg13g2_fill_8 FILLER_0_16_600 ();
 sg13g2_fill_8 FILLER_0_16_608 ();
 sg13g2_fill_8 FILLER_0_16_616 ();
 sg13g2_fill_8 FILLER_0_16_624 ();
 sg13g2_fill_8 FILLER_0_16_632 ();
 sg13g2_fill_8 FILLER_0_16_640 ();
 sg13g2_fill_8 FILLER_0_16_648 ();
 sg13g2_fill_8 FILLER_0_16_656 ();
 sg13g2_fill_8 FILLER_0_16_664 ();
 sg13g2_fill_8 FILLER_0_16_672 ();
 sg13g2_fill_8 FILLER_0_16_680 ();
 sg13g2_fill_8 FILLER_0_16_688 ();
 sg13g2_fill_8 FILLER_0_16_696 ();
 sg13g2_fill_8 FILLER_0_16_704 ();
 sg13g2_fill_8 FILLER_0_16_712 ();
 sg13g2_fill_8 FILLER_0_16_720 ();
 sg13g2_fill_8 FILLER_0_16_728 ();
 sg13g2_fill_8 FILLER_0_16_736 ();
 sg13g2_fill_8 FILLER_0_16_744 ();
 sg13g2_fill_8 FILLER_0_16_752 ();
 sg13g2_fill_8 FILLER_0_16_760 ();
 sg13g2_fill_8 FILLER_0_16_768 ();
 sg13g2_fill_8 FILLER_0_16_776 ();
 sg13g2_fill_8 FILLER_0_16_784 ();
 sg13g2_fill_8 FILLER_0_16_792 ();
 sg13g2_fill_8 FILLER_0_16_800 ();
 sg13g2_fill_8 FILLER_0_16_808 ();
 sg13g2_fill_8 FILLER_0_16_816 ();
 sg13g2_fill_8 FILLER_0_16_824 ();
 sg13g2_fill_8 FILLER_0_16_832 ();
 sg13g2_fill_8 FILLER_0_16_840 ();
 sg13g2_fill_8 FILLER_0_16_848 ();
 sg13g2_fill_8 FILLER_0_16_856 ();
 sg13g2_fill_8 FILLER_0_16_864 ();
 sg13g2_fill_8 FILLER_0_16_872 ();
 sg13g2_fill_8 FILLER_0_16_880 ();
 sg13g2_fill_8 FILLER_0_16_888 ();
 sg13g2_fill_8 FILLER_0_16_896 ();
 sg13g2_fill_8 FILLER_0_16_904 ();
 sg13g2_fill_8 FILLER_0_16_912 ();
 sg13g2_fill_8 FILLER_0_16_920 ();
 sg13g2_fill_8 FILLER_0_16_928 ();
 sg13g2_fill_8 FILLER_0_16_936 ();
 sg13g2_fill_8 FILLER_0_16_944 ();
 sg13g2_fill_8 FILLER_0_16_952 ();
 sg13g2_fill_8 FILLER_0_16_960 ();
 sg13g2_fill_8 FILLER_0_16_968 ();
 sg13g2_fill_8 FILLER_0_16_976 ();
 sg13g2_fill_8 FILLER_0_16_984 ();
 sg13g2_fill_8 FILLER_0_16_992 ();
 sg13g2_fill_8 FILLER_0_16_1000 ();
 sg13g2_fill_8 FILLER_0_16_1008 ();
 sg13g2_fill_8 FILLER_0_16_1016 ();
 sg13g2_fill_8 FILLER_0_16_1024 ();
 sg13g2_fill_8 FILLER_0_16_1032 ();
 sg13g2_fill_8 FILLER_0_16_1040 ();
 sg13g2_fill_8 FILLER_0_16_1048 ();
 sg13g2_fill_8 FILLER_0_16_1056 ();
 sg13g2_fill_8 FILLER_0_16_1064 ();
 sg13g2_fill_8 FILLER_0_16_1072 ();
 sg13g2_fill_8 FILLER_0_16_1080 ();
 sg13g2_fill_8 FILLER_0_16_1088 ();
 sg13g2_fill_8 FILLER_0_16_1096 ();
 sg13g2_fill_8 FILLER_0_16_1104 ();
 sg13g2_fill_8 FILLER_0_16_1112 ();
 sg13g2_fill_8 FILLER_0_16_1120 ();
 sg13g2_fill_8 FILLER_0_16_1128 ();
 sg13g2_fill_8 FILLER_0_16_1136 ();
 sg13g2_fill_8 FILLER_0_16_1144 ();
 sg13g2_fill_8 FILLER_0_16_1152 ();
 sg13g2_fill_8 FILLER_0_16_1160 ();
 sg13g2_fill_8 FILLER_0_16_1168 ();
 sg13g2_fill_8 FILLER_0_16_1176 ();
 sg13g2_fill_8 FILLER_0_16_1184 ();
 sg13g2_fill_8 FILLER_0_16_1192 ();
 sg13g2_fill_8 FILLER_0_16_1200 ();
 sg13g2_fill_8 FILLER_0_16_1208 ();
 sg13g2_fill_8 FILLER_0_16_1216 ();
 sg13g2_fill_4 FILLER_0_16_1224 ();
 sg13g2_fill_8 FILLER_0_17_0 ();
 sg13g2_fill_8 FILLER_0_17_8 ();
 sg13g2_fill_8 FILLER_0_17_16 ();
 sg13g2_fill_8 FILLER_0_17_24 ();
 sg13g2_fill_8 FILLER_0_17_32 ();
 sg13g2_fill_8 FILLER_0_17_40 ();
 sg13g2_fill_8 FILLER_0_17_48 ();
 sg13g2_fill_8 FILLER_0_17_56 ();
 sg13g2_fill_8 FILLER_0_17_64 ();
 sg13g2_fill_8 FILLER_0_17_72 ();
 sg13g2_fill_8 FILLER_0_17_80 ();
 sg13g2_fill_8 FILLER_0_17_88 ();
 sg13g2_fill_8 FILLER_0_17_96 ();
 sg13g2_fill_8 FILLER_0_17_104 ();
 sg13g2_fill_8 FILLER_0_17_112 ();
 sg13g2_fill_8 FILLER_0_17_120 ();
 sg13g2_fill_8 FILLER_0_17_128 ();
 sg13g2_fill_8 FILLER_0_17_136 ();
 sg13g2_fill_8 FILLER_0_17_144 ();
 sg13g2_fill_8 FILLER_0_17_152 ();
 sg13g2_fill_8 FILLER_0_17_160 ();
 sg13g2_fill_8 FILLER_0_17_168 ();
 sg13g2_fill_8 FILLER_0_17_176 ();
 sg13g2_fill_8 FILLER_0_17_184 ();
 sg13g2_fill_8 FILLER_0_17_192 ();
 sg13g2_fill_8 FILLER_0_17_200 ();
 sg13g2_fill_8 FILLER_0_17_208 ();
 sg13g2_fill_8 FILLER_0_17_216 ();
 sg13g2_fill_8 FILLER_0_17_224 ();
 sg13g2_fill_8 FILLER_0_17_232 ();
 sg13g2_fill_8 FILLER_0_17_240 ();
 sg13g2_fill_8 FILLER_0_17_248 ();
 sg13g2_fill_8 FILLER_0_17_256 ();
 sg13g2_fill_8 FILLER_0_17_264 ();
 sg13g2_fill_8 FILLER_0_17_272 ();
 sg13g2_fill_8 FILLER_0_17_280 ();
 sg13g2_fill_8 FILLER_0_17_288 ();
 sg13g2_fill_8 FILLER_0_17_296 ();
 sg13g2_fill_8 FILLER_0_17_304 ();
 sg13g2_fill_8 FILLER_0_17_312 ();
 sg13g2_fill_8 FILLER_0_17_320 ();
 sg13g2_fill_8 FILLER_0_17_328 ();
 sg13g2_fill_8 FILLER_0_17_336 ();
 sg13g2_fill_8 FILLER_0_17_344 ();
 sg13g2_fill_8 FILLER_0_17_352 ();
 sg13g2_fill_8 FILLER_0_17_360 ();
 sg13g2_fill_8 FILLER_0_17_368 ();
 sg13g2_fill_8 FILLER_0_17_376 ();
 sg13g2_fill_8 FILLER_0_17_384 ();
 sg13g2_fill_8 FILLER_0_17_392 ();
 sg13g2_fill_8 FILLER_0_17_400 ();
 sg13g2_fill_8 FILLER_0_17_408 ();
 sg13g2_fill_8 FILLER_0_17_416 ();
 sg13g2_fill_8 FILLER_0_17_424 ();
 sg13g2_fill_8 FILLER_0_17_432 ();
 sg13g2_fill_8 FILLER_0_17_440 ();
 sg13g2_fill_8 FILLER_0_17_448 ();
 sg13g2_fill_8 FILLER_0_17_456 ();
 sg13g2_fill_8 FILLER_0_17_464 ();
 sg13g2_fill_8 FILLER_0_17_472 ();
 sg13g2_fill_8 FILLER_0_17_480 ();
 sg13g2_fill_8 FILLER_0_17_488 ();
 sg13g2_fill_8 FILLER_0_17_496 ();
 sg13g2_fill_8 FILLER_0_17_504 ();
 sg13g2_fill_8 FILLER_0_17_512 ();
 sg13g2_fill_8 FILLER_0_17_520 ();
 sg13g2_fill_8 FILLER_0_17_528 ();
 sg13g2_fill_8 FILLER_0_17_536 ();
 sg13g2_fill_8 FILLER_0_17_544 ();
 sg13g2_fill_8 FILLER_0_17_552 ();
 sg13g2_fill_8 FILLER_0_17_560 ();
 sg13g2_fill_8 FILLER_0_17_568 ();
 sg13g2_fill_8 FILLER_0_17_576 ();
 sg13g2_fill_8 FILLER_0_17_584 ();
 sg13g2_fill_8 FILLER_0_17_592 ();
 sg13g2_fill_8 FILLER_0_17_600 ();
 sg13g2_fill_8 FILLER_0_17_608 ();
 sg13g2_fill_8 FILLER_0_17_616 ();
 sg13g2_fill_8 FILLER_0_17_624 ();
 sg13g2_fill_8 FILLER_0_17_632 ();
 sg13g2_fill_8 FILLER_0_17_640 ();
 sg13g2_fill_8 FILLER_0_17_648 ();
 sg13g2_fill_8 FILLER_0_17_656 ();
 sg13g2_fill_8 FILLER_0_17_664 ();
 sg13g2_fill_8 FILLER_0_17_672 ();
 sg13g2_fill_8 FILLER_0_17_680 ();
 sg13g2_fill_8 FILLER_0_17_688 ();
 sg13g2_fill_8 FILLER_0_17_696 ();
 sg13g2_fill_8 FILLER_0_17_704 ();
 sg13g2_fill_8 FILLER_0_17_712 ();
 sg13g2_fill_8 FILLER_0_17_720 ();
 sg13g2_fill_8 FILLER_0_17_728 ();
 sg13g2_fill_8 FILLER_0_17_736 ();
 sg13g2_fill_8 FILLER_0_17_744 ();
 sg13g2_fill_8 FILLER_0_17_752 ();
 sg13g2_fill_8 FILLER_0_17_760 ();
 sg13g2_fill_8 FILLER_0_17_768 ();
 sg13g2_fill_8 FILLER_0_17_776 ();
 sg13g2_fill_8 FILLER_0_17_784 ();
 sg13g2_fill_8 FILLER_0_17_792 ();
 sg13g2_fill_8 FILLER_0_17_800 ();
 sg13g2_fill_8 FILLER_0_17_808 ();
 sg13g2_fill_8 FILLER_0_17_816 ();
 sg13g2_fill_8 FILLER_0_17_824 ();
 sg13g2_fill_8 FILLER_0_17_832 ();
 sg13g2_fill_8 FILLER_0_17_840 ();
 sg13g2_fill_8 FILLER_0_17_848 ();
 sg13g2_fill_8 FILLER_0_17_856 ();
 sg13g2_fill_8 FILLER_0_17_864 ();
 sg13g2_fill_8 FILLER_0_17_872 ();
 sg13g2_fill_8 FILLER_0_17_880 ();
 sg13g2_fill_8 FILLER_0_17_888 ();
 sg13g2_fill_8 FILLER_0_17_896 ();
 sg13g2_fill_8 FILLER_0_17_904 ();
 sg13g2_fill_8 FILLER_0_17_912 ();
 sg13g2_fill_8 FILLER_0_17_920 ();
 sg13g2_fill_8 FILLER_0_17_928 ();
 sg13g2_fill_8 FILLER_0_17_936 ();
 sg13g2_fill_8 FILLER_0_17_944 ();
 sg13g2_fill_8 FILLER_0_17_952 ();
 sg13g2_fill_8 FILLER_0_17_960 ();
 sg13g2_fill_8 FILLER_0_17_968 ();
 sg13g2_fill_8 FILLER_0_17_976 ();
 sg13g2_fill_8 FILLER_0_17_984 ();
 sg13g2_fill_8 FILLER_0_17_992 ();
 sg13g2_fill_8 FILLER_0_17_1000 ();
 sg13g2_fill_8 FILLER_0_17_1008 ();
 sg13g2_fill_8 FILLER_0_17_1016 ();
 sg13g2_fill_8 FILLER_0_17_1024 ();
 sg13g2_fill_8 FILLER_0_17_1032 ();
 sg13g2_fill_8 FILLER_0_17_1040 ();
 sg13g2_fill_8 FILLER_0_17_1048 ();
 sg13g2_fill_8 FILLER_0_17_1056 ();
 sg13g2_fill_8 FILLER_0_17_1064 ();
 sg13g2_fill_8 FILLER_0_17_1072 ();
 sg13g2_fill_8 FILLER_0_17_1080 ();
 sg13g2_fill_8 FILLER_0_17_1088 ();
 sg13g2_fill_8 FILLER_0_17_1096 ();
 sg13g2_fill_8 FILLER_0_17_1104 ();
 sg13g2_fill_8 FILLER_0_17_1112 ();
 sg13g2_fill_8 FILLER_0_17_1120 ();
 sg13g2_fill_8 FILLER_0_17_1128 ();
 sg13g2_fill_8 FILLER_0_17_1136 ();
 sg13g2_fill_8 FILLER_0_17_1144 ();
 sg13g2_fill_8 FILLER_0_17_1152 ();
 sg13g2_fill_8 FILLER_0_17_1160 ();
 sg13g2_fill_8 FILLER_0_17_1168 ();
 sg13g2_fill_8 FILLER_0_17_1176 ();
 sg13g2_fill_8 FILLER_0_17_1184 ();
 sg13g2_fill_8 FILLER_0_17_1192 ();
 sg13g2_fill_8 FILLER_0_17_1200 ();
 sg13g2_fill_8 FILLER_0_17_1208 ();
 sg13g2_fill_8 FILLER_0_17_1216 ();
 sg13g2_fill_4 FILLER_0_17_1224 ();
 sg13g2_fill_8 FILLER_0_18_0 ();
 sg13g2_fill_8 FILLER_0_18_8 ();
 sg13g2_fill_8 FILLER_0_18_16 ();
 sg13g2_fill_8 FILLER_0_18_24 ();
 sg13g2_fill_8 FILLER_0_18_32 ();
 sg13g2_fill_8 FILLER_0_18_40 ();
 sg13g2_fill_8 FILLER_0_18_48 ();
 sg13g2_fill_8 FILLER_0_18_56 ();
 sg13g2_fill_8 FILLER_0_18_64 ();
 sg13g2_fill_8 FILLER_0_18_72 ();
 sg13g2_fill_8 FILLER_0_18_80 ();
 sg13g2_fill_8 FILLER_0_18_88 ();
 sg13g2_fill_8 FILLER_0_18_96 ();
 sg13g2_fill_8 FILLER_0_18_104 ();
 sg13g2_fill_8 FILLER_0_18_112 ();
 sg13g2_fill_8 FILLER_0_18_120 ();
 sg13g2_fill_8 FILLER_0_18_128 ();
 sg13g2_fill_8 FILLER_0_18_136 ();
 sg13g2_fill_8 FILLER_0_18_144 ();
 sg13g2_fill_8 FILLER_0_18_152 ();
 sg13g2_fill_8 FILLER_0_18_160 ();
 sg13g2_fill_8 FILLER_0_18_168 ();
 sg13g2_fill_8 FILLER_0_18_176 ();
 sg13g2_fill_8 FILLER_0_18_184 ();
 sg13g2_fill_8 FILLER_0_18_192 ();
 sg13g2_fill_8 FILLER_0_18_200 ();
 sg13g2_fill_8 FILLER_0_18_208 ();
 sg13g2_fill_8 FILLER_0_18_216 ();
 sg13g2_fill_8 FILLER_0_18_224 ();
 sg13g2_fill_8 FILLER_0_18_232 ();
 sg13g2_fill_8 FILLER_0_18_240 ();
 sg13g2_fill_8 FILLER_0_18_248 ();
 sg13g2_fill_8 FILLER_0_18_256 ();
 sg13g2_fill_8 FILLER_0_18_264 ();
 sg13g2_fill_8 FILLER_0_18_272 ();
 sg13g2_fill_8 FILLER_0_18_280 ();
 sg13g2_fill_8 FILLER_0_18_288 ();
 sg13g2_fill_8 FILLER_0_18_296 ();
 sg13g2_fill_8 FILLER_0_18_304 ();
 sg13g2_fill_8 FILLER_0_18_312 ();
 sg13g2_fill_8 FILLER_0_18_320 ();
 sg13g2_fill_8 FILLER_0_18_328 ();
 sg13g2_fill_8 FILLER_0_18_336 ();
 sg13g2_fill_8 FILLER_0_18_344 ();
 sg13g2_fill_8 FILLER_0_18_352 ();
 sg13g2_fill_8 FILLER_0_18_360 ();
 sg13g2_fill_8 FILLER_0_18_368 ();
 sg13g2_fill_8 FILLER_0_18_376 ();
 sg13g2_fill_8 FILLER_0_18_384 ();
 sg13g2_fill_8 FILLER_0_18_392 ();
 sg13g2_fill_8 FILLER_0_18_400 ();
 sg13g2_fill_8 FILLER_0_18_408 ();
 sg13g2_fill_8 FILLER_0_18_416 ();
 sg13g2_fill_8 FILLER_0_18_424 ();
 sg13g2_fill_8 FILLER_0_18_432 ();
 sg13g2_fill_8 FILLER_0_18_440 ();
 sg13g2_fill_8 FILLER_0_18_448 ();
 sg13g2_fill_8 FILLER_0_18_456 ();
 sg13g2_fill_8 FILLER_0_18_464 ();
 sg13g2_fill_8 FILLER_0_18_472 ();
 sg13g2_fill_8 FILLER_0_18_480 ();
 sg13g2_fill_8 FILLER_0_18_488 ();
 sg13g2_fill_8 FILLER_0_18_496 ();
 sg13g2_fill_8 FILLER_0_18_504 ();
 sg13g2_fill_8 FILLER_0_18_512 ();
 sg13g2_fill_8 FILLER_0_18_520 ();
 sg13g2_fill_8 FILLER_0_18_528 ();
 sg13g2_fill_8 FILLER_0_18_536 ();
 sg13g2_fill_8 FILLER_0_18_544 ();
 sg13g2_fill_8 FILLER_0_18_552 ();
 sg13g2_fill_8 FILLER_0_18_560 ();
 sg13g2_fill_8 FILLER_0_18_568 ();
 sg13g2_fill_8 FILLER_0_18_576 ();
 sg13g2_fill_8 FILLER_0_18_584 ();
 sg13g2_fill_8 FILLER_0_18_592 ();
 sg13g2_fill_8 FILLER_0_18_600 ();
 sg13g2_fill_8 FILLER_0_18_608 ();
 sg13g2_fill_8 FILLER_0_18_616 ();
 sg13g2_fill_8 FILLER_0_18_624 ();
 sg13g2_fill_8 FILLER_0_18_632 ();
 sg13g2_fill_8 FILLER_0_18_640 ();
 sg13g2_fill_8 FILLER_0_18_648 ();
 sg13g2_fill_8 FILLER_0_18_656 ();
 sg13g2_fill_8 FILLER_0_18_664 ();
 sg13g2_fill_8 FILLER_0_18_672 ();
 sg13g2_fill_8 FILLER_0_18_680 ();
 sg13g2_fill_8 FILLER_0_18_688 ();
 sg13g2_fill_8 FILLER_0_18_696 ();
 sg13g2_fill_8 FILLER_0_18_704 ();
 sg13g2_fill_8 FILLER_0_18_712 ();
 sg13g2_fill_8 FILLER_0_18_720 ();
 sg13g2_fill_8 FILLER_0_18_728 ();
 sg13g2_fill_8 FILLER_0_18_736 ();
 sg13g2_fill_8 FILLER_0_18_744 ();
 sg13g2_fill_8 FILLER_0_18_752 ();
 sg13g2_fill_8 FILLER_0_18_760 ();
 sg13g2_fill_8 FILLER_0_18_768 ();
 sg13g2_fill_8 FILLER_0_18_776 ();
 sg13g2_fill_8 FILLER_0_18_784 ();
 sg13g2_fill_8 FILLER_0_18_792 ();
 sg13g2_fill_8 FILLER_0_18_800 ();
 sg13g2_fill_8 FILLER_0_18_808 ();
 sg13g2_fill_8 FILLER_0_18_816 ();
 sg13g2_fill_8 FILLER_0_18_824 ();
 sg13g2_fill_8 FILLER_0_18_832 ();
 sg13g2_fill_8 FILLER_0_18_840 ();
 sg13g2_fill_8 FILLER_0_18_848 ();
 sg13g2_fill_8 FILLER_0_18_856 ();
 sg13g2_fill_8 FILLER_0_18_864 ();
 sg13g2_fill_8 FILLER_0_18_872 ();
 sg13g2_fill_8 FILLER_0_18_880 ();
 sg13g2_fill_8 FILLER_0_18_888 ();
 sg13g2_fill_8 FILLER_0_18_896 ();
 sg13g2_fill_8 FILLER_0_18_904 ();
 sg13g2_fill_8 FILLER_0_18_912 ();
 sg13g2_fill_8 FILLER_0_18_920 ();
 sg13g2_fill_8 FILLER_0_18_928 ();
 sg13g2_fill_8 FILLER_0_18_936 ();
 sg13g2_fill_8 FILLER_0_18_944 ();
 sg13g2_fill_8 FILLER_0_18_952 ();
 sg13g2_fill_8 FILLER_0_18_960 ();
 sg13g2_fill_8 FILLER_0_18_968 ();
 sg13g2_fill_8 FILLER_0_18_976 ();
 sg13g2_fill_8 FILLER_0_18_984 ();
 sg13g2_fill_8 FILLER_0_18_992 ();
 sg13g2_fill_8 FILLER_0_18_1000 ();
 sg13g2_fill_8 FILLER_0_18_1008 ();
 sg13g2_fill_8 FILLER_0_18_1016 ();
 sg13g2_fill_8 FILLER_0_18_1024 ();
 sg13g2_fill_8 FILLER_0_18_1032 ();
 sg13g2_fill_8 FILLER_0_18_1040 ();
 sg13g2_fill_8 FILLER_0_18_1048 ();
 sg13g2_fill_8 FILLER_0_18_1056 ();
 sg13g2_fill_8 FILLER_0_18_1064 ();
 sg13g2_fill_8 FILLER_0_18_1072 ();
 sg13g2_fill_8 FILLER_0_18_1080 ();
 sg13g2_fill_8 FILLER_0_18_1088 ();
 sg13g2_fill_8 FILLER_0_18_1096 ();
 sg13g2_fill_8 FILLER_0_18_1104 ();
 sg13g2_fill_8 FILLER_0_18_1112 ();
 sg13g2_fill_8 FILLER_0_18_1120 ();
 sg13g2_fill_8 FILLER_0_18_1128 ();
 sg13g2_fill_8 FILLER_0_18_1136 ();
 sg13g2_fill_8 FILLER_0_18_1144 ();
 sg13g2_fill_8 FILLER_0_18_1152 ();
 sg13g2_fill_8 FILLER_0_18_1160 ();
 sg13g2_fill_8 FILLER_0_18_1168 ();
 sg13g2_fill_8 FILLER_0_18_1176 ();
 sg13g2_fill_8 FILLER_0_18_1184 ();
 sg13g2_fill_8 FILLER_0_18_1192 ();
 sg13g2_fill_8 FILLER_0_18_1200 ();
 sg13g2_fill_8 FILLER_0_18_1208 ();
 sg13g2_fill_8 FILLER_0_18_1216 ();
 sg13g2_fill_4 FILLER_0_18_1224 ();
 sg13g2_fill_8 FILLER_0_19_0 ();
 sg13g2_fill_8 FILLER_0_19_8 ();
 sg13g2_fill_8 FILLER_0_19_16 ();
 sg13g2_fill_8 FILLER_0_19_24 ();
 sg13g2_fill_8 FILLER_0_19_32 ();
 sg13g2_fill_8 FILLER_0_19_40 ();
 sg13g2_fill_8 FILLER_0_19_48 ();
 sg13g2_fill_8 FILLER_0_19_56 ();
 sg13g2_fill_8 FILLER_0_19_64 ();
 sg13g2_fill_8 FILLER_0_19_72 ();
 sg13g2_fill_8 FILLER_0_19_80 ();
 sg13g2_fill_8 FILLER_0_19_88 ();
 sg13g2_fill_8 FILLER_0_19_96 ();
 sg13g2_fill_8 FILLER_0_19_104 ();
 sg13g2_fill_8 FILLER_0_19_112 ();
 sg13g2_fill_8 FILLER_0_19_120 ();
 sg13g2_fill_8 FILLER_0_19_128 ();
 sg13g2_fill_8 FILLER_0_19_136 ();
 sg13g2_fill_8 FILLER_0_19_144 ();
 sg13g2_fill_8 FILLER_0_19_152 ();
 sg13g2_fill_8 FILLER_0_19_160 ();
 sg13g2_fill_8 FILLER_0_19_168 ();
 sg13g2_fill_8 FILLER_0_19_176 ();
 sg13g2_fill_8 FILLER_0_19_184 ();
 sg13g2_fill_8 FILLER_0_19_192 ();
 sg13g2_fill_8 FILLER_0_19_200 ();
 sg13g2_fill_8 FILLER_0_19_208 ();
 sg13g2_fill_8 FILLER_0_19_216 ();
 sg13g2_fill_8 FILLER_0_19_224 ();
 sg13g2_fill_8 FILLER_0_19_232 ();
 sg13g2_fill_8 FILLER_0_19_240 ();
 sg13g2_fill_8 FILLER_0_19_248 ();
 sg13g2_fill_8 FILLER_0_19_256 ();
 sg13g2_fill_8 FILLER_0_19_264 ();
 sg13g2_fill_8 FILLER_0_19_272 ();
 sg13g2_fill_8 FILLER_0_19_280 ();
 sg13g2_fill_8 FILLER_0_19_288 ();
 sg13g2_fill_8 FILLER_0_19_296 ();
 sg13g2_fill_8 FILLER_0_19_304 ();
 sg13g2_fill_8 FILLER_0_19_312 ();
 sg13g2_fill_8 FILLER_0_19_320 ();
 sg13g2_fill_8 FILLER_0_19_328 ();
 sg13g2_fill_8 FILLER_0_19_336 ();
 sg13g2_fill_8 FILLER_0_19_344 ();
 sg13g2_fill_8 FILLER_0_19_352 ();
 sg13g2_fill_8 FILLER_0_19_360 ();
 sg13g2_fill_8 FILLER_0_19_368 ();
 sg13g2_fill_8 FILLER_0_19_376 ();
 sg13g2_fill_8 FILLER_0_19_384 ();
 sg13g2_fill_8 FILLER_0_19_392 ();
 sg13g2_fill_8 FILLER_0_19_400 ();
 sg13g2_fill_8 FILLER_0_19_408 ();
 sg13g2_fill_8 FILLER_0_19_416 ();
 sg13g2_fill_8 FILLER_0_19_424 ();
 sg13g2_fill_8 FILLER_0_19_432 ();
 sg13g2_fill_8 FILLER_0_19_440 ();
 sg13g2_fill_8 FILLER_0_19_448 ();
 sg13g2_fill_8 FILLER_0_19_456 ();
 sg13g2_fill_8 FILLER_0_19_464 ();
 sg13g2_fill_8 FILLER_0_19_472 ();
 sg13g2_fill_8 FILLER_0_19_480 ();
 sg13g2_fill_8 FILLER_0_19_488 ();
 sg13g2_fill_8 FILLER_0_19_496 ();
 sg13g2_fill_8 FILLER_0_19_504 ();
 sg13g2_fill_8 FILLER_0_19_512 ();
 sg13g2_fill_8 FILLER_0_19_520 ();
 sg13g2_fill_8 FILLER_0_19_528 ();
 sg13g2_fill_8 FILLER_0_19_536 ();
 sg13g2_fill_8 FILLER_0_19_544 ();
 sg13g2_fill_8 FILLER_0_19_552 ();
 sg13g2_fill_8 FILLER_0_19_560 ();
 sg13g2_fill_8 FILLER_0_19_568 ();
 sg13g2_fill_8 FILLER_0_19_576 ();
 sg13g2_fill_8 FILLER_0_19_584 ();
 sg13g2_fill_8 FILLER_0_19_592 ();
 sg13g2_fill_8 FILLER_0_19_600 ();
 sg13g2_fill_8 FILLER_0_19_608 ();
 sg13g2_fill_8 FILLER_0_19_616 ();
 sg13g2_fill_8 FILLER_0_19_624 ();
 sg13g2_fill_8 FILLER_0_19_632 ();
 sg13g2_fill_8 FILLER_0_19_640 ();
 sg13g2_fill_8 FILLER_0_19_648 ();
 sg13g2_fill_8 FILLER_0_19_656 ();
 sg13g2_fill_8 FILLER_0_19_664 ();
 sg13g2_fill_8 FILLER_0_19_672 ();
 sg13g2_fill_8 FILLER_0_19_680 ();
 sg13g2_fill_8 FILLER_0_19_688 ();
 sg13g2_fill_8 FILLER_0_19_696 ();
 sg13g2_fill_8 FILLER_0_19_704 ();
 sg13g2_fill_8 FILLER_0_19_712 ();
 sg13g2_fill_8 FILLER_0_19_720 ();
 sg13g2_fill_8 FILLER_0_19_728 ();
 sg13g2_fill_8 FILLER_0_19_736 ();
 sg13g2_fill_8 FILLER_0_19_744 ();
 sg13g2_fill_8 FILLER_0_19_752 ();
 sg13g2_fill_8 FILLER_0_19_760 ();
 sg13g2_fill_8 FILLER_0_19_768 ();
 sg13g2_fill_8 FILLER_0_19_776 ();
 sg13g2_fill_8 FILLER_0_19_784 ();
 sg13g2_fill_8 FILLER_0_19_792 ();
 sg13g2_fill_8 FILLER_0_19_800 ();
 sg13g2_fill_8 FILLER_0_19_808 ();
 sg13g2_fill_8 FILLER_0_19_816 ();
 sg13g2_fill_8 FILLER_0_19_824 ();
 sg13g2_fill_8 FILLER_0_19_832 ();
 sg13g2_fill_8 FILLER_0_19_840 ();
 sg13g2_fill_8 FILLER_0_19_848 ();
 sg13g2_fill_8 FILLER_0_19_856 ();
 sg13g2_fill_8 FILLER_0_19_864 ();
 sg13g2_fill_8 FILLER_0_19_872 ();
 sg13g2_fill_8 FILLER_0_19_880 ();
 sg13g2_fill_8 FILLER_0_19_888 ();
 sg13g2_fill_8 FILLER_0_19_896 ();
 sg13g2_fill_8 FILLER_0_19_904 ();
 sg13g2_fill_8 FILLER_0_19_912 ();
 sg13g2_fill_8 FILLER_0_19_920 ();
 sg13g2_fill_8 FILLER_0_19_928 ();
 sg13g2_fill_8 FILLER_0_19_936 ();
 sg13g2_fill_8 FILLER_0_19_944 ();
 sg13g2_fill_8 FILLER_0_19_952 ();
 sg13g2_fill_8 FILLER_0_19_960 ();
 sg13g2_fill_8 FILLER_0_19_968 ();
 sg13g2_fill_8 FILLER_0_19_976 ();
 sg13g2_fill_8 FILLER_0_19_984 ();
 sg13g2_fill_8 FILLER_0_19_992 ();
 sg13g2_fill_8 FILLER_0_19_1000 ();
 sg13g2_fill_8 FILLER_0_19_1008 ();
 sg13g2_fill_8 FILLER_0_19_1016 ();
 sg13g2_fill_8 FILLER_0_19_1024 ();
 sg13g2_fill_8 FILLER_0_19_1032 ();
 sg13g2_fill_8 FILLER_0_19_1040 ();
 sg13g2_fill_8 FILLER_0_19_1048 ();
 sg13g2_fill_8 FILLER_0_19_1056 ();
 sg13g2_fill_8 FILLER_0_19_1064 ();
 sg13g2_fill_8 FILLER_0_19_1072 ();
 sg13g2_fill_8 FILLER_0_19_1080 ();
 sg13g2_fill_8 FILLER_0_19_1088 ();
 sg13g2_fill_8 FILLER_0_19_1096 ();
 sg13g2_fill_8 FILLER_0_19_1104 ();
 sg13g2_fill_8 FILLER_0_19_1112 ();
 sg13g2_fill_8 FILLER_0_19_1120 ();
 sg13g2_fill_8 FILLER_0_19_1128 ();
 sg13g2_fill_8 FILLER_0_19_1136 ();
 sg13g2_fill_8 FILLER_0_19_1144 ();
 sg13g2_fill_8 FILLER_0_19_1152 ();
 sg13g2_fill_8 FILLER_0_19_1160 ();
 sg13g2_fill_8 FILLER_0_19_1168 ();
 sg13g2_fill_8 FILLER_0_19_1176 ();
 sg13g2_fill_8 FILLER_0_19_1184 ();
 sg13g2_fill_8 FILLER_0_19_1192 ();
 sg13g2_fill_8 FILLER_0_19_1200 ();
 sg13g2_fill_8 FILLER_0_19_1208 ();
 sg13g2_fill_8 FILLER_0_19_1216 ();
 sg13g2_fill_4 FILLER_0_19_1224 ();
 sg13g2_fill_8 FILLER_0_20_0 ();
 sg13g2_fill_8 FILLER_0_20_8 ();
 sg13g2_fill_8 FILLER_0_20_16 ();
 sg13g2_fill_8 FILLER_0_20_24 ();
 sg13g2_fill_8 FILLER_0_20_32 ();
 sg13g2_fill_8 FILLER_0_20_40 ();
 sg13g2_fill_8 FILLER_0_20_48 ();
 sg13g2_fill_8 FILLER_0_20_56 ();
 sg13g2_fill_8 FILLER_0_20_64 ();
 sg13g2_fill_8 FILLER_0_20_72 ();
 sg13g2_fill_8 FILLER_0_20_80 ();
 sg13g2_fill_8 FILLER_0_20_88 ();
 sg13g2_fill_8 FILLER_0_20_96 ();
 sg13g2_fill_8 FILLER_0_20_104 ();
 sg13g2_fill_8 FILLER_0_20_112 ();
 sg13g2_fill_8 FILLER_0_20_120 ();
 sg13g2_fill_8 FILLER_0_20_128 ();
 sg13g2_fill_8 FILLER_0_20_136 ();
 sg13g2_fill_8 FILLER_0_20_144 ();
 sg13g2_fill_8 FILLER_0_20_152 ();
 sg13g2_fill_8 FILLER_0_20_160 ();
 sg13g2_fill_8 FILLER_0_20_168 ();
 sg13g2_fill_8 FILLER_0_20_176 ();
 sg13g2_fill_8 FILLER_0_20_184 ();
 sg13g2_fill_8 FILLER_0_20_192 ();
 sg13g2_fill_8 FILLER_0_20_200 ();
 sg13g2_fill_8 FILLER_0_20_208 ();
 sg13g2_fill_8 FILLER_0_20_216 ();
 sg13g2_fill_8 FILLER_0_20_224 ();
 sg13g2_fill_8 FILLER_0_20_232 ();
 sg13g2_fill_8 FILLER_0_20_240 ();
 sg13g2_fill_8 FILLER_0_20_248 ();
 sg13g2_fill_8 FILLER_0_20_256 ();
 sg13g2_fill_8 FILLER_0_20_264 ();
 sg13g2_fill_8 FILLER_0_20_272 ();
 sg13g2_fill_8 FILLER_0_20_280 ();
 sg13g2_fill_8 FILLER_0_20_288 ();
 sg13g2_fill_8 FILLER_0_20_296 ();
 sg13g2_fill_8 FILLER_0_20_304 ();
 sg13g2_fill_8 FILLER_0_20_312 ();
 sg13g2_fill_8 FILLER_0_20_320 ();
 sg13g2_fill_8 FILLER_0_20_328 ();
 sg13g2_fill_8 FILLER_0_20_336 ();
 sg13g2_fill_8 FILLER_0_20_344 ();
 sg13g2_fill_8 FILLER_0_20_352 ();
 sg13g2_fill_8 FILLER_0_20_360 ();
 sg13g2_fill_8 FILLER_0_20_368 ();
 sg13g2_fill_8 FILLER_0_20_376 ();
 sg13g2_fill_8 FILLER_0_20_384 ();
 sg13g2_fill_8 FILLER_0_20_392 ();
 sg13g2_fill_8 FILLER_0_20_400 ();
 sg13g2_fill_8 FILLER_0_20_408 ();
 sg13g2_fill_8 FILLER_0_20_416 ();
 sg13g2_fill_8 FILLER_0_20_424 ();
 sg13g2_fill_8 FILLER_0_20_432 ();
 sg13g2_fill_8 FILLER_0_20_440 ();
 sg13g2_fill_8 FILLER_0_20_448 ();
 sg13g2_fill_8 FILLER_0_20_456 ();
 sg13g2_fill_8 FILLER_0_20_464 ();
 sg13g2_fill_8 FILLER_0_20_472 ();
 sg13g2_fill_8 FILLER_0_20_480 ();
 sg13g2_fill_8 FILLER_0_20_488 ();
 sg13g2_fill_8 FILLER_0_20_496 ();
 sg13g2_fill_8 FILLER_0_20_504 ();
 sg13g2_fill_8 FILLER_0_20_512 ();
 sg13g2_fill_8 FILLER_0_20_520 ();
 sg13g2_fill_8 FILLER_0_20_528 ();
 sg13g2_fill_8 FILLER_0_20_536 ();
 sg13g2_fill_8 FILLER_0_20_544 ();
 sg13g2_fill_8 FILLER_0_20_552 ();
 sg13g2_fill_8 FILLER_0_20_560 ();
 sg13g2_fill_8 FILLER_0_20_568 ();
 sg13g2_fill_8 FILLER_0_20_576 ();
 sg13g2_fill_8 FILLER_0_20_584 ();
 sg13g2_fill_8 FILLER_0_20_592 ();
 sg13g2_fill_8 FILLER_0_20_600 ();
 sg13g2_fill_8 FILLER_0_20_608 ();
 sg13g2_fill_8 FILLER_0_20_616 ();
 sg13g2_fill_8 FILLER_0_20_624 ();
 sg13g2_fill_8 FILLER_0_20_632 ();
 sg13g2_fill_8 FILLER_0_20_640 ();
 sg13g2_fill_8 FILLER_0_20_648 ();
 sg13g2_fill_8 FILLER_0_20_656 ();
 sg13g2_fill_8 FILLER_0_20_664 ();
 sg13g2_fill_8 FILLER_0_20_672 ();
 sg13g2_fill_8 FILLER_0_20_680 ();
 sg13g2_fill_8 FILLER_0_20_688 ();
 sg13g2_fill_8 FILLER_0_20_696 ();
 sg13g2_fill_8 FILLER_0_20_704 ();
 sg13g2_fill_8 FILLER_0_20_712 ();
 sg13g2_fill_8 FILLER_0_20_720 ();
 sg13g2_fill_8 FILLER_0_20_728 ();
 sg13g2_fill_8 FILLER_0_20_736 ();
 sg13g2_fill_8 FILLER_0_20_744 ();
 sg13g2_fill_8 FILLER_0_20_752 ();
 sg13g2_fill_8 FILLER_0_20_760 ();
 sg13g2_fill_8 FILLER_0_20_768 ();
 sg13g2_fill_8 FILLER_0_20_776 ();
 sg13g2_fill_8 FILLER_0_20_784 ();
 sg13g2_fill_8 FILLER_0_20_792 ();
 sg13g2_fill_8 FILLER_0_20_800 ();
 sg13g2_fill_8 FILLER_0_20_808 ();
 sg13g2_fill_8 FILLER_0_20_816 ();
 sg13g2_fill_8 FILLER_0_20_824 ();
 sg13g2_fill_8 FILLER_0_20_832 ();
 sg13g2_fill_8 FILLER_0_20_840 ();
 sg13g2_fill_8 FILLER_0_20_848 ();
 sg13g2_fill_8 FILLER_0_20_856 ();
 sg13g2_fill_8 FILLER_0_20_864 ();
 sg13g2_fill_8 FILLER_0_20_872 ();
 sg13g2_fill_8 FILLER_0_20_880 ();
 sg13g2_fill_8 FILLER_0_20_888 ();
 sg13g2_fill_8 FILLER_0_20_896 ();
 sg13g2_fill_8 FILLER_0_20_904 ();
 sg13g2_fill_8 FILLER_0_20_912 ();
 sg13g2_fill_8 FILLER_0_20_920 ();
 sg13g2_fill_8 FILLER_0_20_928 ();
 sg13g2_fill_8 FILLER_0_20_936 ();
 sg13g2_fill_8 FILLER_0_20_944 ();
 sg13g2_fill_8 FILLER_0_20_952 ();
 sg13g2_fill_8 FILLER_0_20_960 ();
 sg13g2_fill_8 FILLER_0_20_968 ();
 sg13g2_fill_8 FILLER_0_20_976 ();
 sg13g2_fill_8 FILLER_0_20_984 ();
 sg13g2_fill_8 FILLER_0_20_992 ();
 sg13g2_fill_8 FILLER_0_20_1000 ();
 sg13g2_fill_8 FILLER_0_20_1008 ();
 sg13g2_fill_8 FILLER_0_20_1016 ();
 sg13g2_fill_8 FILLER_0_20_1024 ();
 sg13g2_fill_8 FILLER_0_20_1032 ();
 sg13g2_fill_8 FILLER_0_20_1040 ();
 sg13g2_fill_8 FILLER_0_20_1048 ();
 sg13g2_fill_8 FILLER_0_20_1056 ();
 sg13g2_fill_8 FILLER_0_20_1064 ();
 sg13g2_fill_8 FILLER_0_20_1072 ();
 sg13g2_fill_8 FILLER_0_20_1080 ();
 sg13g2_fill_8 FILLER_0_20_1088 ();
 sg13g2_fill_8 FILLER_0_20_1096 ();
 sg13g2_fill_8 FILLER_0_20_1104 ();
 sg13g2_fill_8 FILLER_0_20_1112 ();
 sg13g2_fill_8 FILLER_0_20_1120 ();
 sg13g2_fill_8 FILLER_0_20_1128 ();
 sg13g2_fill_8 FILLER_0_20_1136 ();
 sg13g2_fill_8 FILLER_0_20_1144 ();
 sg13g2_fill_8 FILLER_0_20_1152 ();
 sg13g2_fill_8 FILLER_0_20_1160 ();
 sg13g2_fill_8 FILLER_0_20_1168 ();
 sg13g2_fill_8 FILLER_0_20_1176 ();
 sg13g2_fill_8 FILLER_0_20_1184 ();
 sg13g2_fill_8 FILLER_0_20_1192 ();
 sg13g2_fill_8 FILLER_0_20_1200 ();
 sg13g2_fill_8 FILLER_0_20_1208 ();
 sg13g2_fill_8 FILLER_0_20_1216 ();
 sg13g2_fill_4 FILLER_0_20_1224 ();
 sg13g2_fill_8 FILLER_0_21_0 ();
 sg13g2_fill_8 FILLER_0_21_8 ();
 sg13g2_fill_8 FILLER_0_21_16 ();
 sg13g2_fill_8 FILLER_0_21_24 ();
 sg13g2_fill_8 FILLER_0_21_32 ();
 sg13g2_fill_8 FILLER_0_21_40 ();
 sg13g2_fill_8 FILLER_0_21_48 ();
 sg13g2_fill_8 FILLER_0_21_56 ();
 sg13g2_fill_8 FILLER_0_21_64 ();
 sg13g2_fill_8 FILLER_0_21_72 ();
 sg13g2_fill_8 FILLER_0_21_80 ();
 sg13g2_fill_8 FILLER_0_21_88 ();
 sg13g2_fill_8 FILLER_0_21_96 ();
 sg13g2_fill_8 FILLER_0_21_104 ();
 sg13g2_fill_8 FILLER_0_21_112 ();
 sg13g2_fill_8 FILLER_0_21_120 ();
 sg13g2_fill_8 FILLER_0_21_128 ();
 sg13g2_fill_8 FILLER_0_21_136 ();
 sg13g2_fill_8 FILLER_0_21_144 ();
 sg13g2_fill_8 FILLER_0_21_152 ();
 sg13g2_fill_8 FILLER_0_21_160 ();
 sg13g2_fill_8 FILLER_0_21_168 ();
 sg13g2_fill_4 FILLER_0_21_176 ();
 sg13g2_fill_8 FILLER_0_21_185 ();
 sg13g2_fill_2 FILLER_0_21_193 ();
 sg13g2_fill_1 FILLER_0_21_195 ();
 sg13g2_fill_2 FILLER_0_21_201 ();
 sg13g2_fill_8 FILLER_0_21_208 ();
 sg13g2_fill_8 FILLER_0_21_216 ();
 sg13g2_fill_8 FILLER_0_21_224 ();
 sg13g2_fill_8 FILLER_0_21_232 ();
 sg13g2_fill_8 FILLER_0_21_240 ();
 sg13g2_fill_8 FILLER_0_21_248 ();
 sg13g2_fill_2 FILLER_0_21_256 ();
 sg13g2_fill_8 FILLER_0_21_262 ();
 sg13g2_fill_8 FILLER_0_21_270 ();
 sg13g2_fill_8 FILLER_0_21_278 ();
 sg13g2_fill_8 FILLER_0_21_286 ();
 sg13g2_fill_8 FILLER_0_21_294 ();
 sg13g2_fill_8 FILLER_0_21_302 ();
 sg13g2_fill_8 FILLER_0_21_310 ();
 sg13g2_fill_8 FILLER_0_21_318 ();
 sg13g2_fill_4 FILLER_0_21_326 ();
 sg13g2_fill_2 FILLER_0_21_330 ();
 sg13g2_fill_8 FILLER_0_21_337 ();
 sg13g2_fill_8 FILLER_0_21_345 ();
 sg13g2_fill_8 FILLER_0_21_353 ();
 sg13g2_fill_2 FILLER_0_21_371 ();
 sg13g2_fill_1 FILLER_0_21_373 ();
 sg13g2_fill_1 FILLER_0_21_379 ();
 sg13g2_fill_8 FILLER_0_21_384 ();
 sg13g2_fill_8 FILLER_0_21_392 ();
 sg13g2_fill_8 FILLER_0_21_400 ();
 sg13g2_fill_8 FILLER_0_21_408 ();
 sg13g2_fill_8 FILLER_0_21_416 ();
 sg13g2_fill_8 FILLER_0_21_424 ();
 sg13g2_fill_8 FILLER_0_21_432 ();
 sg13g2_fill_8 FILLER_0_21_440 ();
 sg13g2_fill_8 FILLER_0_21_448 ();
 sg13g2_fill_8 FILLER_0_21_456 ();
 sg13g2_fill_8 FILLER_0_21_464 ();
 sg13g2_fill_8 FILLER_0_21_472 ();
 sg13g2_fill_8 FILLER_0_21_480 ();
 sg13g2_fill_8 FILLER_0_21_488 ();
 sg13g2_fill_8 FILLER_0_21_496 ();
 sg13g2_fill_8 FILLER_0_21_504 ();
 sg13g2_fill_8 FILLER_0_21_512 ();
 sg13g2_fill_8 FILLER_0_21_520 ();
 sg13g2_fill_8 FILLER_0_21_528 ();
 sg13g2_fill_8 FILLER_0_21_536 ();
 sg13g2_fill_8 FILLER_0_21_544 ();
 sg13g2_fill_8 FILLER_0_21_552 ();
 sg13g2_fill_8 FILLER_0_21_560 ();
 sg13g2_fill_8 FILLER_0_21_568 ();
 sg13g2_fill_8 FILLER_0_21_576 ();
 sg13g2_fill_8 FILLER_0_21_584 ();
 sg13g2_fill_8 FILLER_0_21_592 ();
 sg13g2_fill_8 FILLER_0_21_600 ();
 sg13g2_fill_8 FILLER_0_21_608 ();
 sg13g2_fill_8 FILLER_0_21_616 ();
 sg13g2_fill_8 FILLER_0_21_624 ();
 sg13g2_fill_8 FILLER_0_21_632 ();
 sg13g2_fill_8 FILLER_0_21_640 ();
 sg13g2_fill_8 FILLER_0_21_648 ();
 sg13g2_fill_8 FILLER_0_21_656 ();
 sg13g2_fill_8 FILLER_0_21_664 ();
 sg13g2_fill_8 FILLER_0_21_672 ();
 sg13g2_fill_8 FILLER_0_21_680 ();
 sg13g2_fill_8 FILLER_0_21_688 ();
 sg13g2_fill_8 FILLER_0_21_696 ();
 sg13g2_fill_8 FILLER_0_21_704 ();
 sg13g2_fill_8 FILLER_0_21_712 ();
 sg13g2_fill_8 FILLER_0_21_720 ();
 sg13g2_fill_8 FILLER_0_21_728 ();
 sg13g2_fill_8 FILLER_0_21_736 ();
 sg13g2_fill_8 FILLER_0_21_744 ();
 sg13g2_fill_8 FILLER_0_21_752 ();
 sg13g2_fill_8 FILLER_0_21_760 ();
 sg13g2_fill_8 FILLER_0_21_768 ();
 sg13g2_fill_8 FILLER_0_21_776 ();
 sg13g2_fill_8 FILLER_0_21_784 ();
 sg13g2_fill_8 FILLER_0_21_792 ();
 sg13g2_fill_8 FILLER_0_21_800 ();
 sg13g2_fill_8 FILLER_0_21_808 ();
 sg13g2_fill_8 FILLER_0_21_816 ();
 sg13g2_fill_8 FILLER_0_21_824 ();
 sg13g2_fill_8 FILLER_0_21_832 ();
 sg13g2_fill_8 FILLER_0_21_840 ();
 sg13g2_fill_8 FILLER_0_21_848 ();
 sg13g2_fill_8 FILLER_0_21_856 ();
 sg13g2_fill_8 FILLER_0_21_864 ();
 sg13g2_fill_8 FILLER_0_21_872 ();
 sg13g2_fill_8 FILLER_0_21_880 ();
 sg13g2_fill_8 FILLER_0_21_888 ();
 sg13g2_fill_8 FILLER_0_21_896 ();
 sg13g2_fill_8 FILLER_0_21_904 ();
 sg13g2_fill_8 FILLER_0_21_912 ();
 sg13g2_fill_8 FILLER_0_21_920 ();
 sg13g2_fill_8 FILLER_0_21_928 ();
 sg13g2_fill_8 FILLER_0_21_936 ();
 sg13g2_fill_8 FILLER_0_21_944 ();
 sg13g2_fill_8 FILLER_0_21_952 ();
 sg13g2_fill_8 FILLER_0_21_960 ();
 sg13g2_fill_8 FILLER_0_21_968 ();
 sg13g2_fill_8 FILLER_0_21_976 ();
 sg13g2_fill_8 FILLER_0_21_984 ();
 sg13g2_fill_8 FILLER_0_21_992 ();
 sg13g2_fill_8 FILLER_0_21_1000 ();
 sg13g2_fill_8 FILLER_0_21_1008 ();
 sg13g2_fill_8 FILLER_0_21_1016 ();
 sg13g2_fill_8 FILLER_0_21_1024 ();
 sg13g2_fill_8 FILLER_0_21_1032 ();
 sg13g2_fill_8 FILLER_0_21_1040 ();
 sg13g2_fill_8 FILLER_0_21_1048 ();
 sg13g2_fill_8 FILLER_0_21_1056 ();
 sg13g2_fill_8 FILLER_0_21_1064 ();
 sg13g2_fill_8 FILLER_0_21_1072 ();
 sg13g2_fill_8 FILLER_0_21_1080 ();
 sg13g2_fill_8 FILLER_0_21_1088 ();
 sg13g2_fill_8 FILLER_0_21_1096 ();
 sg13g2_fill_8 FILLER_0_21_1104 ();
 sg13g2_fill_8 FILLER_0_21_1112 ();
 sg13g2_fill_8 FILLER_0_21_1120 ();
 sg13g2_fill_8 FILLER_0_21_1128 ();
 sg13g2_fill_8 FILLER_0_21_1136 ();
 sg13g2_fill_8 FILLER_0_21_1144 ();
 sg13g2_fill_8 FILLER_0_21_1152 ();
 sg13g2_fill_8 FILLER_0_21_1160 ();
 sg13g2_fill_8 FILLER_0_21_1168 ();
 sg13g2_fill_8 FILLER_0_21_1176 ();
 sg13g2_fill_8 FILLER_0_21_1184 ();
 sg13g2_fill_8 FILLER_0_21_1192 ();
 sg13g2_fill_8 FILLER_0_21_1200 ();
 sg13g2_fill_8 FILLER_0_21_1208 ();
 sg13g2_fill_8 FILLER_0_21_1216 ();
 sg13g2_fill_4 FILLER_0_21_1224 ();
 sg13g2_fill_8 FILLER_0_22_0 ();
 sg13g2_fill_8 FILLER_0_22_8 ();
 sg13g2_fill_8 FILLER_0_22_16 ();
 sg13g2_fill_8 FILLER_0_22_24 ();
 sg13g2_fill_8 FILLER_0_22_32 ();
 sg13g2_fill_8 FILLER_0_22_40 ();
 sg13g2_fill_8 FILLER_0_22_48 ();
 sg13g2_fill_8 FILLER_0_22_56 ();
 sg13g2_fill_8 FILLER_0_22_64 ();
 sg13g2_fill_8 FILLER_0_22_72 ();
 sg13g2_fill_8 FILLER_0_22_80 ();
 sg13g2_decap_8 FILLER_0_22_88 ();
 sg13g2_fill_8 FILLER_0_22_121 ();
 sg13g2_fill_8 FILLER_0_22_129 ();
 sg13g2_fill_8 FILLER_0_22_137 ();
 sg13g2_fill_8 FILLER_0_22_145 ();
 sg13g2_fill_8 FILLER_0_22_153 ();
 sg13g2_fill_2 FILLER_0_22_161 ();
 sg13g2_fill_1 FILLER_0_22_163 ();
 sg13g2_fill_8 FILLER_0_22_224 ();
 sg13g2_fill_8 FILLER_0_22_232 ();
 sg13g2_fill_8 FILLER_0_22_240 ();
 sg13g2_fill_2 FILLER_0_22_248 ();
 sg13g2_fill_1 FILLER_0_22_250 ();
 sg13g2_fill_1 FILLER_0_22_282 ();
 sg13g2_fill_1 FILLER_0_22_293 ();
 sg13g2_fill_4 FILLER_0_22_298 ();
 sg13g2_fill_2 FILLER_0_22_302 ();
 sg13g2_fill_4 FILLER_0_22_330 ();
 sg13g2_fill_1 FILLER_0_22_360 ();
 sg13g2_fill_1 FILLER_0_22_366 ();
 sg13g2_fill_1 FILLER_0_22_413 ();
 sg13g2_fill_8 FILLER_0_22_418 ();
 sg13g2_fill_8 FILLER_0_22_426 ();
 sg13g2_fill_8 FILLER_0_22_434 ();
 sg13g2_fill_8 FILLER_0_22_442 ();
 sg13g2_fill_8 FILLER_0_22_450 ();
 sg13g2_fill_8 FILLER_0_22_458 ();
 sg13g2_fill_8 FILLER_0_22_466 ();
 sg13g2_fill_8 FILLER_0_22_474 ();
 sg13g2_fill_8 FILLER_0_22_482 ();
 sg13g2_fill_8 FILLER_0_22_490 ();
 sg13g2_fill_8 FILLER_0_22_498 ();
 sg13g2_fill_8 FILLER_0_22_506 ();
 sg13g2_fill_8 FILLER_0_22_514 ();
 sg13g2_fill_8 FILLER_0_22_522 ();
 sg13g2_fill_8 FILLER_0_22_530 ();
 sg13g2_fill_8 FILLER_0_22_538 ();
 sg13g2_fill_8 FILLER_0_22_546 ();
 sg13g2_fill_8 FILLER_0_22_554 ();
 sg13g2_fill_8 FILLER_0_22_562 ();
 sg13g2_fill_8 FILLER_0_22_570 ();
 sg13g2_fill_8 FILLER_0_22_578 ();
 sg13g2_fill_8 FILLER_0_22_586 ();
 sg13g2_fill_8 FILLER_0_22_594 ();
 sg13g2_fill_8 FILLER_0_22_602 ();
 sg13g2_fill_8 FILLER_0_22_610 ();
 sg13g2_fill_8 FILLER_0_22_618 ();
 sg13g2_fill_8 FILLER_0_22_626 ();
 sg13g2_fill_8 FILLER_0_22_634 ();
 sg13g2_fill_8 FILLER_0_22_642 ();
 sg13g2_fill_8 FILLER_0_22_650 ();
 sg13g2_fill_8 FILLER_0_22_658 ();
 sg13g2_fill_8 FILLER_0_22_666 ();
 sg13g2_fill_8 FILLER_0_22_674 ();
 sg13g2_fill_8 FILLER_0_22_682 ();
 sg13g2_fill_8 FILLER_0_22_690 ();
 sg13g2_fill_8 FILLER_0_22_698 ();
 sg13g2_fill_8 FILLER_0_22_706 ();
 sg13g2_fill_8 FILLER_0_22_714 ();
 sg13g2_fill_8 FILLER_0_22_722 ();
 sg13g2_fill_8 FILLER_0_22_730 ();
 sg13g2_fill_8 FILLER_0_22_738 ();
 sg13g2_fill_8 FILLER_0_22_746 ();
 sg13g2_fill_8 FILLER_0_22_754 ();
 sg13g2_fill_8 FILLER_0_22_762 ();
 sg13g2_fill_8 FILLER_0_22_770 ();
 sg13g2_fill_8 FILLER_0_22_778 ();
 sg13g2_fill_8 FILLER_0_22_786 ();
 sg13g2_fill_8 FILLER_0_22_794 ();
 sg13g2_fill_8 FILLER_0_22_802 ();
 sg13g2_fill_8 FILLER_0_22_810 ();
 sg13g2_fill_8 FILLER_0_22_818 ();
 sg13g2_fill_8 FILLER_0_22_826 ();
 sg13g2_fill_8 FILLER_0_22_834 ();
 sg13g2_fill_8 FILLER_0_22_842 ();
 sg13g2_fill_8 FILLER_0_22_850 ();
 sg13g2_fill_8 FILLER_0_22_858 ();
 sg13g2_fill_8 FILLER_0_22_866 ();
 sg13g2_fill_8 FILLER_0_22_874 ();
 sg13g2_fill_8 FILLER_0_22_882 ();
 sg13g2_fill_8 FILLER_0_22_890 ();
 sg13g2_fill_8 FILLER_0_22_898 ();
 sg13g2_fill_8 FILLER_0_22_906 ();
 sg13g2_fill_8 FILLER_0_22_914 ();
 sg13g2_fill_8 FILLER_0_22_922 ();
 sg13g2_fill_8 FILLER_0_22_930 ();
 sg13g2_fill_8 FILLER_0_22_938 ();
 sg13g2_fill_8 FILLER_0_22_946 ();
 sg13g2_fill_8 FILLER_0_22_954 ();
 sg13g2_fill_8 FILLER_0_22_962 ();
 sg13g2_fill_8 FILLER_0_22_970 ();
 sg13g2_fill_8 FILLER_0_22_978 ();
 sg13g2_fill_8 FILLER_0_22_986 ();
 sg13g2_fill_8 FILLER_0_22_994 ();
 sg13g2_fill_8 FILLER_0_22_1002 ();
 sg13g2_fill_8 FILLER_0_22_1010 ();
 sg13g2_fill_8 FILLER_0_22_1018 ();
 sg13g2_fill_8 FILLER_0_22_1026 ();
 sg13g2_fill_8 FILLER_0_22_1034 ();
 sg13g2_fill_8 FILLER_0_22_1042 ();
 sg13g2_fill_8 FILLER_0_22_1050 ();
 sg13g2_fill_8 FILLER_0_22_1058 ();
 sg13g2_fill_8 FILLER_0_22_1066 ();
 sg13g2_fill_8 FILLER_0_22_1074 ();
 sg13g2_fill_8 FILLER_0_22_1082 ();
 sg13g2_fill_8 FILLER_0_22_1090 ();
 sg13g2_fill_8 FILLER_0_22_1098 ();
 sg13g2_fill_8 FILLER_0_22_1106 ();
 sg13g2_fill_8 FILLER_0_22_1114 ();
 sg13g2_fill_8 FILLER_0_22_1122 ();
 sg13g2_fill_8 FILLER_0_22_1130 ();
 sg13g2_fill_8 FILLER_0_22_1138 ();
 sg13g2_fill_8 FILLER_0_22_1146 ();
 sg13g2_fill_8 FILLER_0_22_1154 ();
 sg13g2_fill_8 FILLER_0_22_1162 ();
 sg13g2_fill_8 FILLER_0_22_1170 ();
 sg13g2_fill_8 FILLER_0_22_1178 ();
 sg13g2_fill_8 FILLER_0_22_1186 ();
 sg13g2_fill_8 FILLER_0_22_1194 ();
 sg13g2_fill_8 FILLER_0_22_1202 ();
 sg13g2_fill_8 FILLER_0_22_1210 ();
 sg13g2_fill_8 FILLER_0_22_1218 ();
 sg13g2_fill_2 FILLER_0_22_1226 ();
 sg13g2_fill_8 FILLER_0_23_0 ();
 sg13g2_fill_8 FILLER_0_23_8 ();
 sg13g2_fill_8 FILLER_0_23_16 ();
 sg13g2_fill_8 FILLER_0_23_24 ();
 sg13g2_fill_8 FILLER_0_23_36 ();
 sg13g2_fill_8 FILLER_0_23_44 ();
 sg13g2_fill_8 FILLER_0_23_52 ();
 sg13g2_fill_4 FILLER_0_23_60 ();
 sg13g2_fill_1 FILLER_0_23_64 ();
 sg13g2_fill_8 FILLER_0_23_69 ();
 sg13g2_fill_8 FILLER_0_23_77 ();
 sg13g2_fill_8 FILLER_0_23_90 ();
 sg13g2_fill_1 FILLER_0_23_98 ();
 sg13g2_fill_2 FILLER_0_23_103 ();
 sg13g2_fill_1 FILLER_0_23_115 ();
 sg13g2_fill_4 FILLER_0_23_125 ();
 sg13g2_fill_1 FILLER_0_23_129 ();
 sg13g2_fill_1 FILLER_0_23_135 ();
 sg13g2_fill_2 FILLER_0_23_162 ();
 sg13g2_fill_1 FILLER_0_23_190 ();
 sg13g2_fill_2 FILLER_0_23_201 ();
 sg13g2_fill_1 FILLER_0_23_203 ();
 sg13g2_fill_4 FILLER_0_23_235 ();
 sg13g2_fill_8 FILLER_0_23_243 ();
 sg13g2_fill_2 FILLER_0_23_251 ();
 sg13g2_fill_1 FILLER_0_23_309 ();
 sg13g2_fill_8 FILLER_0_23_429 ();
 sg13g2_fill_8 FILLER_0_23_437 ();
 sg13g2_fill_8 FILLER_0_23_445 ();
 sg13g2_fill_8 FILLER_0_23_453 ();
 sg13g2_fill_8 FILLER_0_23_461 ();
 sg13g2_fill_8 FILLER_0_23_469 ();
 sg13g2_fill_8 FILLER_0_23_477 ();
 sg13g2_fill_8 FILLER_0_23_485 ();
 sg13g2_fill_8 FILLER_0_23_493 ();
 sg13g2_fill_8 FILLER_0_23_501 ();
 sg13g2_fill_8 FILLER_0_23_509 ();
 sg13g2_fill_8 FILLER_0_23_517 ();
 sg13g2_fill_8 FILLER_0_23_525 ();
 sg13g2_fill_8 FILLER_0_23_533 ();
 sg13g2_fill_8 FILLER_0_23_541 ();
 sg13g2_fill_8 FILLER_0_23_549 ();
 sg13g2_fill_8 FILLER_0_23_557 ();
 sg13g2_fill_8 FILLER_0_23_565 ();
 sg13g2_fill_8 FILLER_0_23_573 ();
 sg13g2_fill_8 FILLER_0_23_581 ();
 sg13g2_fill_8 FILLER_0_23_589 ();
 sg13g2_fill_8 FILLER_0_23_597 ();
 sg13g2_fill_8 FILLER_0_23_605 ();
 sg13g2_fill_8 FILLER_0_23_613 ();
 sg13g2_fill_8 FILLER_0_23_621 ();
 sg13g2_fill_8 FILLER_0_23_629 ();
 sg13g2_fill_8 FILLER_0_23_637 ();
 sg13g2_fill_8 FILLER_0_23_645 ();
 sg13g2_fill_8 FILLER_0_23_653 ();
 sg13g2_fill_8 FILLER_0_23_661 ();
 sg13g2_fill_8 FILLER_0_23_669 ();
 sg13g2_fill_8 FILLER_0_23_677 ();
 sg13g2_fill_8 FILLER_0_23_685 ();
 sg13g2_fill_8 FILLER_0_23_693 ();
 sg13g2_fill_8 FILLER_0_23_701 ();
 sg13g2_fill_8 FILLER_0_23_709 ();
 sg13g2_fill_8 FILLER_0_23_717 ();
 sg13g2_fill_8 FILLER_0_23_725 ();
 sg13g2_fill_8 FILLER_0_23_733 ();
 sg13g2_fill_8 FILLER_0_23_741 ();
 sg13g2_fill_8 FILLER_0_23_749 ();
 sg13g2_fill_8 FILLER_0_23_757 ();
 sg13g2_fill_8 FILLER_0_23_765 ();
 sg13g2_fill_8 FILLER_0_23_773 ();
 sg13g2_fill_8 FILLER_0_23_781 ();
 sg13g2_fill_8 FILLER_0_23_789 ();
 sg13g2_fill_8 FILLER_0_23_797 ();
 sg13g2_fill_8 FILLER_0_23_805 ();
 sg13g2_fill_8 FILLER_0_23_813 ();
 sg13g2_fill_8 FILLER_0_23_821 ();
 sg13g2_fill_8 FILLER_0_23_829 ();
 sg13g2_fill_8 FILLER_0_23_837 ();
 sg13g2_fill_8 FILLER_0_23_845 ();
 sg13g2_fill_8 FILLER_0_23_853 ();
 sg13g2_fill_8 FILLER_0_23_861 ();
 sg13g2_fill_8 FILLER_0_23_869 ();
 sg13g2_fill_8 FILLER_0_23_877 ();
 sg13g2_fill_8 FILLER_0_23_885 ();
 sg13g2_fill_8 FILLER_0_23_893 ();
 sg13g2_fill_8 FILLER_0_23_901 ();
 sg13g2_fill_8 FILLER_0_23_909 ();
 sg13g2_fill_8 FILLER_0_23_917 ();
 sg13g2_fill_8 FILLER_0_23_925 ();
 sg13g2_fill_8 FILLER_0_23_933 ();
 sg13g2_fill_8 FILLER_0_23_941 ();
 sg13g2_fill_8 FILLER_0_23_949 ();
 sg13g2_fill_8 FILLER_0_23_957 ();
 sg13g2_fill_8 FILLER_0_23_965 ();
 sg13g2_fill_8 FILLER_0_23_973 ();
 sg13g2_fill_8 FILLER_0_23_981 ();
 sg13g2_fill_8 FILLER_0_23_989 ();
 sg13g2_fill_8 FILLER_0_23_997 ();
 sg13g2_fill_8 FILLER_0_23_1005 ();
 sg13g2_fill_8 FILLER_0_23_1013 ();
 sg13g2_fill_8 FILLER_0_23_1021 ();
 sg13g2_fill_8 FILLER_0_23_1029 ();
 sg13g2_fill_8 FILLER_0_23_1037 ();
 sg13g2_fill_8 FILLER_0_23_1045 ();
 sg13g2_fill_8 FILLER_0_23_1053 ();
 sg13g2_fill_8 FILLER_0_23_1061 ();
 sg13g2_fill_8 FILLER_0_23_1069 ();
 sg13g2_fill_8 FILLER_0_23_1077 ();
 sg13g2_fill_8 FILLER_0_23_1085 ();
 sg13g2_fill_8 FILLER_0_23_1093 ();
 sg13g2_fill_8 FILLER_0_23_1101 ();
 sg13g2_fill_8 FILLER_0_23_1109 ();
 sg13g2_fill_8 FILLER_0_23_1117 ();
 sg13g2_fill_8 FILLER_0_23_1125 ();
 sg13g2_fill_8 FILLER_0_23_1133 ();
 sg13g2_fill_8 FILLER_0_23_1141 ();
 sg13g2_fill_8 FILLER_0_23_1149 ();
 sg13g2_fill_8 FILLER_0_23_1157 ();
 sg13g2_fill_8 FILLER_0_23_1165 ();
 sg13g2_fill_8 FILLER_0_23_1173 ();
 sg13g2_fill_8 FILLER_0_23_1181 ();
 sg13g2_fill_8 FILLER_0_23_1189 ();
 sg13g2_fill_8 FILLER_0_23_1197 ();
 sg13g2_fill_8 FILLER_0_23_1205 ();
 sg13g2_fill_8 FILLER_0_23_1213 ();
 sg13g2_decap_8 FILLER_0_23_1221 ();
 sg13g2_fill_8 FILLER_0_24_0 ();
 sg13g2_decap_8 FILLER_0_24_8 ();
 sg13g2_fill_2 FILLER_0_24_51 ();
 sg13g2_fill_1 FILLER_0_24_84 ();
 sg13g2_fill_2 FILLER_0_24_111 ();
 sg13g2_fill_2 FILLER_0_24_139 ();
 sg13g2_fill_2 FILLER_0_24_199 ();
 sg13g2_fill_2 FILLER_0_24_205 ();
 sg13g2_fill_1 FILLER_0_24_207 ();
 sg13g2_fill_2 FILLER_0_24_218 ();
 sg13g2_fill_1 FILLER_0_24_220 ();
 sg13g2_fill_2 FILLER_0_24_231 ();
 sg13g2_fill_4 FILLER_0_24_259 ();
 sg13g2_fill_2 FILLER_0_24_318 ();
 sg13g2_fill_1 FILLER_0_24_320 ();
 sg13g2_fill_2 FILLER_0_24_356 ();
 sg13g2_fill_1 FILLER_0_24_358 ();
 sg13g2_fill_2 FILLER_0_24_395 ();
 sg13g2_fill_1 FILLER_0_24_397 ();
 sg13g2_fill_8 FILLER_0_24_434 ();
 sg13g2_fill_8 FILLER_0_24_442 ();
 sg13g2_fill_8 FILLER_0_24_450 ();
 sg13g2_fill_8 FILLER_0_24_458 ();
 sg13g2_fill_8 FILLER_0_24_466 ();
 sg13g2_fill_8 FILLER_0_24_474 ();
 sg13g2_fill_8 FILLER_0_24_482 ();
 sg13g2_fill_8 FILLER_0_24_490 ();
 sg13g2_fill_8 FILLER_0_24_498 ();
 sg13g2_fill_8 FILLER_0_24_506 ();
 sg13g2_fill_8 FILLER_0_24_514 ();
 sg13g2_fill_8 FILLER_0_24_522 ();
 sg13g2_fill_8 FILLER_0_24_530 ();
 sg13g2_fill_8 FILLER_0_24_538 ();
 sg13g2_fill_8 FILLER_0_24_546 ();
 sg13g2_fill_8 FILLER_0_24_554 ();
 sg13g2_fill_8 FILLER_0_24_562 ();
 sg13g2_fill_8 FILLER_0_24_570 ();
 sg13g2_fill_8 FILLER_0_24_578 ();
 sg13g2_fill_8 FILLER_0_24_586 ();
 sg13g2_fill_8 FILLER_0_24_594 ();
 sg13g2_fill_8 FILLER_0_24_602 ();
 sg13g2_fill_8 FILLER_0_24_610 ();
 sg13g2_fill_8 FILLER_0_24_618 ();
 sg13g2_fill_8 FILLER_0_24_626 ();
 sg13g2_fill_8 FILLER_0_24_634 ();
 sg13g2_fill_8 FILLER_0_24_642 ();
 sg13g2_fill_8 FILLER_0_24_650 ();
 sg13g2_fill_8 FILLER_0_24_658 ();
 sg13g2_fill_8 FILLER_0_24_666 ();
 sg13g2_fill_8 FILLER_0_24_674 ();
 sg13g2_fill_8 FILLER_0_24_682 ();
 sg13g2_fill_8 FILLER_0_24_690 ();
 sg13g2_fill_8 FILLER_0_24_698 ();
 sg13g2_fill_8 FILLER_0_24_706 ();
 sg13g2_fill_8 FILLER_0_24_714 ();
 sg13g2_fill_8 FILLER_0_24_722 ();
 sg13g2_fill_8 FILLER_0_24_730 ();
 sg13g2_fill_8 FILLER_0_24_738 ();
 sg13g2_fill_8 FILLER_0_24_746 ();
 sg13g2_fill_8 FILLER_0_24_754 ();
 sg13g2_fill_8 FILLER_0_24_762 ();
 sg13g2_fill_8 FILLER_0_24_770 ();
 sg13g2_fill_8 FILLER_0_24_778 ();
 sg13g2_fill_8 FILLER_0_24_786 ();
 sg13g2_fill_8 FILLER_0_24_794 ();
 sg13g2_fill_8 FILLER_0_24_802 ();
 sg13g2_fill_8 FILLER_0_24_810 ();
 sg13g2_fill_8 FILLER_0_24_818 ();
 sg13g2_fill_8 FILLER_0_24_826 ();
 sg13g2_fill_8 FILLER_0_24_834 ();
 sg13g2_fill_8 FILLER_0_24_842 ();
 sg13g2_fill_8 FILLER_0_24_850 ();
 sg13g2_fill_8 FILLER_0_24_858 ();
 sg13g2_fill_8 FILLER_0_24_866 ();
 sg13g2_fill_8 FILLER_0_24_874 ();
 sg13g2_fill_8 FILLER_0_24_882 ();
 sg13g2_fill_8 FILLER_0_24_890 ();
 sg13g2_fill_8 FILLER_0_24_898 ();
 sg13g2_fill_8 FILLER_0_24_906 ();
 sg13g2_fill_8 FILLER_0_24_914 ();
 sg13g2_fill_8 FILLER_0_24_922 ();
 sg13g2_fill_8 FILLER_0_24_930 ();
 sg13g2_fill_8 FILLER_0_24_938 ();
 sg13g2_fill_8 FILLER_0_24_946 ();
 sg13g2_fill_8 FILLER_0_24_954 ();
 sg13g2_fill_8 FILLER_0_24_962 ();
 sg13g2_fill_8 FILLER_0_24_970 ();
 sg13g2_fill_8 FILLER_0_24_978 ();
 sg13g2_fill_8 FILLER_0_24_986 ();
 sg13g2_fill_8 FILLER_0_24_994 ();
 sg13g2_fill_8 FILLER_0_24_1002 ();
 sg13g2_fill_8 FILLER_0_24_1010 ();
 sg13g2_fill_8 FILLER_0_24_1018 ();
 sg13g2_fill_8 FILLER_0_24_1026 ();
 sg13g2_fill_8 FILLER_0_24_1034 ();
 sg13g2_fill_8 FILLER_0_24_1042 ();
 sg13g2_fill_8 FILLER_0_24_1050 ();
 sg13g2_fill_8 FILLER_0_24_1058 ();
 sg13g2_fill_8 FILLER_0_24_1066 ();
 sg13g2_fill_8 FILLER_0_24_1074 ();
 sg13g2_fill_8 FILLER_0_24_1082 ();
 sg13g2_fill_8 FILLER_0_24_1090 ();
 sg13g2_fill_8 FILLER_0_24_1098 ();
 sg13g2_fill_8 FILLER_0_24_1106 ();
 sg13g2_fill_8 FILLER_0_24_1114 ();
 sg13g2_fill_8 FILLER_0_24_1122 ();
 sg13g2_fill_8 FILLER_0_24_1130 ();
 sg13g2_fill_8 FILLER_0_24_1138 ();
 sg13g2_fill_8 FILLER_0_24_1146 ();
 sg13g2_fill_8 FILLER_0_24_1154 ();
 sg13g2_fill_8 FILLER_0_24_1162 ();
 sg13g2_fill_8 FILLER_0_24_1170 ();
 sg13g2_fill_8 FILLER_0_24_1178 ();
 sg13g2_fill_8 FILLER_0_24_1186 ();
 sg13g2_fill_8 FILLER_0_24_1194 ();
 sg13g2_fill_8 FILLER_0_24_1202 ();
 sg13g2_fill_8 FILLER_0_24_1210 ();
 sg13g2_fill_8 FILLER_0_24_1218 ();
 sg13g2_fill_2 FILLER_0_24_1226 ();
 sg13g2_fill_1 FILLER_0_25_0 ();
 sg13g2_fill_2 FILLER_0_25_27 ();
 sg13g2_fill_1 FILLER_0_25_33 ();
 sg13g2_fill_2 FILLER_0_25_103 ();
 sg13g2_fill_1 FILLER_0_25_105 ();
 sg13g2_fill_2 FILLER_0_25_150 ();
 sg13g2_fill_8 FILLER_0_25_156 ();
 sg13g2_fill_2 FILLER_0_25_164 ();
 sg13g2_fill_1 FILLER_0_25_166 ();
 sg13g2_fill_8 FILLER_0_25_191 ();
 sg13g2_fill_8 FILLER_0_25_199 ();
 sg13g2_fill_8 FILLER_0_25_207 ();
 sg13g2_fill_2 FILLER_0_25_215 ();
 sg13g2_fill_1 FILLER_0_25_217 ();
 sg13g2_fill_1 FILLER_0_25_284 ();
 sg13g2_fill_2 FILLER_0_25_290 ();
 sg13g2_fill_1 FILLER_0_25_297 ();
 sg13g2_fill_1 FILLER_0_25_308 ();
 sg13g2_fill_1 FILLER_0_25_324 ();
 sg13g2_fill_4 FILLER_0_25_337 ();
 sg13g2_fill_4 FILLER_0_25_345 ();
 sg13g2_fill_1 FILLER_0_25_349 ();
 sg13g2_decap_8 FILLER_0_25_354 ();
 sg13g2_fill_8 FILLER_0_25_373 ();
 sg13g2_fill_2 FILLER_0_25_381 ();
 sg13g2_fill_2 FILLER_0_25_387 ();
 sg13g2_fill_4 FILLER_0_25_399 ();
 sg13g2_decap_8 FILLER_0_25_408 ();
 sg13g2_fill_8 FILLER_0_25_419 ();
 sg13g2_fill_8 FILLER_0_25_427 ();
 sg13g2_fill_8 FILLER_0_25_435 ();
 sg13g2_fill_8 FILLER_0_25_443 ();
 sg13g2_fill_8 FILLER_0_25_451 ();
 sg13g2_fill_8 FILLER_0_25_459 ();
 sg13g2_fill_8 FILLER_0_25_467 ();
 sg13g2_fill_8 FILLER_0_25_475 ();
 sg13g2_fill_8 FILLER_0_25_483 ();
 sg13g2_fill_8 FILLER_0_25_491 ();
 sg13g2_fill_8 FILLER_0_25_499 ();
 sg13g2_fill_2 FILLER_0_25_507 ();
 sg13g2_fill_1 FILLER_0_25_509 ();
 sg13g2_fill_8 FILLER_0_25_536 ();
 sg13g2_fill_8 FILLER_0_25_544 ();
 sg13g2_fill_8 FILLER_0_25_552 ();
 sg13g2_fill_8 FILLER_0_25_560 ();
 sg13g2_fill_8 FILLER_0_25_568 ();
 sg13g2_fill_8 FILLER_0_25_576 ();
 sg13g2_fill_8 FILLER_0_25_584 ();
 sg13g2_fill_8 FILLER_0_25_592 ();
 sg13g2_fill_8 FILLER_0_25_600 ();
 sg13g2_fill_8 FILLER_0_25_608 ();
 sg13g2_fill_8 FILLER_0_25_616 ();
 sg13g2_fill_8 FILLER_0_25_624 ();
 sg13g2_fill_8 FILLER_0_25_632 ();
 sg13g2_fill_8 FILLER_0_25_640 ();
 sg13g2_fill_8 FILLER_0_25_648 ();
 sg13g2_fill_8 FILLER_0_25_656 ();
 sg13g2_fill_8 FILLER_0_25_664 ();
 sg13g2_fill_8 FILLER_0_25_672 ();
 sg13g2_fill_8 FILLER_0_25_680 ();
 sg13g2_fill_8 FILLER_0_25_688 ();
 sg13g2_fill_8 FILLER_0_25_696 ();
 sg13g2_fill_8 FILLER_0_25_704 ();
 sg13g2_fill_8 FILLER_0_25_712 ();
 sg13g2_fill_8 FILLER_0_25_720 ();
 sg13g2_fill_8 FILLER_0_25_728 ();
 sg13g2_fill_8 FILLER_0_25_736 ();
 sg13g2_fill_8 FILLER_0_25_744 ();
 sg13g2_fill_8 FILLER_0_25_752 ();
 sg13g2_fill_8 FILLER_0_25_760 ();
 sg13g2_fill_8 FILLER_0_25_768 ();
 sg13g2_fill_8 FILLER_0_25_776 ();
 sg13g2_fill_8 FILLER_0_25_784 ();
 sg13g2_fill_8 FILLER_0_25_792 ();
 sg13g2_fill_8 FILLER_0_25_800 ();
 sg13g2_fill_8 FILLER_0_25_808 ();
 sg13g2_fill_8 FILLER_0_25_816 ();
 sg13g2_fill_8 FILLER_0_25_824 ();
 sg13g2_fill_8 FILLER_0_25_832 ();
 sg13g2_fill_8 FILLER_0_25_840 ();
 sg13g2_fill_8 FILLER_0_25_848 ();
 sg13g2_fill_8 FILLER_0_25_856 ();
 sg13g2_fill_8 FILLER_0_25_864 ();
 sg13g2_fill_8 FILLER_0_25_872 ();
 sg13g2_fill_8 FILLER_0_25_880 ();
 sg13g2_fill_8 FILLER_0_25_888 ();
 sg13g2_fill_8 FILLER_0_25_896 ();
 sg13g2_fill_8 FILLER_0_25_904 ();
 sg13g2_fill_8 FILLER_0_25_912 ();
 sg13g2_fill_8 FILLER_0_25_920 ();
 sg13g2_fill_8 FILLER_0_25_928 ();
 sg13g2_fill_8 FILLER_0_25_936 ();
 sg13g2_fill_8 FILLER_0_25_944 ();
 sg13g2_fill_8 FILLER_0_25_952 ();
 sg13g2_fill_8 FILLER_0_25_960 ();
 sg13g2_fill_8 FILLER_0_25_968 ();
 sg13g2_fill_8 FILLER_0_25_976 ();
 sg13g2_fill_8 FILLER_0_25_984 ();
 sg13g2_fill_8 FILLER_0_25_992 ();
 sg13g2_fill_8 FILLER_0_25_1000 ();
 sg13g2_fill_8 FILLER_0_25_1008 ();
 sg13g2_fill_8 FILLER_0_25_1016 ();
 sg13g2_fill_8 FILLER_0_25_1024 ();
 sg13g2_fill_8 FILLER_0_25_1032 ();
 sg13g2_fill_8 FILLER_0_25_1040 ();
 sg13g2_fill_8 FILLER_0_25_1048 ();
 sg13g2_fill_8 FILLER_0_25_1056 ();
 sg13g2_fill_8 FILLER_0_25_1064 ();
 sg13g2_fill_8 FILLER_0_25_1072 ();
 sg13g2_fill_8 FILLER_0_25_1080 ();
 sg13g2_fill_8 FILLER_0_25_1088 ();
 sg13g2_fill_8 FILLER_0_25_1096 ();
 sg13g2_fill_8 FILLER_0_25_1104 ();
 sg13g2_fill_8 FILLER_0_25_1112 ();
 sg13g2_fill_8 FILLER_0_25_1120 ();
 sg13g2_fill_8 FILLER_0_25_1128 ();
 sg13g2_fill_8 FILLER_0_25_1136 ();
 sg13g2_fill_8 FILLER_0_25_1144 ();
 sg13g2_fill_8 FILLER_0_25_1152 ();
 sg13g2_fill_8 FILLER_0_25_1160 ();
 sg13g2_fill_8 FILLER_0_25_1168 ();
 sg13g2_fill_8 FILLER_0_25_1176 ();
 sg13g2_fill_8 FILLER_0_25_1184 ();
 sg13g2_fill_8 FILLER_0_25_1192 ();
 sg13g2_fill_8 FILLER_0_25_1200 ();
 sg13g2_fill_8 FILLER_0_25_1208 ();
 sg13g2_fill_8 FILLER_0_25_1216 ();
 sg13g2_fill_4 FILLER_0_25_1224 ();
 sg13g2_fill_2 FILLER_0_26_5 ();
 sg13g2_fill_1 FILLER_0_26_11 ();
 sg13g2_fill_1 FILLER_0_26_22 ();
 sg13g2_fill_1 FILLER_0_26_28 ();
 sg13g2_fill_1 FILLER_0_26_54 ();
 sg13g2_fill_4 FILLER_0_26_80 ();
 sg13g2_fill_1 FILLER_0_26_84 ();
 sg13g2_fill_8 FILLER_0_26_119 ();
 sg13g2_decap_8 FILLER_0_26_127 ();
 sg13g2_fill_8 FILLER_0_26_144 ();
 sg13g2_fill_8 FILLER_0_26_152 ();
 sg13g2_fill_8 FILLER_0_26_160 ();
 sg13g2_fill_2 FILLER_0_26_194 ();
 sg13g2_fill_2 FILLER_0_26_222 ();
 sg13g2_fill_1 FILLER_0_26_224 ();
 sg13g2_fill_8 FILLER_0_26_252 ();
 sg13g2_fill_4 FILLER_0_26_260 ();
 sg13g2_fill_8 FILLER_0_26_279 ();
 sg13g2_fill_8 FILLER_0_26_287 ();
 sg13g2_decap_8 FILLER_0_26_295 ();
 sg13g2_fill_2 FILLER_0_26_310 ();
 sg13g2_fill_8 FILLER_0_26_316 ();
 sg13g2_fill_4 FILLER_0_26_329 ();
 sg13g2_fill_8 FILLER_0_26_337 ();
 sg13g2_fill_8 FILLER_0_26_345 ();
 sg13g2_fill_8 FILLER_0_26_353 ();
 sg13g2_fill_4 FILLER_0_26_361 ();
 sg13g2_fill_8 FILLER_0_26_373 ();
 sg13g2_fill_8 FILLER_0_26_381 ();
 sg13g2_fill_2 FILLER_0_26_389 ();
 sg13g2_fill_8 FILLER_0_26_431 ();
 sg13g2_fill_8 FILLER_0_26_439 ();
 sg13g2_fill_8 FILLER_0_26_447 ();
 sg13g2_fill_4 FILLER_0_26_455 ();
 sg13g2_fill_8 FILLER_0_26_467 ();
 sg13g2_fill_8 FILLER_0_26_475 ();
 sg13g2_fill_8 FILLER_0_26_483 ();
 sg13g2_fill_8 FILLER_0_26_491 ();
 sg13g2_fill_8 FILLER_0_26_499 ();
 sg13g2_fill_8 FILLER_0_26_507 ();
 sg13g2_fill_2 FILLER_0_26_515 ();
 sg13g2_fill_1 FILLER_0_26_517 ();
 sg13g2_fill_8 FILLER_0_26_567 ();
 sg13g2_fill_8 FILLER_0_26_575 ();
 sg13g2_fill_8 FILLER_0_26_583 ();
 sg13g2_fill_8 FILLER_0_26_591 ();
 sg13g2_fill_8 FILLER_0_26_599 ();
 sg13g2_fill_8 FILLER_0_26_607 ();
 sg13g2_fill_8 FILLER_0_26_615 ();
 sg13g2_fill_8 FILLER_0_26_623 ();
 sg13g2_fill_8 FILLER_0_26_631 ();
 sg13g2_fill_8 FILLER_0_26_639 ();
 sg13g2_fill_8 FILLER_0_26_647 ();
 sg13g2_fill_8 FILLER_0_26_655 ();
 sg13g2_fill_8 FILLER_0_26_663 ();
 sg13g2_fill_8 FILLER_0_26_671 ();
 sg13g2_fill_8 FILLER_0_26_679 ();
 sg13g2_fill_8 FILLER_0_26_687 ();
 sg13g2_fill_8 FILLER_0_26_695 ();
 sg13g2_fill_8 FILLER_0_26_703 ();
 sg13g2_fill_8 FILLER_0_26_711 ();
 sg13g2_fill_8 FILLER_0_26_719 ();
 sg13g2_fill_8 FILLER_0_26_727 ();
 sg13g2_fill_8 FILLER_0_26_735 ();
 sg13g2_fill_8 FILLER_0_26_743 ();
 sg13g2_fill_8 FILLER_0_26_751 ();
 sg13g2_fill_8 FILLER_0_26_759 ();
 sg13g2_fill_8 FILLER_0_26_767 ();
 sg13g2_fill_8 FILLER_0_26_775 ();
 sg13g2_fill_8 FILLER_0_26_783 ();
 sg13g2_fill_8 FILLER_0_26_791 ();
 sg13g2_fill_8 FILLER_0_26_799 ();
 sg13g2_fill_8 FILLER_0_26_807 ();
 sg13g2_fill_8 FILLER_0_26_815 ();
 sg13g2_fill_8 FILLER_0_26_823 ();
 sg13g2_fill_8 FILLER_0_26_831 ();
 sg13g2_fill_8 FILLER_0_26_839 ();
 sg13g2_fill_8 FILLER_0_26_847 ();
 sg13g2_fill_8 FILLER_0_26_855 ();
 sg13g2_fill_8 FILLER_0_26_863 ();
 sg13g2_fill_8 FILLER_0_26_871 ();
 sg13g2_fill_8 FILLER_0_26_879 ();
 sg13g2_fill_8 FILLER_0_26_887 ();
 sg13g2_fill_8 FILLER_0_26_895 ();
 sg13g2_fill_8 FILLER_0_26_903 ();
 sg13g2_fill_8 FILLER_0_26_911 ();
 sg13g2_fill_8 FILLER_0_26_919 ();
 sg13g2_fill_8 FILLER_0_26_927 ();
 sg13g2_fill_8 FILLER_0_26_935 ();
 sg13g2_fill_8 FILLER_0_26_943 ();
 sg13g2_fill_8 FILLER_0_26_951 ();
 sg13g2_fill_8 FILLER_0_26_959 ();
 sg13g2_fill_8 FILLER_0_26_967 ();
 sg13g2_fill_8 FILLER_0_26_975 ();
 sg13g2_fill_8 FILLER_0_26_983 ();
 sg13g2_fill_8 FILLER_0_26_991 ();
 sg13g2_fill_8 FILLER_0_26_999 ();
 sg13g2_fill_8 FILLER_0_26_1007 ();
 sg13g2_fill_8 FILLER_0_26_1015 ();
 sg13g2_fill_8 FILLER_0_26_1023 ();
 sg13g2_fill_8 FILLER_0_26_1031 ();
 sg13g2_fill_8 FILLER_0_26_1039 ();
 sg13g2_fill_8 FILLER_0_26_1047 ();
 sg13g2_fill_8 FILLER_0_26_1055 ();
 sg13g2_fill_8 FILLER_0_26_1063 ();
 sg13g2_fill_8 FILLER_0_26_1071 ();
 sg13g2_fill_8 FILLER_0_26_1079 ();
 sg13g2_fill_8 FILLER_0_26_1087 ();
 sg13g2_fill_8 FILLER_0_26_1095 ();
 sg13g2_fill_8 FILLER_0_26_1103 ();
 sg13g2_fill_8 FILLER_0_26_1111 ();
 sg13g2_fill_8 FILLER_0_26_1119 ();
 sg13g2_fill_8 FILLER_0_26_1127 ();
 sg13g2_fill_8 FILLER_0_26_1135 ();
 sg13g2_fill_8 FILLER_0_26_1143 ();
 sg13g2_fill_8 FILLER_0_26_1151 ();
 sg13g2_fill_8 FILLER_0_26_1159 ();
 sg13g2_fill_8 FILLER_0_26_1167 ();
 sg13g2_fill_8 FILLER_0_26_1175 ();
 sg13g2_fill_8 FILLER_0_26_1183 ();
 sg13g2_fill_8 FILLER_0_26_1191 ();
 sg13g2_fill_8 FILLER_0_26_1199 ();
 sg13g2_fill_8 FILLER_0_26_1207 ();
 sg13g2_fill_8 FILLER_0_26_1215 ();
 sg13g2_fill_4 FILLER_0_26_1223 ();
 sg13g2_fill_1 FILLER_0_26_1227 ();
 sg13g2_decap_8 FILLER_0_27_0 ();
 sg13g2_fill_4 FILLER_0_27_50 ();
 sg13g2_fill_1 FILLER_0_27_54 ();
 sg13g2_fill_4 FILLER_0_27_60 ();
 sg13g2_fill_4 FILLER_0_27_78 ();
 sg13g2_fill_1 FILLER_0_27_82 ();
 sg13g2_fill_8 FILLER_0_27_106 ();
 sg13g2_fill_8 FILLER_0_27_114 ();
 sg13g2_fill_4 FILLER_0_27_122 ();
 sg13g2_fill_1 FILLER_0_27_126 ();
 sg13g2_fill_4 FILLER_0_27_135 ();
 sg13g2_fill_8 FILLER_0_27_153 ();
 sg13g2_fill_4 FILLER_0_27_161 ();
 sg13g2_fill_2 FILLER_0_27_206 ();
 sg13g2_fill_8 FILLER_0_27_220 ();
 sg13g2_fill_8 FILLER_0_27_268 ();
 sg13g2_fill_4 FILLER_0_27_276 ();
 sg13g2_fill_1 FILLER_0_27_316 ();
 sg13g2_fill_1 FILLER_0_27_327 ();
 sg13g2_fill_2 FILLER_0_27_332 ();
 sg13g2_fill_2 FILLER_0_27_339 ();
 sg13g2_fill_2 FILLER_0_27_345 ();
 sg13g2_fill_1 FILLER_0_27_347 ();
 sg13g2_fill_1 FILLER_0_27_378 ();
 sg13g2_fill_2 FILLER_0_27_383 ();
 sg13g2_fill_1 FILLER_0_27_403 ();
 sg13g2_fill_8 FILLER_0_27_434 ();
 sg13g2_fill_8 FILLER_0_27_442 ();
 sg13g2_fill_8 FILLER_0_27_450 ();
 sg13g2_fill_8 FILLER_0_27_458 ();
 sg13g2_fill_8 FILLER_0_27_466 ();
 sg13g2_fill_8 FILLER_0_27_474 ();
 sg13g2_fill_8 FILLER_0_27_482 ();
 sg13g2_fill_8 FILLER_0_27_490 ();
 sg13g2_fill_1 FILLER_0_27_498 ();
 sg13g2_fill_2 FILLER_0_27_540 ();
 sg13g2_fill_1 FILLER_0_27_542 ();
 sg13g2_fill_8 FILLER_0_27_578 ();
 sg13g2_fill_8 FILLER_0_27_586 ();
 sg13g2_fill_8 FILLER_0_27_594 ();
 sg13g2_fill_8 FILLER_0_27_602 ();
 sg13g2_fill_8 FILLER_0_27_610 ();
 sg13g2_fill_8 FILLER_0_27_618 ();
 sg13g2_fill_8 FILLER_0_27_626 ();
 sg13g2_fill_8 FILLER_0_27_634 ();
 sg13g2_fill_8 FILLER_0_27_642 ();
 sg13g2_fill_8 FILLER_0_27_650 ();
 sg13g2_fill_8 FILLER_0_27_658 ();
 sg13g2_fill_8 FILLER_0_27_666 ();
 sg13g2_fill_8 FILLER_0_27_674 ();
 sg13g2_fill_8 FILLER_0_27_682 ();
 sg13g2_fill_8 FILLER_0_27_690 ();
 sg13g2_fill_8 FILLER_0_27_698 ();
 sg13g2_fill_8 FILLER_0_27_706 ();
 sg13g2_fill_8 FILLER_0_27_714 ();
 sg13g2_fill_8 FILLER_0_27_722 ();
 sg13g2_fill_8 FILLER_0_27_730 ();
 sg13g2_fill_8 FILLER_0_27_738 ();
 sg13g2_fill_8 FILLER_0_27_746 ();
 sg13g2_fill_8 FILLER_0_27_754 ();
 sg13g2_fill_8 FILLER_0_27_762 ();
 sg13g2_fill_8 FILLER_0_27_770 ();
 sg13g2_fill_8 FILLER_0_27_778 ();
 sg13g2_fill_8 FILLER_0_27_786 ();
 sg13g2_fill_8 FILLER_0_27_794 ();
 sg13g2_fill_8 FILLER_0_27_802 ();
 sg13g2_fill_8 FILLER_0_27_810 ();
 sg13g2_fill_8 FILLER_0_27_818 ();
 sg13g2_fill_8 FILLER_0_27_826 ();
 sg13g2_fill_8 FILLER_0_27_834 ();
 sg13g2_fill_8 FILLER_0_27_842 ();
 sg13g2_fill_8 FILLER_0_27_850 ();
 sg13g2_fill_8 FILLER_0_27_858 ();
 sg13g2_fill_8 FILLER_0_27_866 ();
 sg13g2_fill_8 FILLER_0_27_874 ();
 sg13g2_fill_8 FILLER_0_27_882 ();
 sg13g2_fill_8 FILLER_0_27_890 ();
 sg13g2_fill_8 FILLER_0_27_898 ();
 sg13g2_fill_8 FILLER_0_27_906 ();
 sg13g2_fill_8 FILLER_0_27_914 ();
 sg13g2_fill_8 FILLER_0_27_922 ();
 sg13g2_fill_8 FILLER_0_27_930 ();
 sg13g2_fill_8 FILLER_0_27_938 ();
 sg13g2_fill_8 FILLER_0_27_946 ();
 sg13g2_fill_8 FILLER_0_27_954 ();
 sg13g2_fill_8 FILLER_0_27_962 ();
 sg13g2_fill_8 FILLER_0_27_970 ();
 sg13g2_fill_8 FILLER_0_27_978 ();
 sg13g2_fill_8 FILLER_0_27_986 ();
 sg13g2_fill_8 FILLER_0_27_994 ();
 sg13g2_fill_8 FILLER_0_27_1002 ();
 sg13g2_fill_8 FILLER_0_27_1010 ();
 sg13g2_fill_8 FILLER_0_27_1018 ();
 sg13g2_fill_8 FILLER_0_27_1026 ();
 sg13g2_fill_8 FILLER_0_27_1034 ();
 sg13g2_fill_8 FILLER_0_27_1042 ();
 sg13g2_fill_8 FILLER_0_27_1050 ();
 sg13g2_fill_8 FILLER_0_27_1058 ();
 sg13g2_fill_8 FILLER_0_27_1066 ();
 sg13g2_fill_8 FILLER_0_27_1074 ();
 sg13g2_fill_8 FILLER_0_27_1082 ();
 sg13g2_fill_8 FILLER_0_27_1090 ();
 sg13g2_fill_8 FILLER_0_27_1098 ();
 sg13g2_fill_8 FILLER_0_27_1106 ();
 sg13g2_fill_8 FILLER_0_27_1114 ();
 sg13g2_fill_8 FILLER_0_27_1122 ();
 sg13g2_fill_8 FILLER_0_27_1130 ();
 sg13g2_fill_8 FILLER_0_27_1138 ();
 sg13g2_fill_8 FILLER_0_27_1146 ();
 sg13g2_fill_8 FILLER_0_27_1154 ();
 sg13g2_fill_8 FILLER_0_27_1162 ();
 sg13g2_fill_8 FILLER_0_27_1170 ();
 sg13g2_fill_8 FILLER_0_27_1178 ();
 sg13g2_fill_8 FILLER_0_27_1186 ();
 sg13g2_fill_8 FILLER_0_27_1194 ();
 sg13g2_fill_8 FILLER_0_27_1202 ();
 sg13g2_fill_8 FILLER_0_27_1210 ();
 sg13g2_fill_8 FILLER_0_27_1218 ();
 sg13g2_fill_2 FILLER_0_27_1226 ();
 sg13g2_fill_8 FILLER_0_28_0 ();
 sg13g2_decap_8 FILLER_0_28_8 ();
 sg13g2_fill_8 FILLER_0_28_19 ();
 sg13g2_fill_2 FILLER_0_28_27 ();
 sg13g2_fill_8 FILLER_0_28_39 ();
 sg13g2_decap_8 FILLER_0_28_47 ();
 sg13g2_fill_2 FILLER_0_28_80 ();
 sg13g2_fill_4 FILLER_0_28_87 ();
 sg13g2_fill_4 FILLER_0_28_95 ();
 sg13g2_fill_2 FILLER_0_28_125 ();
 sg13g2_fill_1 FILLER_0_28_127 ();
 sg13g2_fill_8 FILLER_0_28_164 ();
 sg13g2_decap_8 FILLER_0_28_172 ();
 sg13g2_fill_8 FILLER_0_28_183 ();
 sg13g2_fill_8 FILLER_0_28_191 ();
 sg13g2_fill_8 FILLER_0_28_199 ();
 sg13g2_fill_8 FILLER_0_28_207 ();
 sg13g2_fill_8 FILLER_0_28_215 ();
 sg13g2_decap_8 FILLER_0_28_223 ();
 sg13g2_fill_2 FILLER_0_28_245 ();
 sg13g2_fill_2 FILLER_0_28_281 ();
 sg13g2_fill_2 FILLER_0_28_293 ();
 sg13g2_fill_1 FILLER_0_28_295 ();
 sg13g2_fill_4 FILLER_0_28_300 ();
 sg13g2_fill_8 FILLER_0_28_426 ();
 sg13g2_fill_8 FILLER_0_28_434 ();
 sg13g2_fill_8 FILLER_0_28_442 ();
 sg13g2_fill_8 FILLER_0_28_450 ();
 sg13g2_fill_8 FILLER_0_28_458 ();
 sg13g2_fill_8 FILLER_0_28_466 ();
 sg13g2_fill_8 FILLER_0_28_474 ();
 sg13g2_fill_8 FILLER_0_28_482 ();
 sg13g2_fill_8 FILLER_0_28_490 ();
 sg13g2_fill_8 FILLER_0_28_498 ();
 sg13g2_fill_2 FILLER_0_28_506 ();
 sg13g2_fill_1 FILLER_0_28_508 ();
 sg13g2_fill_1 FILLER_0_28_538 ();
 sg13g2_fill_1 FILLER_0_28_543 ();
 sg13g2_fill_1 FILLER_0_28_559 ();
 sg13g2_fill_8 FILLER_0_28_586 ();
 sg13g2_fill_8 FILLER_0_28_594 ();
 sg13g2_fill_8 FILLER_0_28_602 ();
 sg13g2_fill_8 FILLER_0_28_610 ();
 sg13g2_fill_8 FILLER_0_28_618 ();
 sg13g2_fill_8 FILLER_0_28_626 ();
 sg13g2_fill_8 FILLER_0_28_634 ();
 sg13g2_fill_8 FILLER_0_28_642 ();
 sg13g2_fill_8 FILLER_0_28_650 ();
 sg13g2_fill_8 FILLER_0_28_658 ();
 sg13g2_fill_8 FILLER_0_28_666 ();
 sg13g2_fill_8 FILLER_0_28_674 ();
 sg13g2_fill_8 FILLER_0_28_682 ();
 sg13g2_fill_8 FILLER_0_28_690 ();
 sg13g2_fill_8 FILLER_0_28_698 ();
 sg13g2_fill_8 FILLER_0_28_706 ();
 sg13g2_fill_8 FILLER_0_28_714 ();
 sg13g2_fill_8 FILLER_0_28_722 ();
 sg13g2_fill_8 FILLER_0_28_730 ();
 sg13g2_fill_8 FILLER_0_28_738 ();
 sg13g2_fill_8 FILLER_0_28_746 ();
 sg13g2_fill_8 FILLER_0_28_754 ();
 sg13g2_fill_8 FILLER_0_28_762 ();
 sg13g2_fill_8 FILLER_0_28_770 ();
 sg13g2_fill_8 FILLER_0_28_778 ();
 sg13g2_fill_8 FILLER_0_28_786 ();
 sg13g2_fill_8 FILLER_0_28_794 ();
 sg13g2_fill_8 FILLER_0_28_802 ();
 sg13g2_fill_8 FILLER_0_28_810 ();
 sg13g2_fill_8 FILLER_0_28_818 ();
 sg13g2_fill_8 FILLER_0_28_826 ();
 sg13g2_fill_8 FILLER_0_28_834 ();
 sg13g2_fill_8 FILLER_0_28_842 ();
 sg13g2_fill_8 FILLER_0_28_850 ();
 sg13g2_fill_8 FILLER_0_28_858 ();
 sg13g2_fill_8 FILLER_0_28_866 ();
 sg13g2_fill_8 FILLER_0_28_874 ();
 sg13g2_fill_8 FILLER_0_28_882 ();
 sg13g2_fill_8 FILLER_0_28_890 ();
 sg13g2_fill_8 FILLER_0_28_898 ();
 sg13g2_fill_8 FILLER_0_28_906 ();
 sg13g2_fill_8 FILLER_0_28_914 ();
 sg13g2_fill_8 FILLER_0_28_922 ();
 sg13g2_fill_8 FILLER_0_28_930 ();
 sg13g2_fill_8 FILLER_0_28_938 ();
 sg13g2_fill_8 FILLER_0_28_946 ();
 sg13g2_fill_8 FILLER_0_28_954 ();
 sg13g2_fill_8 FILLER_0_28_962 ();
 sg13g2_fill_8 FILLER_0_28_970 ();
 sg13g2_fill_8 FILLER_0_28_978 ();
 sg13g2_fill_8 FILLER_0_28_986 ();
 sg13g2_fill_8 FILLER_0_28_994 ();
 sg13g2_fill_8 FILLER_0_28_1002 ();
 sg13g2_fill_8 FILLER_0_28_1010 ();
 sg13g2_fill_8 FILLER_0_28_1018 ();
 sg13g2_fill_8 FILLER_0_28_1026 ();
 sg13g2_fill_8 FILLER_0_28_1034 ();
 sg13g2_fill_8 FILLER_0_28_1042 ();
 sg13g2_fill_8 FILLER_0_28_1050 ();
 sg13g2_fill_8 FILLER_0_28_1058 ();
 sg13g2_fill_8 FILLER_0_28_1066 ();
 sg13g2_fill_8 FILLER_0_28_1074 ();
 sg13g2_fill_8 FILLER_0_28_1082 ();
 sg13g2_fill_8 FILLER_0_28_1090 ();
 sg13g2_fill_8 FILLER_0_28_1098 ();
 sg13g2_fill_8 FILLER_0_28_1106 ();
 sg13g2_fill_8 FILLER_0_28_1114 ();
 sg13g2_fill_8 FILLER_0_28_1122 ();
 sg13g2_fill_8 FILLER_0_28_1130 ();
 sg13g2_fill_8 FILLER_0_28_1138 ();
 sg13g2_fill_8 FILLER_0_28_1146 ();
 sg13g2_fill_8 FILLER_0_28_1154 ();
 sg13g2_fill_8 FILLER_0_28_1162 ();
 sg13g2_fill_8 FILLER_0_28_1170 ();
 sg13g2_fill_8 FILLER_0_28_1178 ();
 sg13g2_fill_8 FILLER_0_28_1186 ();
 sg13g2_fill_8 FILLER_0_28_1194 ();
 sg13g2_fill_8 FILLER_0_28_1202 ();
 sg13g2_fill_8 FILLER_0_28_1210 ();
 sg13g2_fill_8 FILLER_0_28_1218 ();
 sg13g2_fill_2 FILLER_0_28_1226 ();
 sg13g2_fill_8 FILLER_0_29_0 ();
 sg13g2_fill_1 FILLER_0_29_39 ();
 sg13g2_fill_1 FILLER_0_29_44 ();
 sg13g2_fill_2 FILLER_0_29_53 ();
 sg13g2_fill_2 FILLER_0_29_81 ();
 sg13g2_fill_1 FILLER_0_29_83 ();
 sg13g2_fill_2 FILLER_0_29_172 ();
 sg13g2_fill_1 FILLER_0_29_174 ();
 sg13g2_fill_1 FILLER_0_29_205 ();
 sg13g2_fill_2 FILLER_0_29_232 ();
 sg13g2_fill_2 FILLER_0_29_274 ();
 sg13g2_fill_1 FILLER_0_29_276 ();
 sg13g2_fill_2 FILLER_0_29_287 ();
 sg13g2_fill_4 FILLER_0_29_298 ();
 sg13g2_fill_2 FILLER_0_29_302 ();
 sg13g2_fill_4 FILLER_0_29_308 ();
 sg13g2_fill_1 FILLER_0_29_312 ();
 sg13g2_fill_2 FILLER_0_29_347 ();
 sg13g2_fill_1 FILLER_0_29_349 ();
 sg13g2_fill_1 FILLER_0_29_354 ();
 sg13g2_fill_1 FILLER_0_29_360 ();
 sg13g2_fill_2 FILLER_0_29_366 ();
 sg13g2_fill_1 FILLER_0_29_378 ();
 sg13g2_fill_8 FILLER_0_29_420 ();
 sg13g2_fill_4 FILLER_0_29_428 ();
 sg13g2_fill_2 FILLER_0_29_432 ();
 sg13g2_fill_4 FILLER_0_29_438 ();
 sg13g2_fill_8 FILLER_0_29_452 ();
 sg13g2_fill_2 FILLER_0_29_460 ();
 sg13g2_decap_8 FILLER_0_29_466 ();
 sg13g2_fill_8 FILLER_0_29_482 ();
 sg13g2_fill_8 FILLER_0_29_490 ();
 sg13g2_fill_8 FILLER_0_29_498 ();
 sg13g2_decap_8 FILLER_0_29_506 ();
 sg13g2_fill_8 FILLER_0_29_536 ();
 sg13g2_fill_4 FILLER_0_29_544 ();
 sg13g2_fill_2 FILLER_0_29_548 ();
 sg13g2_fill_8 FILLER_0_29_586 ();
 sg13g2_fill_8 FILLER_0_29_594 ();
 sg13g2_fill_8 FILLER_0_29_602 ();
 sg13g2_fill_8 FILLER_0_29_610 ();
 sg13g2_fill_8 FILLER_0_29_618 ();
 sg13g2_fill_8 FILLER_0_29_626 ();
 sg13g2_fill_8 FILLER_0_29_634 ();
 sg13g2_fill_8 FILLER_0_29_642 ();
 sg13g2_fill_8 FILLER_0_29_650 ();
 sg13g2_fill_8 FILLER_0_29_658 ();
 sg13g2_fill_8 FILLER_0_29_666 ();
 sg13g2_fill_8 FILLER_0_29_674 ();
 sg13g2_fill_8 FILLER_0_29_682 ();
 sg13g2_fill_8 FILLER_0_29_690 ();
 sg13g2_fill_8 FILLER_0_29_698 ();
 sg13g2_fill_8 FILLER_0_29_706 ();
 sg13g2_fill_8 FILLER_0_29_714 ();
 sg13g2_fill_8 FILLER_0_29_722 ();
 sg13g2_fill_8 FILLER_0_29_730 ();
 sg13g2_fill_8 FILLER_0_29_738 ();
 sg13g2_fill_8 FILLER_0_29_746 ();
 sg13g2_fill_8 FILLER_0_29_754 ();
 sg13g2_fill_8 FILLER_0_29_762 ();
 sg13g2_fill_8 FILLER_0_29_770 ();
 sg13g2_fill_8 FILLER_0_29_778 ();
 sg13g2_fill_8 FILLER_0_29_786 ();
 sg13g2_fill_8 FILLER_0_29_794 ();
 sg13g2_fill_8 FILLER_0_29_802 ();
 sg13g2_fill_8 FILLER_0_29_810 ();
 sg13g2_fill_8 FILLER_0_29_818 ();
 sg13g2_fill_8 FILLER_0_29_826 ();
 sg13g2_fill_8 FILLER_0_29_834 ();
 sg13g2_fill_8 FILLER_0_29_842 ();
 sg13g2_fill_8 FILLER_0_29_850 ();
 sg13g2_fill_8 FILLER_0_29_858 ();
 sg13g2_fill_8 FILLER_0_29_866 ();
 sg13g2_fill_8 FILLER_0_29_874 ();
 sg13g2_fill_8 FILLER_0_29_882 ();
 sg13g2_fill_8 FILLER_0_29_890 ();
 sg13g2_fill_8 FILLER_0_29_898 ();
 sg13g2_fill_8 FILLER_0_29_906 ();
 sg13g2_fill_8 FILLER_0_29_914 ();
 sg13g2_fill_8 FILLER_0_29_922 ();
 sg13g2_fill_8 FILLER_0_29_930 ();
 sg13g2_fill_8 FILLER_0_29_938 ();
 sg13g2_fill_8 FILLER_0_29_946 ();
 sg13g2_fill_8 FILLER_0_29_954 ();
 sg13g2_fill_8 FILLER_0_29_962 ();
 sg13g2_fill_8 FILLER_0_29_970 ();
 sg13g2_fill_8 FILLER_0_29_978 ();
 sg13g2_fill_8 FILLER_0_29_986 ();
 sg13g2_fill_8 FILLER_0_29_994 ();
 sg13g2_fill_8 FILLER_0_29_1002 ();
 sg13g2_fill_8 FILLER_0_29_1010 ();
 sg13g2_fill_8 FILLER_0_29_1018 ();
 sg13g2_fill_8 FILLER_0_29_1026 ();
 sg13g2_fill_8 FILLER_0_29_1034 ();
 sg13g2_fill_8 FILLER_0_29_1042 ();
 sg13g2_fill_8 FILLER_0_29_1050 ();
 sg13g2_fill_8 FILLER_0_29_1058 ();
 sg13g2_fill_8 FILLER_0_29_1066 ();
 sg13g2_fill_8 FILLER_0_29_1074 ();
 sg13g2_fill_8 FILLER_0_29_1082 ();
 sg13g2_fill_8 FILLER_0_29_1090 ();
 sg13g2_fill_8 FILLER_0_29_1098 ();
 sg13g2_fill_8 FILLER_0_29_1106 ();
 sg13g2_fill_8 FILLER_0_29_1114 ();
 sg13g2_fill_8 FILLER_0_29_1122 ();
 sg13g2_fill_8 FILLER_0_29_1130 ();
 sg13g2_fill_8 FILLER_0_29_1138 ();
 sg13g2_fill_8 FILLER_0_29_1146 ();
 sg13g2_fill_8 FILLER_0_29_1154 ();
 sg13g2_fill_8 FILLER_0_29_1162 ();
 sg13g2_fill_8 FILLER_0_29_1170 ();
 sg13g2_fill_8 FILLER_0_29_1178 ();
 sg13g2_fill_8 FILLER_0_29_1186 ();
 sg13g2_fill_8 FILLER_0_29_1194 ();
 sg13g2_fill_8 FILLER_0_29_1202 ();
 sg13g2_fill_8 FILLER_0_29_1210 ();
 sg13g2_fill_8 FILLER_0_29_1218 ();
 sg13g2_fill_2 FILLER_0_29_1226 ();
 sg13g2_fill_1 FILLER_0_30_0 ();
 sg13g2_fill_1 FILLER_0_30_5 ();
 sg13g2_fill_2 FILLER_0_30_67 ();
 sg13g2_fill_1 FILLER_0_30_79 ();
 sg13g2_fill_1 FILLER_0_30_90 ();
 sg13g2_fill_1 FILLER_0_30_95 ();
 sg13g2_fill_2 FILLER_0_30_106 ();
 sg13g2_decap_8 FILLER_0_30_112 ();
 sg13g2_fill_4 FILLER_0_30_123 ();
 sg13g2_decap_8 FILLER_0_30_147 ();
 sg13g2_fill_4 FILLER_0_30_158 ();
 sg13g2_fill_8 FILLER_0_30_203 ();
 sg13g2_fill_4 FILLER_0_30_211 ();
 sg13g2_fill_4 FILLER_0_30_223 ();
 sg13g2_fill_2 FILLER_0_30_227 ();
 sg13g2_fill_8 FILLER_0_30_244 ();
 sg13g2_fill_4 FILLER_0_30_252 ();
 sg13g2_fill_2 FILLER_0_30_256 ();
 sg13g2_fill_4 FILLER_0_30_281 ();
 sg13g2_fill_1 FILLER_0_30_285 ();
 sg13g2_fill_2 FILLER_0_30_322 ();
 sg13g2_fill_4 FILLER_0_30_338 ();
 sg13g2_fill_2 FILLER_0_30_368 ();
 sg13g2_fill_1 FILLER_0_30_370 ();
 sg13g2_fill_8 FILLER_0_30_375 ();
 sg13g2_fill_4 FILLER_0_30_383 ();
 sg13g2_fill_2 FILLER_0_30_387 ();
 sg13g2_fill_4 FILLER_0_30_394 ();
 sg13g2_fill_2 FILLER_0_30_398 ();
 sg13g2_fill_4 FILLER_0_30_404 ();
 sg13g2_fill_8 FILLER_0_30_412 ();
 sg13g2_fill_4 FILLER_0_30_420 ();
 sg13g2_fill_2 FILLER_0_30_424 ();
 sg13g2_fill_2 FILLER_0_30_462 ();
 sg13g2_fill_1 FILLER_0_30_464 ();
 sg13g2_fill_8 FILLER_0_30_496 ();
 sg13g2_fill_2 FILLER_0_30_504 ();
 sg13g2_fill_2 FILLER_0_30_541 ();
 sg13g2_fill_4 FILLER_0_30_557 ();
 sg13g2_fill_1 FILLER_0_30_566 ();
 sg13g2_fill_8 FILLER_0_30_571 ();
 sg13g2_fill_8 FILLER_0_30_579 ();
 sg13g2_fill_8 FILLER_0_30_587 ();
 sg13g2_fill_8 FILLER_0_30_595 ();
 sg13g2_fill_8 FILLER_0_30_603 ();
 sg13g2_fill_8 FILLER_0_30_611 ();
 sg13g2_fill_8 FILLER_0_30_619 ();
 sg13g2_fill_8 FILLER_0_30_627 ();
 sg13g2_fill_8 FILLER_0_30_635 ();
 sg13g2_fill_8 FILLER_0_30_643 ();
 sg13g2_fill_8 FILLER_0_30_651 ();
 sg13g2_fill_8 FILLER_0_30_659 ();
 sg13g2_fill_8 FILLER_0_30_667 ();
 sg13g2_fill_8 FILLER_0_30_675 ();
 sg13g2_fill_8 FILLER_0_30_683 ();
 sg13g2_fill_8 FILLER_0_30_691 ();
 sg13g2_fill_8 FILLER_0_30_699 ();
 sg13g2_fill_8 FILLER_0_30_707 ();
 sg13g2_fill_8 FILLER_0_30_715 ();
 sg13g2_fill_8 FILLER_0_30_723 ();
 sg13g2_fill_8 FILLER_0_30_731 ();
 sg13g2_fill_8 FILLER_0_30_739 ();
 sg13g2_fill_8 FILLER_0_30_747 ();
 sg13g2_fill_8 FILLER_0_30_755 ();
 sg13g2_fill_8 FILLER_0_30_763 ();
 sg13g2_fill_8 FILLER_0_30_771 ();
 sg13g2_fill_8 FILLER_0_30_779 ();
 sg13g2_fill_8 FILLER_0_30_787 ();
 sg13g2_fill_8 FILLER_0_30_795 ();
 sg13g2_fill_8 FILLER_0_30_803 ();
 sg13g2_fill_8 FILLER_0_30_811 ();
 sg13g2_fill_8 FILLER_0_30_819 ();
 sg13g2_fill_8 FILLER_0_30_827 ();
 sg13g2_fill_8 FILLER_0_30_835 ();
 sg13g2_fill_8 FILLER_0_30_843 ();
 sg13g2_fill_8 FILLER_0_30_851 ();
 sg13g2_fill_8 FILLER_0_30_859 ();
 sg13g2_fill_8 FILLER_0_30_867 ();
 sg13g2_fill_8 FILLER_0_30_875 ();
 sg13g2_fill_8 FILLER_0_30_883 ();
 sg13g2_fill_8 FILLER_0_30_891 ();
 sg13g2_fill_8 FILLER_0_30_899 ();
 sg13g2_fill_8 FILLER_0_30_907 ();
 sg13g2_fill_8 FILLER_0_30_915 ();
 sg13g2_fill_8 FILLER_0_30_923 ();
 sg13g2_fill_8 FILLER_0_30_931 ();
 sg13g2_fill_8 FILLER_0_30_939 ();
 sg13g2_fill_8 FILLER_0_30_947 ();
 sg13g2_fill_8 FILLER_0_30_955 ();
 sg13g2_fill_8 FILLER_0_30_963 ();
 sg13g2_fill_8 FILLER_0_30_971 ();
 sg13g2_fill_8 FILLER_0_30_979 ();
 sg13g2_fill_8 FILLER_0_30_987 ();
 sg13g2_fill_8 FILLER_0_30_995 ();
 sg13g2_fill_8 FILLER_0_30_1003 ();
 sg13g2_fill_8 FILLER_0_30_1011 ();
 sg13g2_fill_8 FILLER_0_30_1019 ();
 sg13g2_fill_8 FILLER_0_30_1027 ();
 sg13g2_fill_8 FILLER_0_30_1035 ();
 sg13g2_fill_8 FILLER_0_30_1043 ();
 sg13g2_fill_8 FILLER_0_30_1051 ();
 sg13g2_fill_8 FILLER_0_30_1059 ();
 sg13g2_fill_8 FILLER_0_30_1067 ();
 sg13g2_fill_8 FILLER_0_30_1075 ();
 sg13g2_fill_8 FILLER_0_30_1083 ();
 sg13g2_fill_8 FILLER_0_30_1091 ();
 sg13g2_fill_8 FILLER_0_30_1099 ();
 sg13g2_fill_8 FILLER_0_30_1107 ();
 sg13g2_fill_8 FILLER_0_30_1115 ();
 sg13g2_fill_8 FILLER_0_30_1123 ();
 sg13g2_fill_8 FILLER_0_30_1131 ();
 sg13g2_fill_8 FILLER_0_30_1139 ();
 sg13g2_fill_8 FILLER_0_30_1147 ();
 sg13g2_fill_8 FILLER_0_30_1155 ();
 sg13g2_fill_8 FILLER_0_30_1163 ();
 sg13g2_fill_8 FILLER_0_30_1171 ();
 sg13g2_fill_8 FILLER_0_30_1179 ();
 sg13g2_fill_8 FILLER_0_30_1187 ();
 sg13g2_fill_8 FILLER_0_30_1195 ();
 sg13g2_fill_8 FILLER_0_30_1203 ();
 sg13g2_fill_8 FILLER_0_30_1211 ();
 sg13g2_fill_8 FILLER_0_30_1219 ();
 sg13g2_fill_1 FILLER_0_30_1227 ();
 sg13g2_fill_2 FILLER_0_31_0 ();
 sg13g2_fill_1 FILLER_0_31_28 ();
 sg13g2_fill_8 FILLER_0_31_73 ();
 sg13g2_fill_8 FILLER_0_31_81 ();
 sg13g2_fill_4 FILLER_0_31_89 ();
 sg13g2_fill_8 FILLER_0_31_102 ();
 sg13g2_fill_8 FILLER_0_31_110 ();
 sg13g2_fill_4 FILLER_0_31_118 ();
 sg13g2_fill_4 FILLER_0_31_157 ();
 sg13g2_fill_1 FILLER_0_31_161 ();
 sg13g2_fill_1 FILLER_0_31_166 ();
 sg13g2_fill_8 FILLER_0_31_203 ();
 sg13g2_fill_1 FILLER_0_31_211 ();
 sg13g2_fill_8 FILLER_0_31_248 ();
 sg13g2_fill_8 FILLER_0_31_256 ();
 sg13g2_decap_8 FILLER_0_31_264 ();
 sg13g2_fill_8 FILLER_0_31_302 ();
 sg13g2_fill_4 FILLER_0_31_310 ();
 sg13g2_fill_1 FILLER_0_31_314 ();
 sg13g2_fill_2 FILLER_0_31_319 ();
 sg13g2_fill_2 FILLER_0_31_339 ();
 sg13g2_fill_2 FILLER_0_31_349 ();
 sg13g2_fill_1 FILLER_0_31_351 ();
 sg13g2_fill_2 FILLER_0_31_356 ();
 sg13g2_fill_1 FILLER_0_31_358 ();
 sg13g2_fill_8 FILLER_0_31_390 ();
 sg13g2_fill_8 FILLER_0_31_398 ();
 sg13g2_fill_8 FILLER_0_31_406 ();
 sg13g2_fill_8 FILLER_0_31_414 ();
 sg13g2_fill_1 FILLER_0_31_539 ();
 sg13g2_fill_8 FILLER_0_31_571 ();
 sg13g2_fill_8 FILLER_0_31_579 ();
 sg13g2_fill_8 FILLER_0_31_587 ();
 sg13g2_fill_8 FILLER_0_31_595 ();
 sg13g2_fill_8 FILLER_0_31_603 ();
 sg13g2_fill_8 FILLER_0_31_611 ();
 sg13g2_fill_8 FILLER_0_31_619 ();
 sg13g2_fill_8 FILLER_0_31_627 ();
 sg13g2_fill_8 FILLER_0_31_635 ();
 sg13g2_fill_8 FILLER_0_31_643 ();
 sg13g2_fill_8 FILLER_0_31_651 ();
 sg13g2_fill_8 FILLER_0_31_659 ();
 sg13g2_fill_8 FILLER_0_31_667 ();
 sg13g2_fill_8 FILLER_0_31_675 ();
 sg13g2_fill_8 FILLER_0_31_683 ();
 sg13g2_fill_8 FILLER_0_31_691 ();
 sg13g2_fill_8 FILLER_0_31_699 ();
 sg13g2_fill_8 FILLER_0_31_707 ();
 sg13g2_fill_8 FILLER_0_31_715 ();
 sg13g2_fill_8 FILLER_0_31_723 ();
 sg13g2_fill_8 FILLER_0_31_731 ();
 sg13g2_fill_8 FILLER_0_31_739 ();
 sg13g2_fill_8 FILLER_0_31_747 ();
 sg13g2_fill_8 FILLER_0_31_755 ();
 sg13g2_fill_8 FILLER_0_31_763 ();
 sg13g2_fill_8 FILLER_0_31_771 ();
 sg13g2_fill_8 FILLER_0_31_779 ();
 sg13g2_fill_8 FILLER_0_31_787 ();
 sg13g2_fill_8 FILLER_0_31_795 ();
 sg13g2_fill_8 FILLER_0_31_803 ();
 sg13g2_fill_8 FILLER_0_31_811 ();
 sg13g2_fill_8 FILLER_0_31_819 ();
 sg13g2_fill_8 FILLER_0_31_827 ();
 sg13g2_fill_8 FILLER_0_31_835 ();
 sg13g2_fill_8 FILLER_0_31_843 ();
 sg13g2_fill_8 FILLER_0_31_851 ();
 sg13g2_fill_8 FILLER_0_31_859 ();
 sg13g2_fill_8 FILLER_0_31_867 ();
 sg13g2_fill_8 FILLER_0_31_875 ();
 sg13g2_fill_8 FILLER_0_31_883 ();
 sg13g2_fill_8 FILLER_0_31_891 ();
 sg13g2_fill_8 FILLER_0_31_899 ();
 sg13g2_fill_8 FILLER_0_31_907 ();
 sg13g2_fill_8 FILLER_0_31_915 ();
 sg13g2_fill_8 FILLER_0_31_923 ();
 sg13g2_fill_8 FILLER_0_31_931 ();
 sg13g2_fill_8 FILLER_0_31_939 ();
 sg13g2_fill_8 FILLER_0_31_947 ();
 sg13g2_fill_8 FILLER_0_31_955 ();
 sg13g2_fill_8 FILLER_0_31_963 ();
 sg13g2_fill_8 FILLER_0_31_971 ();
 sg13g2_fill_8 FILLER_0_31_979 ();
 sg13g2_fill_8 FILLER_0_31_987 ();
 sg13g2_fill_8 FILLER_0_31_995 ();
 sg13g2_fill_8 FILLER_0_31_1003 ();
 sg13g2_fill_8 FILLER_0_31_1011 ();
 sg13g2_fill_8 FILLER_0_31_1019 ();
 sg13g2_fill_8 FILLER_0_31_1027 ();
 sg13g2_fill_8 FILLER_0_31_1035 ();
 sg13g2_fill_8 FILLER_0_31_1043 ();
 sg13g2_fill_8 FILLER_0_31_1051 ();
 sg13g2_fill_8 FILLER_0_31_1059 ();
 sg13g2_fill_8 FILLER_0_31_1067 ();
 sg13g2_fill_8 FILLER_0_31_1075 ();
 sg13g2_fill_8 FILLER_0_31_1083 ();
 sg13g2_fill_8 FILLER_0_31_1091 ();
 sg13g2_fill_8 FILLER_0_31_1099 ();
 sg13g2_fill_8 FILLER_0_31_1107 ();
 sg13g2_fill_8 FILLER_0_31_1115 ();
 sg13g2_fill_8 FILLER_0_31_1123 ();
 sg13g2_fill_8 FILLER_0_31_1131 ();
 sg13g2_fill_8 FILLER_0_31_1139 ();
 sg13g2_fill_8 FILLER_0_31_1147 ();
 sg13g2_fill_8 FILLER_0_31_1155 ();
 sg13g2_fill_8 FILLER_0_31_1163 ();
 sg13g2_fill_8 FILLER_0_31_1171 ();
 sg13g2_fill_8 FILLER_0_31_1179 ();
 sg13g2_fill_8 FILLER_0_31_1187 ();
 sg13g2_fill_8 FILLER_0_31_1195 ();
 sg13g2_fill_8 FILLER_0_31_1203 ();
 sg13g2_fill_8 FILLER_0_31_1211 ();
 sg13g2_fill_8 FILLER_0_31_1219 ();
 sg13g2_fill_1 FILLER_0_31_1227 ();
 sg13g2_fill_4 FILLER_0_32_0 ();
 sg13g2_fill_1 FILLER_0_32_13 ();
 sg13g2_fill_1 FILLER_0_32_39 ();
 sg13g2_fill_1 FILLER_0_32_45 ();
 sg13g2_fill_4 FILLER_0_32_64 ();
 sg13g2_fill_2 FILLER_0_32_68 ();
 sg13g2_fill_1 FILLER_0_32_106 ();
 sg13g2_fill_2 FILLER_0_32_117 ();
 sg13g2_fill_1 FILLER_0_32_119 ();
 sg13g2_fill_1 FILLER_0_32_129 ();
 sg13g2_fill_2 FILLER_0_32_140 ();
 sg13g2_fill_8 FILLER_0_32_146 ();
 sg13g2_fill_4 FILLER_0_32_154 ();
 sg13g2_fill_2 FILLER_0_32_162 ();
 sg13g2_fill_1 FILLER_0_32_164 ();
 sg13g2_fill_2 FILLER_0_32_183 ();
 sg13g2_fill_2 FILLER_0_32_195 ();
 sg13g2_fill_1 FILLER_0_32_223 ();
 sg13g2_fill_1 FILLER_0_32_250 ();
 sg13g2_fill_1 FILLER_0_32_281 ();
 sg13g2_fill_2 FILLER_0_32_308 ();
 sg13g2_decap_8 FILLER_0_32_336 ();
 sg13g2_fill_2 FILLER_0_32_357 ();
 sg13g2_fill_4 FILLER_0_32_369 ();
 sg13g2_fill_8 FILLER_0_32_399 ();
 sg13g2_fill_8 FILLER_0_32_407 ();
 sg13g2_fill_2 FILLER_0_32_415 ();
 sg13g2_fill_1 FILLER_0_32_479 ();
 sg13g2_fill_2 FILLER_0_32_484 ();
 sg13g2_fill_8 FILLER_0_32_496 ();
 sg13g2_fill_2 FILLER_0_32_504 ();
 sg13g2_fill_4 FILLER_0_32_532 ();
 sg13g2_fill_4 FILLER_0_32_569 ();
 sg13g2_fill_8 FILLER_0_32_583 ();
 sg13g2_fill_8 FILLER_0_32_591 ();
 sg13g2_fill_8 FILLER_0_32_599 ();
 sg13g2_fill_8 FILLER_0_32_607 ();
 sg13g2_fill_8 FILLER_0_32_615 ();
 sg13g2_fill_8 FILLER_0_32_623 ();
 sg13g2_fill_8 FILLER_0_32_631 ();
 sg13g2_fill_8 FILLER_0_32_639 ();
 sg13g2_fill_8 FILLER_0_32_647 ();
 sg13g2_fill_8 FILLER_0_32_655 ();
 sg13g2_fill_8 FILLER_0_32_663 ();
 sg13g2_fill_8 FILLER_0_32_671 ();
 sg13g2_fill_8 FILLER_0_32_679 ();
 sg13g2_fill_8 FILLER_0_32_687 ();
 sg13g2_fill_8 FILLER_0_32_695 ();
 sg13g2_fill_8 FILLER_0_32_703 ();
 sg13g2_fill_8 FILLER_0_32_711 ();
 sg13g2_fill_8 FILLER_0_32_719 ();
 sg13g2_fill_8 FILLER_0_32_727 ();
 sg13g2_fill_8 FILLER_0_32_735 ();
 sg13g2_fill_8 FILLER_0_32_743 ();
 sg13g2_fill_8 FILLER_0_32_751 ();
 sg13g2_fill_8 FILLER_0_32_759 ();
 sg13g2_fill_8 FILLER_0_32_767 ();
 sg13g2_fill_8 FILLER_0_32_775 ();
 sg13g2_fill_8 FILLER_0_32_783 ();
 sg13g2_fill_8 FILLER_0_32_791 ();
 sg13g2_fill_8 FILLER_0_32_799 ();
 sg13g2_fill_8 FILLER_0_32_807 ();
 sg13g2_fill_8 FILLER_0_32_815 ();
 sg13g2_fill_8 FILLER_0_32_823 ();
 sg13g2_fill_8 FILLER_0_32_831 ();
 sg13g2_fill_8 FILLER_0_32_839 ();
 sg13g2_fill_8 FILLER_0_32_847 ();
 sg13g2_fill_8 FILLER_0_32_855 ();
 sg13g2_fill_8 FILLER_0_32_863 ();
 sg13g2_fill_8 FILLER_0_32_871 ();
 sg13g2_fill_8 FILLER_0_32_879 ();
 sg13g2_fill_8 FILLER_0_32_887 ();
 sg13g2_fill_8 FILLER_0_32_895 ();
 sg13g2_fill_8 FILLER_0_32_903 ();
 sg13g2_fill_8 FILLER_0_32_911 ();
 sg13g2_fill_8 FILLER_0_32_919 ();
 sg13g2_fill_8 FILLER_0_32_927 ();
 sg13g2_fill_8 FILLER_0_32_935 ();
 sg13g2_fill_8 FILLER_0_32_943 ();
 sg13g2_fill_8 FILLER_0_32_951 ();
 sg13g2_fill_8 FILLER_0_32_959 ();
 sg13g2_fill_8 FILLER_0_32_967 ();
 sg13g2_fill_8 FILLER_0_32_975 ();
 sg13g2_fill_8 FILLER_0_32_983 ();
 sg13g2_fill_8 FILLER_0_32_991 ();
 sg13g2_fill_8 FILLER_0_32_999 ();
 sg13g2_fill_8 FILLER_0_32_1007 ();
 sg13g2_fill_8 FILLER_0_32_1015 ();
 sg13g2_fill_8 FILLER_0_32_1023 ();
 sg13g2_fill_8 FILLER_0_32_1031 ();
 sg13g2_fill_8 FILLER_0_32_1039 ();
 sg13g2_fill_8 FILLER_0_32_1047 ();
 sg13g2_fill_8 FILLER_0_32_1055 ();
 sg13g2_fill_8 FILLER_0_32_1063 ();
 sg13g2_fill_8 FILLER_0_32_1071 ();
 sg13g2_fill_8 FILLER_0_32_1079 ();
 sg13g2_fill_8 FILLER_0_32_1087 ();
 sg13g2_fill_8 FILLER_0_32_1095 ();
 sg13g2_fill_8 FILLER_0_32_1103 ();
 sg13g2_fill_8 FILLER_0_32_1111 ();
 sg13g2_fill_8 FILLER_0_32_1119 ();
 sg13g2_fill_8 FILLER_0_32_1127 ();
 sg13g2_fill_8 FILLER_0_32_1135 ();
 sg13g2_fill_8 FILLER_0_32_1143 ();
 sg13g2_fill_8 FILLER_0_32_1151 ();
 sg13g2_fill_8 FILLER_0_32_1159 ();
 sg13g2_fill_8 FILLER_0_32_1167 ();
 sg13g2_fill_8 FILLER_0_32_1175 ();
 sg13g2_fill_8 FILLER_0_32_1183 ();
 sg13g2_fill_8 FILLER_0_32_1191 ();
 sg13g2_fill_8 FILLER_0_32_1199 ();
 sg13g2_fill_8 FILLER_0_32_1207 ();
 sg13g2_fill_8 FILLER_0_32_1215 ();
 sg13g2_fill_4 FILLER_0_32_1223 ();
 sg13g2_fill_1 FILLER_0_32_1227 ();
 sg13g2_fill_8 FILLER_0_33_0 ();
 sg13g2_fill_8 FILLER_0_33_8 ();
 sg13g2_fill_2 FILLER_0_33_16 ();
 sg13g2_fill_1 FILLER_0_33_18 ();
 sg13g2_fill_8 FILLER_0_33_152 ();
 sg13g2_fill_4 FILLER_0_33_160 ();
 sg13g2_fill_1 FILLER_0_33_164 ();
 sg13g2_fill_4 FILLER_0_33_174 ();
 sg13g2_fill_4 FILLER_0_33_182 ();
 sg13g2_fill_1 FILLER_0_33_186 ();
 sg13g2_fill_8 FILLER_0_33_211 ();
 sg13g2_fill_4 FILLER_0_33_219 ();
 sg13g2_fill_2 FILLER_0_33_223 ();
 sg13g2_fill_2 FILLER_0_33_234 ();
 sg13g2_fill_4 FILLER_0_33_262 ();
 sg13g2_fill_4 FILLER_0_33_274 ();
 sg13g2_fill_4 FILLER_0_33_304 ();
 sg13g2_fill_8 FILLER_0_33_312 ();
 sg13g2_fill_4 FILLER_0_33_320 ();
 sg13g2_fill_1 FILLER_0_33_324 ();
 sg13g2_fill_2 FILLER_0_33_356 ();
 sg13g2_fill_2 FILLER_0_33_445 ();
 sg13g2_fill_1 FILLER_0_33_447 ();
 sg13g2_fill_8 FILLER_0_33_460 ();
 sg13g2_fill_1 FILLER_0_33_468 ();
 sg13g2_fill_2 FILLER_0_33_474 ();
 sg13g2_fill_8 FILLER_0_33_486 ();
 sg13g2_fill_8 FILLER_0_33_494 ();
 sg13g2_fill_2 FILLER_0_33_502 ();
 sg13g2_fill_1 FILLER_0_33_504 ();
 sg13g2_fill_2 FILLER_0_33_514 ();
 sg13g2_fill_8 FILLER_0_33_526 ();
 sg13g2_decap_8 FILLER_0_33_534 ();
 sg13g2_fill_2 FILLER_0_33_571 ();
 sg13g2_fill_8 FILLER_0_33_604 ();
 sg13g2_fill_8 FILLER_0_33_612 ();
 sg13g2_fill_8 FILLER_0_33_620 ();
 sg13g2_fill_8 FILLER_0_33_628 ();
 sg13g2_fill_8 FILLER_0_33_636 ();
 sg13g2_fill_8 FILLER_0_33_644 ();
 sg13g2_fill_8 FILLER_0_33_652 ();
 sg13g2_fill_8 FILLER_0_33_660 ();
 sg13g2_fill_8 FILLER_0_33_668 ();
 sg13g2_fill_8 FILLER_0_33_676 ();
 sg13g2_fill_8 FILLER_0_33_684 ();
 sg13g2_fill_8 FILLER_0_33_692 ();
 sg13g2_fill_8 FILLER_0_33_700 ();
 sg13g2_fill_8 FILLER_0_33_708 ();
 sg13g2_fill_8 FILLER_0_33_716 ();
 sg13g2_fill_8 FILLER_0_33_724 ();
 sg13g2_fill_8 FILLER_0_33_732 ();
 sg13g2_fill_8 FILLER_0_33_740 ();
 sg13g2_fill_8 FILLER_0_33_748 ();
 sg13g2_fill_8 FILLER_0_33_756 ();
 sg13g2_fill_8 FILLER_0_33_764 ();
 sg13g2_fill_8 FILLER_0_33_772 ();
 sg13g2_fill_8 FILLER_0_33_780 ();
 sg13g2_fill_8 FILLER_0_33_788 ();
 sg13g2_fill_8 FILLER_0_33_796 ();
 sg13g2_fill_8 FILLER_0_33_804 ();
 sg13g2_fill_8 FILLER_0_33_812 ();
 sg13g2_fill_8 FILLER_0_33_820 ();
 sg13g2_fill_8 FILLER_0_33_828 ();
 sg13g2_fill_8 FILLER_0_33_836 ();
 sg13g2_fill_8 FILLER_0_33_844 ();
 sg13g2_fill_8 FILLER_0_33_852 ();
 sg13g2_fill_8 FILLER_0_33_860 ();
 sg13g2_fill_8 FILLER_0_33_868 ();
 sg13g2_fill_8 FILLER_0_33_876 ();
 sg13g2_fill_8 FILLER_0_33_884 ();
 sg13g2_fill_8 FILLER_0_33_892 ();
 sg13g2_fill_8 FILLER_0_33_900 ();
 sg13g2_fill_8 FILLER_0_33_908 ();
 sg13g2_fill_8 FILLER_0_33_916 ();
 sg13g2_fill_8 FILLER_0_33_924 ();
 sg13g2_fill_8 FILLER_0_33_932 ();
 sg13g2_fill_8 FILLER_0_33_940 ();
 sg13g2_fill_8 FILLER_0_33_948 ();
 sg13g2_fill_8 FILLER_0_33_956 ();
 sg13g2_fill_8 FILLER_0_33_964 ();
 sg13g2_fill_8 FILLER_0_33_972 ();
 sg13g2_fill_8 FILLER_0_33_980 ();
 sg13g2_fill_8 FILLER_0_33_988 ();
 sg13g2_fill_8 FILLER_0_33_996 ();
 sg13g2_fill_8 FILLER_0_33_1004 ();
 sg13g2_fill_8 FILLER_0_33_1012 ();
 sg13g2_fill_8 FILLER_0_33_1020 ();
 sg13g2_fill_8 FILLER_0_33_1028 ();
 sg13g2_fill_8 FILLER_0_33_1036 ();
 sg13g2_fill_8 FILLER_0_33_1044 ();
 sg13g2_fill_8 FILLER_0_33_1052 ();
 sg13g2_fill_8 FILLER_0_33_1060 ();
 sg13g2_fill_8 FILLER_0_33_1068 ();
 sg13g2_fill_8 FILLER_0_33_1076 ();
 sg13g2_fill_8 FILLER_0_33_1084 ();
 sg13g2_fill_8 FILLER_0_33_1092 ();
 sg13g2_fill_8 FILLER_0_33_1100 ();
 sg13g2_fill_8 FILLER_0_33_1108 ();
 sg13g2_fill_8 FILLER_0_33_1116 ();
 sg13g2_fill_8 FILLER_0_33_1124 ();
 sg13g2_fill_8 FILLER_0_33_1132 ();
 sg13g2_fill_8 FILLER_0_33_1140 ();
 sg13g2_fill_8 FILLER_0_33_1148 ();
 sg13g2_fill_8 FILLER_0_33_1156 ();
 sg13g2_fill_8 FILLER_0_33_1164 ();
 sg13g2_fill_8 FILLER_0_33_1172 ();
 sg13g2_fill_8 FILLER_0_33_1180 ();
 sg13g2_fill_8 FILLER_0_33_1188 ();
 sg13g2_fill_8 FILLER_0_33_1196 ();
 sg13g2_fill_8 FILLER_0_33_1204 ();
 sg13g2_fill_8 FILLER_0_33_1212 ();
 sg13g2_fill_8 FILLER_0_33_1220 ();
 sg13g2_fill_8 FILLER_0_34_0 ();
 sg13g2_fill_4 FILLER_0_34_8 ();
 sg13g2_fill_1 FILLER_0_34_12 ();
 sg13g2_fill_1 FILLER_0_34_48 ();
 sg13g2_fill_8 FILLER_0_34_53 ();
 sg13g2_fill_8 FILLER_0_34_61 ();
 sg13g2_fill_8 FILLER_0_34_69 ();
 sg13g2_fill_8 FILLER_0_34_81 ();
 sg13g2_fill_1 FILLER_0_34_89 ();
 sg13g2_fill_1 FILLER_0_34_95 ();
 sg13g2_fill_2 FILLER_0_34_122 ();
 sg13g2_fill_1 FILLER_0_34_124 ();
 sg13g2_fill_2 FILLER_0_34_155 ();
 sg13g2_fill_1 FILLER_0_34_157 ();
 sg13g2_fill_2 FILLER_0_34_162 ();
 sg13g2_fill_1 FILLER_0_34_164 ();
 sg13g2_fill_2 FILLER_0_34_191 ();
 sg13g2_fill_1 FILLER_0_34_203 ();
 sg13g2_fill_8 FILLER_0_34_209 ();
 sg13g2_fill_8 FILLER_0_34_217 ();
 sg13g2_fill_8 FILLER_0_34_225 ();
 sg13g2_fill_1 FILLER_0_34_233 ();
 sg13g2_fill_1 FILLER_0_34_268 ();
 sg13g2_fill_2 FILLER_0_34_284 ();
 sg13g2_fill_8 FILLER_0_34_290 ();
 sg13g2_fill_2 FILLER_0_34_298 ();
 sg13g2_fill_1 FILLER_0_34_300 ();
 sg13g2_fill_4 FILLER_0_34_332 ();
 sg13g2_fill_1 FILLER_0_34_336 ();
 sg13g2_fill_8 FILLER_0_34_341 ();
 sg13g2_fill_1 FILLER_0_34_359 ();
 sg13g2_fill_2 FILLER_0_34_364 ();
 sg13g2_fill_1 FILLER_0_34_366 ();
 sg13g2_fill_4 FILLER_0_34_377 ();
 sg13g2_fill_2 FILLER_0_34_381 ();
 sg13g2_fill_2 FILLER_0_34_387 ();
 sg13g2_fill_1 FILLER_0_34_393 ();
 sg13g2_fill_1 FILLER_0_34_420 ();
 sg13g2_fill_8 FILLER_0_34_448 ();
 sg13g2_fill_4 FILLER_0_34_456 ();
 sg13g2_fill_1 FILLER_0_34_460 ();
 sg13g2_fill_8 FILLER_0_34_487 ();
 sg13g2_fill_8 FILLER_0_34_495 ();
 sg13g2_fill_8 FILLER_0_34_503 ();
 sg13g2_fill_2 FILLER_0_34_511 ();
 sg13g2_fill_1 FILLER_0_34_513 ();
 sg13g2_fill_2 FILLER_0_34_575 ();
 sg13g2_fill_1 FILLER_0_34_577 ();
 sg13g2_fill_4 FILLER_0_34_608 ();
 sg13g2_fill_1 FILLER_0_34_612 ();
 sg13g2_fill_8 FILLER_0_34_621 ();
 sg13g2_fill_8 FILLER_0_34_629 ();
 sg13g2_fill_8 FILLER_0_34_637 ();
 sg13g2_fill_8 FILLER_0_34_645 ();
 sg13g2_fill_8 FILLER_0_34_653 ();
 sg13g2_fill_8 FILLER_0_34_661 ();
 sg13g2_fill_8 FILLER_0_34_669 ();
 sg13g2_fill_8 FILLER_0_34_677 ();
 sg13g2_fill_8 FILLER_0_34_685 ();
 sg13g2_fill_8 FILLER_0_34_693 ();
 sg13g2_fill_8 FILLER_0_34_701 ();
 sg13g2_fill_8 FILLER_0_34_709 ();
 sg13g2_fill_8 FILLER_0_34_717 ();
 sg13g2_fill_8 FILLER_0_34_725 ();
 sg13g2_fill_8 FILLER_0_34_733 ();
 sg13g2_fill_8 FILLER_0_34_741 ();
 sg13g2_fill_8 FILLER_0_34_749 ();
 sg13g2_fill_8 FILLER_0_34_757 ();
 sg13g2_fill_8 FILLER_0_34_765 ();
 sg13g2_fill_8 FILLER_0_34_773 ();
 sg13g2_fill_8 FILLER_0_34_781 ();
 sg13g2_fill_8 FILLER_0_34_789 ();
 sg13g2_fill_8 FILLER_0_34_797 ();
 sg13g2_fill_8 FILLER_0_34_805 ();
 sg13g2_fill_8 FILLER_0_34_813 ();
 sg13g2_fill_8 FILLER_0_34_821 ();
 sg13g2_fill_8 FILLER_0_34_829 ();
 sg13g2_fill_8 FILLER_0_34_837 ();
 sg13g2_fill_8 FILLER_0_34_845 ();
 sg13g2_fill_8 FILLER_0_34_853 ();
 sg13g2_fill_8 FILLER_0_34_861 ();
 sg13g2_fill_8 FILLER_0_34_869 ();
 sg13g2_fill_8 FILLER_0_34_877 ();
 sg13g2_fill_8 FILLER_0_34_885 ();
 sg13g2_fill_8 FILLER_0_34_893 ();
 sg13g2_fill_8 FILLER_0_34_901 ();
 sg13g2_fill_8 FILLER_0_34_909 ();
 sg13g2_fill_8 FILLER_0_34_917 ();
 sg13g2_fill_8 FILLER_0_34_925 ();
 sg13g2_fill_8 FILLER_0_34_933 ();
 sg13g2_fill_8 FILLER_0_34_941 ();
 sg13g2_fill_8 FILLER_0_34_949 ();
 sg13g2_fill_8 FILLER_0_34_957 ();
 sg13g2_fill_8 FILLER_0_34_965 ();
 sg13g2_fill_8 FILLER_0_34_973 ();
 sg13g2_fill_8 FILLER_0_34_981 ();
 sg13g2_fill_8 FILLER_0_34_989 ();
 sg13g2_fill_8 FILLER_0_34_997 ();
 sg13g2_fill_8 FILLER_0_34_1005 ();
 sg13g2_fill_8 FILLER_0_34_1013 ();
 sg13g2_fill_8 FILLER_0_34_1021 ();
 sg13g2_fill_8 FILLER_0_34_1029 ();
 sg13g2_fill_8 FILLER_0_34_1037 ();
 sg13g2_fill_8 FILLER_0_34_1045 ();
 sg13g2_fill_8 FILLER_0_34_1053 ();
 sg13g2_fill_8 FILLER_0_34_1061 ();
 sg13g2_fill_8 FILLER_0_34_1069 ();
 sg13g2_fill_8 FILLER_0_34_1077 ();
 sg13g2_fill_8 FILLER_0_34_1085 ();
 sg13g2_fill_8 FILLER_0_34_1093 ();
 sg13g2_fill_8 FILLER_0_34_1101 ();
 sg13g2_fill_8 FILLER_0_34_1109 ();
 sg13g2_fill_8 FILLER_0_34_1117 ();
 sg13g2_fill_8 FILLER_0_34_1125 ();
 sg13g2_fill_8 FILLER_0_34_1133 ();
 sg13g2_fill_8 FILLER_0_34_1141 ();
 sg13g2_fill_8 FILLER_0_34_1149 ();
 sg13g2_fill_8 FILLER_0_34_1157 ();
 sg13g2_fill_8 FILLER_0_34_1165 ();
 sg13g2_fill_8 FILLER_0_34_1173 ();
 sg13g2_fill_8 FILLER_0_34_1181 ();
 sg13g2_fill_8 FILLER_0_34_1189 ();
 sg13g2_fill_8 FILLER_0_34_1197 ();
 sg13g2_fill_8 FILLER_0_34_1205 ();
 sg13g2_fill_8 FILLER_0_34_1213 ();
 sg13g2_decap_8 FILLER_0_34_1221 ();
 sg13g2_fill_1 FILLER_0_35_0 ();
 sg13g2_fill_2 FILLER_0_35_27 ();
 sg13g2_fill_1 FILLER_0_35_60 ();
 sg13g2_fill_4 FILLER_0_35_88 ();
 sg13g2_fill_1 FILLER_0_35_92 ();
 sg13g2_fill_4 FILLER_0_35_97 ();
 sg13g2_fill_2 FILLER_0_35_101 ();
 sg13g2_fill_1 FILLER_0_35_107 ();
 sg13g2_fill_4 FILLER_0_35_120 ();
 sg13g2_fill_2 FILLER_0_35_124 ();
 sg13g2_fill_2 FILLER_0_35_131 ();
 sg13g2_decap_8 FILLER_0_35_147 ();
 sg13g2_fill_2 FILLER_0_35_180 ();
 sg13g2_fill_2 FILLER_0_35_192 ();
 sg13g2_fill_1 FILLER_0_35_194 ();
 sg13g2_fill_8 FILLER_0_35_226 ();
 sg13g2_fill_4 FILLER_0_35_234 ();
 sg13g2_fill_1 FILLER_0_35_238 ();
 sg13g2_fill_4 FILLER_0_35_243 ();
 sg13g2_fill_1 FILLER_0_35_247 ();
 sg13g2_decap_8 FILLER_0_35_256 ();
 sg13g2_fill_8 FILLER_0_35_267 ();
 sg13g2_fill_8 FILLER_0_35_275 ();
 sg13g2_fill_2 FILLER_0_35_283 ();
 sg13g2_fill_1 FILLER_0_35_285 ();
 sg13g2_fill_4 FILLER_0_35_301 ();
 sg13g2_fill_2 FILLER_0_35_305 ();
 sg13g2_fill_4 FILLER_0_35_315 ();
 sg13g2_fill_8 FILLER_0_35_329 ();
 sg13g2_fill_8 FILLER_0_35_337 ();
 sg13g2_fill_1 FILLER_0_35_345 ();
 sg13g2_fill_8 FILLER_0_35_377 ();
 sg13g2_fill_8 FILLER_0_35_385 ();
 sg13g2_fill_8 FILLER_0_35_393 ();
 sg13g2_fill_2 FILLER_0_35_401 ();
 sg13g2_fill_1 FILLER_0_35_412 ();
 sg13g2_fill_1 FILLER_0_35_417 ();
 sg13g2_fill_2 FILLER_0_35_433 ();
 sg13g2_fill_2 FILLER_0_35_461 ();
 sg13g2_fill_1 FILLER_0_35_463 ();
 sg13g2_fill_4 FILLER_0_35_490 ();
 sg13g2_fill_1 FILLER_0_35_494 ();
 sg13g2_fill_2 FILLER_0_35_531 ();
 sg13g2_fill_1 FILLER_0_35_533 ();
 sg13g2_fill_4 FILLER_0_35_547 ();
 sg13g2_fill_1 FILLER_0_35_551 ();
 sg13g2_fill_8 FILLER_0_35_556 ();
 sg13g2_fill_8 FILLER_0_35_564 ();
 sg13g2_fill_4 FILLER_0_35_572 ();
 sg13g2_fill_2 FILLER_0_35_576 ();
 sg13g2_fill_8 FILLER_0_35_597 ();
 sg13g2_fill_8 FILLER_0_35_605 ();
 sg13g2_fill_8 FILLER_0_35_613 ();
 sg13g2_fill_8 FILLER_0_35_621 ();
 sg13g2_fill_8 FILLER_0_35_629 ();
 sg13g2_fill_8 FILLER_0_35_637 ();
 sg13g2_fill_8 FILLER_0_35_645 ();
 sg13g2_fill_8 FILLER_0_35_653 ();
 sg13g2_fill_8 FILLER_0_35_661 ();
 sg13g2_fill_8 FILLER_0_35_669 ();
 sg13g2_fill_8 FILLER_0_35_677 ();
 sg13g2_fill_8 FILLER_0_35_685 ();
 sg13g2_fill_8 FILLER_0_35_693 ();
 sg13g2_fill_8 FILLER_0_35_701 ();
 sg13g2_fill_8 FILLER_0_35_709 ();
 sg13g2_fill_8 FILLER_0_35_717 ();
 sg13g2_fill_8 FILLER_0_35_725 ();
 sg13g2_fill_8 FILLER_0_35_733 ();
 sg13g2_fill_8 FILLER_0_35_741 ();
 sg13g2_fill_8 FILLER_0_35_749 ();
 sg13g2_fill_8 FILLER_0_35_757 ();
 sg13g2_fill_8 FILLER_0_35_765 ();
 sg13g2_fill_8 FILLER_0_35_773 ();
 sg13g2_fill_8 FILLER_0_35_781 ();
 sg13g2_fill_8 FILLER_0_35_789 ();
 sg13g2_fill_8 FILLER_0_35_797 ();
 sg13g2_fill_8 FILLER_0_35_805 ();
 sg13g2_fill_8 FILLER_0_35_813 ();
 sg13g2_fill_8 FILLER_0_35_821 ();
 sg13g2_fill_8 FILLER_0_35_829 ();
 sg13g2_fill_8 FILLER_0_35_837 ();
 sg13g2_fill_8 FILLER_0_35_845 ();
 sg13g2_fill_8 FILLER_0_35_853 ();
 sg13g2_fill_8 FILLER_0_35_861 ();
 sg13g2_fill_8 FILLER_0_35_869 ();
 sg13g2_fill_8 FILLER_0_35_877 ();
 sg13g2_fill_8 FILLER_0_35_885 ();
 sg13g2_fill_8 FILLER_0_35_893 ();
 sg13g2_fill_8 FILLER_0_35_901 ();
 sg13g2_fill_8 FILLER_0_35_909 ();
 sg13g2_fill_8 FILLER_0_35_917 ();
 sg13g2_fill_8 FILLER_0_35_925 ();
 sg13g2_fill_8 FILLER_0_35_933 ();
 sg13g2_fill_8 FILLER_0_35_941 ();
 sg13g2_fill_8 FILLER_0_35_949 ();
 sg13g2_fill_8 FILLER_0_35_957 ();
 sg13g2_fill_8 FILLER_0_35_965 ();
 sg13g2_fill_8 FILLER_0_35_973 ();
 sg13g2_fill_8 FILLER_0_35_981 ();
 sg13g2_fill_8 FILLER_0_35_989 ();
 sg13g2_fill_8 FILLER_0_35_997 ();
 sg13g2_fill_8 FILLER_0_35_1005 ();
 sg13g2_fill_8 FILLER_0_35_1013 ();
 sg13g2_fill_8 FILLER_0_35_1021 ();
 sg13g2_fill_8 FILLER_0_35_1029 ();
 sg13g2_fill_8 FILLER_0_35_1037 ();
 sg13g2_fill_8 FILLER_0_35_1045 ();
 sg13g2_fill_8 FILLER_0_35_1053 ();
 sg13g2_fill_8 FILLER_0_35_1061 ();
 sg13g2_fill_8 FILLER_0_35_1069 ();
 sg13g2_fill_8 FILLER_0_35_1077 ();
 sg13g2_fill_8 FILLER_0_35_1085 ();
 sg13g2_fill_8 FILLER_0_35_1093 ();
 sg13g2_fill_8 FILLER_0_35_1101 ();
 sg13g2_fill_8 FILLER_0_35_1109 ();
 sg13g2_fill_8 FILLER_0_35_1117 ();
 sg13g2_fill_8 FILLER_0_35_1125 ();
 sg13g2_fill_8 FILLER_0_35_1133 ();
 sg13g2_fill_8 FILLER_0_35_1141 ();
 sg13g2_fill_8 FILLER_0_35_1149 ();
 sg13g2_fill_8 FILLER_0_35_1157 ();
 sg13g2_fill_8 FILLER_0_35_1165 ();
 sg13g2_fill_8 FILLER_0_35_1173 ();
 sg13g2_fill_8 FILLER_0_35_1181 ();
 sg13g2_fill_8 FILLER_0_35_1189 ();
 sg13g2_fill_8 FILLER_0_35_1197 ();
 sg13g2_fill_8 FILLER_0_35_1205 ();
 sg13g2_fill_8 FILLER_0_35_1213 ();
 sg13g2_decap_8 FILLER_0_35_1221 ();
 sg13g2_fill_4 FILLER_0_36_0 ();
 sg13g2_fill_1 FILLER_0_36_4 ();
 sg13g2_fill_1 FILLER_0_36_22 ();
 sg13g2_fill_1 FILLER_0_36_33 ();
 sg13g2_fill_2 FILLER_0_36_44 ();
 sg13g2_decap_8 FILLER_0_36_56 ();
 sg13g2_fill_8 FILLER_0_36_89 ();
 sg13g2_fill_8 FILLER_0_36_97 ();
 sg13g2_fill_4 FILLER_0_36_105 ();
 sg13g2_fill_1 FILLER_0_36_109 ();
 sg13g2_fill_4 FILLER_0_36_120 ();
 sg13g2_fill_2 FILLER_0_36_149 ();
 sg13g2_fill_1 FILLER_0_36_151 ();
 sg13g2_fill_1 FILLER_0_36_204 ();
 sg13g2_fill_1 FILLER_0_36_231 ();
 sg13g2_fill_4 FILLER_0_36_263 ();
 sg13g2_fill_1 FILLER_0_36_267 ();
 sg13g2_fill_1 FILLER_0_36_277 ();
 sg13g2_fill_2 FILLER_0_36_282 ();
 sg13g2_fill_4 FILLER_0_36_294 ();
 sg13g2_fill_4 FILLER_0_36_324 ();
 sg13g2_fill_2 FILLER_0_36_328 ();
 sg13g2_fill_4 FILLER_0_36_403 ();
 sg13g2_fill_1 FILLER_0_36_412 ();
 sg13g2_fill_1 FILLER_0_36_423 ();
 sg13g2_fill_1 FILLER_0_36_434 ();
 sg13g2_fill_2 FILLER_0_36_461 ();
 sg13g2_fill_2 FILLER_0_36_467 ();
 sg13g2_fill_2 FILLER_0_36_479 ();
 sg13g2_fill_2 FILLER_0_36_507 ();
 sg13g2_fill_1 FILLER_0_36_509 ();
 sg13g2_fill_2 FILLER_0_36_546 ();
 sg13g2_fill_1 FILLER_0_36_548 ();
 sg13g2_fill_8 FILLER_0_36_593 ();
 sg13g2_fill_8 FILLER_0_36_601 ();
 sg13g2_fill_8 FILLER_0_36_609 ();
 sg13g2_fill_8 FILLER_0_36_617 ();
 sg13g2_fill_8 FILLER_0_36_625 ();
 sg13g2_fill_8 FILLER_0_36_633 ();
 sg13g2_fill_8 FILLER_0_36_641 ();
 sg13g2_fill_8 FILLER_0_36_649 ();
 sg13g2_fill_8 FILLER_0_36_657 ();
 sg13g2_fill_8 FILLER_0_36_665 ();
 sg13g2_fill_8 FILLER_0_36_673 ();
 sg13g2_fill_8 FILLER_0_36_681 ();
 sg13g2_fill_8 FILLER_0_36_689 ();
 sg13g2_fill_8 FILLER_0_36_697 ();
 sg13g2_fill_8 FILLER_0_36_705 ();
 sg13g2_fill_8 FILLER_0_36_713 ();
 sg13g2_fill_8 FILLER_0_36_721 ();
 sg13g2_fill_8 FILLER_0_36_729 ();
 sg13g2_fill_8 FILLER_0_36_737 ();
 sg13g2_fill_8 FILLER_0_36_745 ();
 sg13g2_fill_8 FILLER_0_36_753 ();
 sg13g2_fill_8 FILLER_0_36_761 ();
 sg13g2_fill_8 FILLER_0_36_769 ();
 sg13g2_fill_8 FILLER_0_36_777 ();
 sg13g2_fill_8 FILLER_0_36_785 ();
 sg13g2_fill_8 FILLER_0_36_793 ();
 sg13g2_fill_8 FILLER_0_36_801 ();
 sg13g2_fill_8 FILLER_0_36_809 ();
 sg13g2_fill_8 FILLER_0_36_817 ();
 sg13g2_fill_8 FILLER_0_36_825 ();
 sg13g2_fill_8 FILLER_0_36_833 ();
 sg13g2_fill_8 FILLER_0_36_841 ();
 sg13g2_fill_8 FILLER_0_36_849 ();
 sg13g2_fill_8 FILLER_0_36_857 ();
 sg13g2_fill_8 FILLER_0_36_865 ();
 sg13g2_fill_8 FILLER_0_36_873 ();
 sg13g2_fill_8 FILLER_0_36_881 ();
 sg13g2_fill_8 FILLER_0_36_889 ();
 sg13g2_fill_8 FILLER_0_36_897 ();
 sg13g2_fill_8 FILLER_0_36_905 ();
 sg13g2_fill_8 FILLER_0_36_913 ();
 sg13g2_fill_8 FILLER_0_36_921 ();
 sg13g2_fill_8 FILLER_0_36_929 ();
 sg13g2_fill_8 FILLER_0_36_937 ();
 sg13g2_fill_8 FILLER_0_36_945 ();
 sg13g2_fill_8 FILLER_0_36_953 ();
 sg13g2_fill_8 FILLER_0_36_961 ();
 sg13g2_fill_8 FILLER_0_36_969 ();
 sg13g2_fill_8 FILLER_0_36_977 ();
 sg13g2_fill_8 FILLER_0_36_985 ();
 sg13g2_fill_8 FILLER_0_36_993 ();
 sg13g2_fill_8 FILLER_0_36_1001 ();
 sg13g2_fill_8 FILLER_0_36_1009 ();
 sg13g2_fill_8 FILLER_0_36_1017 ();
 sg13g2_fill_8 FILLER_0_36_1025 ();
 sg13g2_fill_8 FILLER_0_36_1033 ();
 sg13g2_fill_8 FILLER_0_36_1041 ();
 sg13g2_fill_8 FILLER_0_36_1049 ();
 sg13g2_fill_8 FILLER_0_36_1057 ();
 sg13g2_fill_8 FILLER_0_36_1065 ();
 sg13g2_fill_8 FILLER_0_36_1073 ();
 sg13g2_fill_8 FILLER_0_36_1081 ();
 sg13g2_fill_8 FILLER_0_36_1089 ();
 sg13g2_fill_8 FILLER_0_36_1097 ();
 sg13g2_fill_8 FILLER_0_36_1105 ();
 sg13g2_fill_8 FILLER_0_36_1113 ();
 sg13g2_fill_8 FILLER_0_36_1121 ();
 sg13g2_fill_8 FILLER_0_36_1129 ();
 sg13g2_fill_8 FILLER_0_36_1137 ();
 sg13g2_fill_8 FILLER_0_36_1145 ();
 sg13g2_fill_8 FILLER_0_36_1153 ();
 sg13g2_fill_8 FILLER_0_36_1161 ();
 sg13g2_fill_8 FILLER_0_36_1169 ();
 sg13g2_fill_8 FILLER_0_36_1177 ();
 sg13g2_fill_8 FILLER_0_36_1185 ();
 sg13g2_fill_8 FILLER_0_36_1193 ();
 sg13g2_fill_8 FILLER_0_36_1201 ();
 sg13g2_fill_8 FILLER_0_36_1209 ();
 sg13g2_fill_8 FILLER_0_36_1217 ();
 sg13g2_fill_2 FILLER_0_36_1225 ();
 sg13g2_fill_1 FILLER_0_36_1227 ();
 sg13g2_decap_8 FILLER_0_37_0 ();
 sg13g2_fill_2 FILLER_0_37_11 ();
 sg13g2_fill_1 FILLER_0_37_13 ();
 sg13g2_fill_2 FILLER_0_37_33 ();
 sg13g2_fill_4 FILLER_0_37_39 ();
 sg13g2_fill_1 FILLER_0_37_43 ();
 sg13g2_fill_8 FILLER_0_37_78 ();
 sg13g2_fill_2 FILLER_0_37_86 ();
 sg13g2_fill_1 FILLER_0_37_88 ();
 sg13g2_fill_2 FILLER_0_37_115 ();
 sg13g2_fill_4 FILLER_0_37_152 ();
 sg13g2_fill_2 FILLER_0_37_165 ();
 sg13g2_fill_1 FILLER_0_37_167 ();
 sg13g2_fill_2 FILLER_0_37_173 ();
 sg13g2_fill_1 FILLER_0_37_193 ();
 sg13g2_fill_8 FILLER_0_37_224 ();
 sg13g2_fill_2 FILLER_0_37_232 ();
 sg13g2_fill_1 FILLER_0_37_234 ();
 sg13g2_fill_8 FILLER_0_37_349 ();
 sg13g2_fill_1 FILLER_0_37_357 ();
 sg13g2_fill_8 FILLER_0_37_378 ();
 sg13g2_fill_8 FILLER_0_37_386 ();
 sg13g2_fill_2 FILLER_0_37_394 ();
 sg13g2_fill_2 FILLER_0_37_451 ();
 sg13g2_fill_1 FILLER_0_37_461 ();
 sg13g2_fill_1 FILLER_0_37_466 ();
 sg13g2_fill_1 FILLER_0_37_495 ();
 sg13g2_fill_2 FILLER_0_37_500 ();
 sg13g2_fill_1 FILLER_0_37_526 ();
 sg13g2_fill_1 FILLER_0_37_531 ();
 sg13g2_fill_2 FILLER_0_37_536 ();
 sg13g2_fill_2 FILLER_0_37_542 ();
 sg13g2_fill_1 FILLER_0_37_549 ();
 sg13g2_fill_2 FILLER_0_37_554 ();
 sg13g2_fill_2 FILLER_0_37_561 ();
 sg13g2_fill_2 FILLER_0_37_589 ();
 sg13g2_fill_8 FILLER_0_37_631 ();
 sg13g2_fill_8 FILLER_0_37_639 ();
 sg13g2_fill_8 FILLER_0_37_647 ();
 sg13g2_fill_8 FILLER_0_37_655 ();
 sg13g2_fill_8 FILLER_0_37_663 ();
 sg13g2_fill_8 FILLER_0_37_671 ();
 sg13g2_fill_8 FILLER_0_37_679 ();
 sg13g2_fill_8 FILLER_0_37_687 ();
 sg13g2_fill_8 FILLER_0_37_695 ();
 sg13g2_fill_8 FILLER_0_37_703 ();
 sg13g2_fill_8 FILLER_0_37_711 ();
 sg13g2_fill_8 FILLER_0_37_719 ();
 sg13g2_fill_8 FILLER_0_37_727 ();
 sg13g2_fill_8 FILLER_0_37_735 ();
 sg13g2_fill_8 FILLER_0_37_743 ();
 sg13g2_fill_8 FILLER_0_37_751 ();
 sg13g2_fill_8 FILLER_0_37_759 ();
 sg13g2_fill_8 FILLER_0_37_767 ();
 sg13g2_fill_8 FILLER_0_37_775 ();
 sg13g2_fill_8 FILLER_0_37_783 ();
 sg13g2_fill_8 FILLER_0_37_791 ();
 sg13g2_fill_8 FILLER_0_37_799 ();
 sg13g2_fill_8 FILLER_0_37_807 ();
 sg13g2_fill_8 FILLER_0_37_815 ();
 sg13g2_fill_8 FILLER_0_37_823 ();
 sg13g2_fill_8 FILLER_0_37_831 ();
 sg13g2_fill_8 FILLER_0_37_839 ();
 sg13g2_fill_8 FILLER_0_37_847 ();
 sg13g2_fill_8 FILLER_0_37_855 ();
 sg13g2_fill_8 FILLER_0_37_863 ();
 sg13g2_fill_8 FILLER_0_37_871 ();
 sg13g2_fill_8 FILLER_0_37_879 ();
 sg13g2_fill_8 FILLER_0_37_887 ();
 sg13g2_fill_8 FILLER_0_37_895 ();
 sg13g2_fill_8 FILLER_0_37_903 ();
 sg13g2_fill_8 FILLER_0_37_911 ();
 sg13g2_fill_8 FILLER_0_37_919 ();
 sg13g2_fill_8 FILLER_0_37_927 ();
 sg13g2_fill_8 FILLER_0_37_935 ();
 sg13g2_fill_8 FILLER_0_37_943 ();
 sg13g2_fill_8 FILLER_0_37_951 ();
 sg13g2_fill_8 FILLER_0_37_959 ();
 sg13g2_fill_8 FILLER_0_37_967 ();
 sg13g2_fill_8 FILLER_0_37_975 ();
 sg13g2_fill_8 FILLER_0_37_983 ();
 sg13g2_fill_8 FILLER_0_37_991 ();
 sg13g2_fill_8 FILLER_0_37_999 ();
 sg13g2_fill_8 FILLER_0_37_1007 ();
 sg13g2_fill_8 FILLER_0_37_1015 ();
 sg13g2_fill_8 FILLER_0_37_1023 ();
 sg13g2_fill_8 FILLER_0_37_1031 ();
 sg13g2_fill_8 FILLER_0_37_1039 ();
 sg13g2_fill_8 FILLER_0_37_1047 ();
 sg13g2_fill_8 FILLER_0_37_1055 ();
 sg13g2_fill_8 FILLER_0_37_1063 ();
 sg13g2_fill_8 FILLER_0_37_1071 ();
 sg13g2_fill_8 FILLER_0_37_1079 ();
 sg13g2_fill_8 FILLER_0_37_1087 ();
 sg13g2_fill_8 FILLER_0_37_1095 ();
 sg13g2_fill_8 FILLER_0_37_1103 ();
 sg13g2_fill_8 FILLER_0_37_1111 ();
 sg13g2_fill_8 FILLER_0_37_1119 ();
 sg13g2_fill_8 FILLER_0_37_1127 ();
 sg13g2_fill_8 FILLER_0_37_1135 ();
 sg13g2_fill_8 FILLER_0_37_1143 ();
 sg13g2_fill_8 FILLER_0_37_1151 ();
 sg13g2_fill_8 FILLER_0_37_1159 ();
 sg13g2_fill_8 FILLER_0_37_1167 ();
 sg13g2_fill_8 FILLER_0_37_1175 ();
 sg13g2_fill_8 FILLER_0_37_1183 ();
 sg13g2_fill_8 FILLER_0_37_1191 ();
 sg13g2_fill_8 FILLER_0_37_1199 ();
 sg13g2_fill_8 FILLER_0_37_1207 ();
 sg13g2_fill_8 FILLER_0_37_1215 ();
 sg13g2_fill_4 FILLER_0_37_1223 ();
 sg13g2_fill_1 FILLER_0_37_1227 ();
 sg13g2_fill_1 FILLER_0_38_0 ();
 sg13g2_fill_2 FILLER_0_38_37 ();
 sg13g2_fill_4 FILLER_0_38_49 ();
 sg13g2_decap_8 FILLER_0_38_58 ();
 sg13g2_fill_8 FILLER_0_38_79 ();
 sg13g2_fill_2 FILLER_0_38_113 ();
 sg13g2_fill_1 FILLER_0_38_115 ();
 sg13g2_fill_1 FILLER_0_38_121 ();
 sg13g2_fill_8 FILLER_0_38_153 ();
 sg13g2_fill_8 FILLER_0_38_161 ();
 sg13g2_fill_2 FILLER_0_38_169 ();
 sg13g2_fill_4 FILLER_0_38_175 ();
 sg13g2_fill_2 FILLER_0_38_208 ();
 sg13g2_fill_1 FILLER_0_38_210 ();
 sg13g2_fill_8 FILLER_0_38_215 ();
 sg13g2_fill_8 FILLER_0_38_223 ();
 sg13g2_fill_8 FILLER_0_38_231 ();
 sg13g2_fill_4 FILLER_0_38_263 ();
 sg13g2_fill_1 FILLER_0_38_267 ();
 sg13g2_fill_2 FILLER_0_38_313 ();
 sg13g2_fill_1 FILLER_0_38_315 ();
 sg13g2_fill_2 FILLER_0_38_326 ();
 sg13g2_fill_1 FILLER_0_38_328 ();
 sg13g2_fill_1 FILLER_0_38_365 ();
 sg13g2_fill_2 FILLER_0_38_397 ();
 sg13g2_fill_2 FILLER_0_38_439 ();
 sg13g2_fill_1 FILLER_0_38_441 ();
 sg13g2_fill_8 FILLER_0_38_451 ();
 sg13g2_decap_8 FILLER_0_38_459 ();
 sg13g2_fill_1 FILLER_0_38_478 ();
 sg13g2_decap_8 FILLER_0_38_501 ();
 sg13g2_fill_2 FILLER_0_38_544 ();
 sg13g2_fill_2 FILLER_0_38_568 ();
 sg13g2_fill_8 FILLER_0_38_627 ();
 sg13g2_fill_8 FILLER_0_38_635 ();
 sg13g2_fill_8 FILLER_0_38_643 ();
 sg13g2_fill_8 FILLER_0_38_651 ();
 sg13g2_fill_8 FILLER_0_38_659 ();
 sg13g2_fill_8 FILLER_0_38_667 ();
 sg13g2_fill_8 FILLER_0_38_675 ();
 sg13g2_fill_8 FILLER_0_38_683 ();
 sg13g2_fill_8 FILLER_0_38_691 ();
 sg13g2_fill_8 FILLER_0_38_699 ();
 sg13g2_fill_8 FILLER_0_38_707 ();
 sg13g2_fill_8 FILLER_0_38_715 ();
 sg13g2_fill_8 FILLER_0_38_723 ();
 sg13g2_fill_8 FILLER_0_38_731 ();
 sg13g2_fill_8 FILLER_0_38_739 ();
 sg13g2_fill_8 FILLER_0_38_747 ();
 sg13g2_fill_8 FILLER_0_38_755 ();
 sg13g2_fill_8 FILLER_0_38_763 ();
 sg13g2_fill_4 FILLER_0_38_771 ();
 sg13g2_fill_2 FILLER_0_38_775 ();
 sg13g2_fill_8 FILLER_0_38_781 ();
 sg13g2_fill_8 FILLER_0_38_789 ();
 sg13g2_fill_8 FILLER_0_38_797 ();
 sg13g2_fill_8 FILLER_0_38_805 ();
 sg13g2_fill_8 FILLER_0_38_813 ();
 sg13g2_fill_8 FILLER_0_38_821 ();
 sg13g2_fill_8 FILLER_0_38_829 ();
 sg13g2_fill_8 FILLER_0_38_837 ();
 sg13g2_fill_8 FILLER_0_38_845 ();
 sg13g2_fill_8 FILLER_0_38_853 ();
 sg13g2_fill_8 FILLER_0_38_861 ();
 sg13g2_fill_8 FILLER_0_38_869 ();
 sg13g2_fill_8 FILLER_0_38_877 ();
 sg13g2_fill_8 FILLER_0_38_885 ();
 sg13g2_fill_8 FILLER_0_38_893 ();
 sg13g2_fill_8 FILLER_0_38_901 ();
 sg13g2_fill_8 FILLER_0_38_909 ();
 sg13g2_fill_8 FILLER_0_38_917 ();
 sg13g2_fill_8 FILLER_0_38_925 ();
 sg13g2_fill_8 FILLER_0_38_933 ();
 sg13g2_fill_8 FILLER_0_38_941 ();
 sg13g2_fill_8 FILLER_0_38_949 ();
 sg13g2_fill_8 FILLER_0_38_957 ();
 sg13g2_fill_8 FILLER_0_38_965 ();
 sg13g2_fill_8 FILLER_0_38_973 ();
 sg13g2_fill_8 FILLER_0_38_981 ();
 sg13g2_fill_8 FILLER_0_38_989 ();
 sg13g2_fill_8 FILLER_0_38_997 ();
 sg13g2_fill_8 FILLER_0_38_1005 ();
 sg13g2_fill_8 FILLER_0_38_1013 ();
 sg13g2_fill_8 FILLER_0_38_1021 ();
 sg13g2_fill_8 FILLER_0_38_1029 ();
 sg13g2_fill_8 FILLER_0_38_1037 ();
 sg13g2_fill_8 FILLER_0_38_1045 ();
 sg13g2_fill_8 FILLER_0_38_1053 ();
 sg13g2_fill_8 FILLER_0_38_1061 ();
 sg13g2_fill_8 FILLER_0_38_1069 ();
 sg13g2_fill_8 FILLER_0_38_1077 ();
 sg13g2_fill_8 FILLER_0_38_1085 ();
 sg13g2_fill_8 FILLER_0_38_1093 ();
 sg13g2_fill_8 FILLER_0_38_1101 ();
 sg13g2_fill_8 FILLER_0_38_1109 ();
 sg13g2_fill_8 FILLER_0_38_1117 ();
 sg13g2_fill_8 FILLER_0_38_1125 ();
 sg13g2_fill_8 FILLER_0_38_1133 ();
 sg13g2_fill_8 FILLER_0_38_1141 ();
 sg13g2_fill_8 FILLER_0_38_1149 ();
 sg13g2_fill_8 FILLER_0_38_1157 ();
 sg13g2_fill_8 FILLER_0_38_1165 ();
 sg13g2_fill_8 FILLER_0_38_1173 ();
 sg13g2_fill_8 FILLER_0_38_1181 ();
 sg13g2_fill_8 FILLER_0_38_1189 ();
 sg13g2_fill_8 FILLER_0_38_1197 ();
 sg13g2_fill_8 FILLER_0_38_1205 ();
 sg13g2_fill_8 FILLER_0_38_1213 ();
 sg13g2_decap_8 FILLER_0_38_1221 ();
 sg13g2_fill_2 FILLER_0_39_0 ();
 sg13g2_fill_4 FILLER_0_39_28 ();
 sg13g2_fill_4 FILLER_0_39_119 ();
 sg13g2_fill_2 FILLER_0_39_123 ();
 sg13g2_fill_2 FILLER_0_39_130 ();
 sg13g2_fill_8 FILLER_0_39_140 ();
 sg13g2_fill_8 FILLER_0_39_148 ();
 sg13g2_fill_2 FILLER_0_39_156 ();
 sg13g2_fill_1 FILLER_0_39_188 ();
 sg13g2_fill_1 FILLER_0_39_220 ();
 sg13g2_fill_8 FILLER_0_39_261 ();
 sg13g2_fill_8 FILLER_0_39_269 ();
 sg13g2_fill_8 FILLER_0_39_277 ();
 sg13g2_fill_8 FILLER_0_39_285 ();
 sg13g2_fill_2 FILLER_0_39_293 ();
 sg13g2_fill_2 FILLER_0_39_307 ();
 sg13g2_fill_8 FILLER_0_39_313 ();
 sg13g2_fill_2 FILLER_0_39_326 ();
 sg13g2_fill_1 FILLER_0_39_338 ();
 sg13g2_fill_1 FILLER_0_39_349 ();
 sg13g2_fill_2 FILLER_0_39_376 ();
 sg13g2_fill_1 FILLER_0_39_378 ();
 sg13g2_fill_1 FILLER_0_39_383 ();
 sg13g2_fill_8 FILLER_0_39_388 ();
 sg13g2_fill_4 FILLER_0_39_396 ();
 sg13g2_fill_2 FILLER_0_39_400 ();
 sg13g2_fill_8 FILLER_0_39_410 ();
 sg13g2_fill_8 FILLER_0_39_418 ();
 sg13g2_fill_4 FILLER_0_39_426 ();
 sg13g2_fill_1 FILLER_0_39_430 ();
 sg13g2_fill_2 FILLER_0_39_475 ();
 sg13g2_fill_8 FILLER_0_39_508 ();
 sg13g2_fill_2 FILLER_0_39_516 ();
 sg13g2_fill_1 FILLER_0_39_523 ();
 sg13g2_fill_1 FILLER_0_39_528 ();
 sg13g2_fill_4 FILLER_0_39_533 ();
 sg13g2_fill_1 FILLER_0_39_537 ();
 sg13g2_fill_1 FILLER_0_39_564 ();
 sg13g2_fill_2 FILLER_0_39_594 ();
 sg13g2_fill_8 FILLER_0_39_620 ();
 sg13g2_fill_8 FILLER_0_39_628 ();
 sg13g2_fill_8 FILLER_0_39_636 ();
 sg13g2_fill_8 FILLER_0_39_644 ();
 sg13g2_fill_8 FILLER_0_39_652 ();
 sg13g2_fill_8 FILLER_0_39_660 ();
 sg13g2_fill_8 FILLER_0_39_668 ();
 sg13g2_fill_8 FILLER_0_39_676 ();
 sg13g2_fill_8 FILLER_0_39_684 ();
 sg13g2_fill_8 FILLER_0_39_692 ();
 sg13g2_fill_8 FILLER_0_39_700 ();
 sg13g2_fill_8 FILLER_0_39_708 ();
 sg13g2_fill_8 FILLER_0_39_716 ();
 sg13g2_fill_8 FILLER_0_39_724 ();
 sg13g2_fill_8 FILLER_0_39_732 ();
 sg13g2_fill_8 FILLER_0_39_740 ();
 sg13g2_fill_8 FILLER_0_39_748 ();
 sg13g2_fill_8 FILLER_0_39_756 ();
 sg13g2_fill_4 FILLER_0_39_764 ();
 sg13g2_fill_2 FILLER_0_39_768 ();
 sg13g2_fill_8 FILLER_0_39_822 ();
 sg13g2_fill_8 FILLER_0_39_830 ();
 sg13g2_fill_8 FILLER_0_39_838 ();
 sg13g2_fill_8 FILLER_0_39_846 ();
 sg13g2_fill_8 FILLER_0_39_854 ();
 sg13g2_fill_8 FILLER_0_39_862 ();
 sg13g2_fill_8 FILLER_0_39_870 ();
 sg13g2_fill_8 FILLER_0_39_878 ();
 sg13g2_fill_8 FILLER_0_39_886 ();
 sg13g2_fill_8 FILLER_0_39_894 ();
 sg13g2_fill_8 FILLER_0_39_902 ();
 sg13g2_fill_8 FILLER_0_39_910 ();
 sg13g2_fill_8 FILLER_0_39_918 ();
 sg13g2_fill_8 FILLER_0_39_926 ();
 sg13g2_fill_8 FILLER_0_39_934 ();
 sg13g2_fill_8 FILLER_0_39_942 ();
 sg13g2_fill_8 FILLER_0_39_950 ();
 sg13g2_fill_8 FILLER_0_39_958 ();
 sg13g2_fill_8 FILLER_0_39_966 ();
 sg13g2_fill_8 FILLER_0_39_974 ();
 sg13g2_fill_8 FILLER_0_39_982 ();
 sg13g2_fill_8 FILLER_0_39_990 ();
 sg13g2_fill_8 FILLER_0_39_998 ();
 sg13g2_fill_8 FILLER_0_39_1006 ();
 sg13g2_fill_8 FILLER_0_39_1014 ();
 sg13g2_fill_8 FILLER_0_39_1022 ();
 sg13g2_fill_8 FILLER_0_39_1030 ();
 sg13g2_fill_8 FILLER_0_39_1038 ();
 sg13g2_fill_8 FILLER_0_39_1046 ();
 sg13g2_fill_8 FILLER_0_39_1054 ();
 sg13g2_fill_8 FILLER_0_39_1062 ();
 sg13g2_fill_8 FILLER_0_39_1070 ();
 sg13g2_fill_8 FILLER_0_39_1078 ();
 sg13g2_fill_8 FILLER_0_39_1086 ();
 sg13g2_fill_8 FILLER_0_39_1094 ();
 sg13g2_fill_8 FILLER_0_39_1102 ();
 sg13g2_fill_8 FILLER_0_39_1110 ();
 sg13g2_fill_8 FILLER_0_39_1118 ();
 sg13g2_fill_8 FILLER_0_39_1126 ();
 sg13g2_fill_8 FILLER_0_39_1134 ();
 sg13g2_fill_8 FILLER_0_39_1142 ();
 sg13g2_fill_8 FILLER_0_39_1150 ();
 sg13g2_fill_8 FILLER_0_39_1158 ();
 sg13g2_fill_8 FILLER_0_39_1166 ();
 sg13g2_fill_8 FILLER_0_39_1174 ();
 sg13g2_fill_8 FILLER_0_39_1182 ();
 sg13g2_fill_8 FILLER_0_39_1190 ();
 sg13g2_fill_8 FILLER_0_39_1198 ();
 sg13g2_fill_8 FILLER_0_39_1206 ();
 sg13g2_fill_8 FILLER_0_39_1214 ();
 sg13g2_fill_4 FILLER_0_39_1222 ();
 sg13g2_fill_2 FILLER_0_39_1226 ();
 sg13g2_fill_8 FILLER_0_40_0 ();
 sg13g2_fill_1 FILLER_0_40_8 ();
 sg13g2_fill_8 FILLER_0_40_13 ();
 sg13g2_fill_2 FILLER_0_40_21 ();
 sg13g2_fill_8 FILLER_0_40_33 ();
 sg13g2_fill_2 FILLER_0_40_50 ();
 sg13g2_fill_4 FILLER_0_40_61 ();
 sg13g2_fill_8 FILLER_0_40_79 ();
 sg13g2_fill_4 FILLER_0_40_87 ();
 sg13g2_fill_1 FILLER_0_40_91 ();
 sg13g2_fill_4 FILLER_0_40_96 ();
 sg13g2_fill_2 FILLER_0_40_100 ();
 sg13g2_fill_1 FILLER_0_40_117 ();
 sg13g2_fill_2 FILLER_0_40_154 ();
 sg13g2_fill_1 FILLER_0_40_156 ();
 sg13g2_fill_1 FILLER_0_40_192 ();
 sg13g2_fill_4 FILLER_0_40_224 ();
 sg13g2_fill_2 FILLER_0_40_228 ();
 sg13g2_fill_1 FILLER_0_40_235 ();
 sg13g2_fill_1 FILLER_0_40_241 ();
 sg13g2_fill_2 FILLER_0_40_268 ();
 sg13g2_fill_1 FILLER_0_40_296 ();
 sg13g2_fill_2 FILLER_0_40_307 ();
 sg13g2_fill_8 FILLER_0_40_324 ();
 sg13g2_fill_8 FILLER_0_40_332 ();
 sg13g2_fill_1 FILLER_0_40_340 ();
 sg13g2_fill_8 FILLER_0_40_345 ();
 sg13g2_fill_4 FILLER_0_40_353 ();
 sg13g2_fill_1 FILLER_0_40_357 ();
 sg13g2_fill_8 FILLER_0_40_362 ();
 sg13g2_fill_8 FILLER_0_40_370 ();
 sg13g2_fill_8 FILLER_0_40_378 ();
 sg13g2_fill_8 FILLER_0_40_394 ();
 sg13g2_fill_4 FILLER_0_40_402 ();
 sg13g2_fill_2 FILLER_0_40_406 ();
 sg13g2_decap_8 FILLER_0_40_449 ();
 sg13g2_fill_8 FILLER_0_40_482 ();
 sg13g2_fill_4 FILLER_0_40_490 ();
 sg13g2_fill_8 FILLER_0_40_499 ();
 sg13g2_fill_8 FILLER_0_40_507 ();
 sg13g2_fill_1 FILLER_0_40_515 ();
 sg13g2_fill_8 FILLER_0_40_520 ();
 sg13g2_fill_8 FILLER_0_40_528 ();
 sg13g2_fill_8 FILLER_0_40_536 ();
 sg13g2_fill_1 FILLER_0_40_544 ();
 sg13g2_fill_1 FILLER_0_40_549 ();
 sg13g2_fill_8 FILLER_0_40_569 ();
 sg13g2_decap_8 FILLER_0_40_577 ();
 sg13g2_fill_8 FILLER_0_40_596 ();
 sg13g2_fill_2 FILLER_0_40_604 ();
 sg13g2_fill_8 FILLER_0_40_616 ();
 sg13g2_fill_8 FILLER_0_40_624 ();
 sg13g2_fill_8 FILLER_0_40_632 ();
 sg13g2_fill_8 FILLER_0_40_640 ();
 sg13g2_fill_8 FILLER_0_40_648 ();
 sg13g2_fill_8 FILLER_0_40_656 ();
 sg13g2_fill_8 FILLER_0_40_664 ();
 sg13g2_fill_8 FILLER_0_40_672 ();
 sg13g2_fill_8 FILLER_0_40_680 ();
 sg13g2_fill_8 FILLER_0_40_688 ();
 sg13g2_fill_8 FILLER_0_40_696 ();
 sg13g2_fill_8 FILLER_0_40_704 ();
 sg13g2_fill_4 FILLER_0_40_712 ();
 sg13g2_fill_1 FILLER_0_40_716 ();
 sg13g2_fill_8 FILLER_0_40_727 ();
 sg13g2_fill_8 FILLER_0_40_735 ();
 sg13g2_fill_4 FILLER_0_40_743 ();
 sg13g2_fill_1 FILLER_0_40_747 ();
 sg13g2_fill_8 FILLER_0_40_752 ();
 sg13g2_fill_8 FILLER_0_40_760 ();
 sg13g2_fill_2 FILLER_0_40_768 ();
 sg13g2_fill_4 FILLER_0_40_775 ();
 sg13g2_fill_1 FILLER_0_40_779 ();
 sg13g2_fill_8 FILLER_0_40_814 ();
 sg13g2_fill_1 FILLER_0_40_822 ();
 sg13g2_fill_8 FILLER_0_40_849 ();
 sg13g2_fill_8 FILLER_0_40_857 ();
 sg13g2_fill_8 FILLER_0_40_865 ();
 sg13g2_fill_8 FILLER_0_40_873 ();
 sg13g2_fill_8 FILLER_0_40_881 ();
 sg13g2_fill_8 FILLER_0_40_889 ();
 sg13g2_fill_8 FILLER_0_40_897 ();
 sg13g2_fill_8 FILLER_0_40_905 ();
 sg13g2_fill_8 FILLER_0_40_913 ();
 sg13g2_fill_8 FILLER_0_40_921 ();
 sg13g2_fill_8 FILLER_0_40_929 ();
 sg13g2_fill_8 FILLER_0_40_937 ();
 sg13g2_fill_8 FILLER_0_40_945 ();
 sg13g2_fill_8 FILLER_0_40_953 ();
 sg13g2_fill_8 FILLER_0_40_961 ();
 sg13g2_fill_8 FILLER_0_40_969 ();
 sg13g2_fill_8 FILLER_0_40_977 ();
 sg13g2_fill_8 FILLER_0_40_985 ();
 sg13g2_fill_8 FILLER_0_40_993 ();
 sg13g2_fill_8 FILLER_0_40_1001 ();
 sg13g2_fill_8 FILLER_0_40_1009 ();
 sg13g2_fill_8 FILLER_0_40_1017 ();
 sg13g2_fill_8 FILLER_0_40_1025 ();
 sg13g2_fill_8 FILLER_0_40_1033 ();
 sg13g2_fill_8 FILLER_0_40_1041 ();
 sg13g2_fill_8 FILLER_0_40_1049 ();
 sg13g2_fill_8 FILLER_0_40_1057 ();
 sg13g2_fill_8 FILLER_0_40_1065 ();
 sg13g2_fill_8 FILLER_0_40_1073 ();
 sg13g2_fill_8 FILLER_0_40_1081 ();
 sg13g2_fill_8 FILLER_0_40_1089 ();
 sg13g2_fill_8 FILLER_0_40_1097 ();
 sg13g2_fill_8 FILLER_0_40_1105 ();
 sg13g2_fill_8 FILLER_0_40_1113 ();
 sg13g2_fill_8 FILLER_0_40_1121 ();
 sg13g2_fill_8 FILLER_0_40_1129 ();
 sg13g2_fill_8 FILLER_0_40_1137 ();
 sg13g2_fill_8 FILLER_0_40_1145 ();
 sg13g2_fill_8 FILLER_0_40_1153 ();
 sg13g2_fill_8 FILLER_0_40_1161 ();
 sg13g2_fill_8 FILLER_0_40_1169 ();
 sg13g2_fill_8 FILLER_0_40_1177 ();
 sg13g2_fill_8 FILLER_0_40_1185 ();
 sg13g2_fill_8 FILLER_0_40_1193 ();
 sg13g2_fill_8 FILLER_0_40_1201 ();
 sg13g2_fill_8 FILLER_0_40_1209 ();
 sg13g2_fill_8 FILLER_0_40_1217 ();
 sg13g2_fill_2 FILLER_0_40_1225 ();
 sg13g2_fill_1 FILLER_0_40_1227 ();
 sg13g2_fill_8 FILLER_0_41_0 ();
 sg13g2_fill_8 FILLER_0_41_8 ();
 sg13g2_fill_1 FILLER_0_41_16 ();
 sg13g2_fill_4 FILLER_0_41_22 ();
 sg13g2_fill_8 FILLER_0_41_36 ();
 sg13g2_fill_4 FILLER_0_41_44 ();
 sg13g2_fill_4 FILLER_0_41_53 ();
 sg13g2_fill_2 FILLER_0_41_57 ();
 sg13g2_fill_1 FILLER_0_41_121 ();
 sg13g2_fill_8 FILLER_0_41_126 ();
 sg13g2_fill_1 FILLER_0_41_134 ();
 sg13g2_fill_8 FILLER_0_41_139 ();
 sg13g2_fill_1 FILLER_0_41_147 ();
 sg13g2_fill_4 FILLER_0_41_158 ();
 sg13g2_fill_1 FILLER_0_41_162 ();
 sg13g2_fill_1 FILLER_0_41_178 ();
 sg13g2_fill_1 FILLER_0_41_189 ();
 sg13g2_fill_1 FILLER_0_41_200 ();
 sg13g2_fill_2 FILLER_0_41_211 ();
 sg13g2_decap_8 FILLER_0_41_217 ();
 sg13g2_fill_2 FILLER_0_41_284 ();
 sg13g2_fill_2 FILLER_0_41_312 ();
 sg13g2_fill_1 FILLER_0_41_314 ();
 sg13g2_fill_2 FILLER_0_41_341 ();
 sg13g2_fill_1 FILLER_0_41_343 ();
 sg13g2_fill_2 FILLER_0_41_349 ();
 sg13g2_fill_4 FILLER_0_41_361 ();
 sg13g2_fill_8 FILLER_0_41_396 ();
 sg13g2_decap_8 FILLER_0_41_404 ();
 sg13g2_fill_1 FILLER_0_41_420 ();
 sg13g2_fill_1 FILLER_0_41_452 ();
 sg13g2_fill_4 FILLER_0_41_457 ();
 sg13g2_fill_8 FILLER_0_41_465 ();
 sg13g2_fill_2 FILLER_0_41_473 ();
 sg13g2_fill_1 FILLER_0_41_475 ();
 sg13g2_fill_2 FILLER_0_41_506 ();
 sg13g2_fill_1 FILLER_0_41_508 ();
 sg13g2_fill_8 FILLER_0_41_535 ();
 sg13g2_decap_8 FILLER_0_41_573 ();
 sg13g2_fill_8 FILLER_0_41_584 ();
 sg13g2_fill_8 FILLER_0_41_592 ();
 sg13g2_fill_2 FILLER_0_41_600 ();
 sg13g2_fill_8 FILLER_0_41_633 ();
 sg13g2_fill_8 FILLER_0_41_641 ();
 sg13g2_fill_8 FILLER_0_41_649 ();
 sg13g2_fill_8 FILLER_0_41_657 ();
 sg13g2_fill_8 FILLER_0_41_665 ();
 sg13g2_fill_8 FILLER_0_41_673 ();
 sg13g2_fill_8 FILLER_0_41_681 ();
 sg13g2_fill_8 FILLER_0_41_689 ();
 sg13g2_fill_2 FILLER_0_41_697 ();
 sg13g2_fill_1 FILLER_0_41_699 ();
 sg13g2_fill_4 FILLER_0_41_772 ();
 sg13g2_fill_2 FILLER_0_41_827 ();
 sg13g2_fill_8 FILLER_0_41_833 ();
 sg13g2_fill_8 FILLER_0_41_841 ();
 sg13g2_fill_8 FILLER_0_41_849 ();
 sg13g2_fill_8 FILLER_0_41_857 ();
 sg13g2_fill_8 FILLER_0_41_865 ();
 sg13g2_fill_8 FILLER_0_41_873 ();
 sg13g2_fill_8 FILLER_0_41_881 ();
 sg13g2_fill_8 FILLER_0_41_889 ();
 sg13g2_fill_8 FILLER_0_41_897 ();
 sg13g2_fill_8 FILLER_0_41_905 ();
 sg13g2_fill_8 FILLER_0_41_913 ();
 sg13g2_fill_8 FILLER_0_41_921 ();
 sg13g2_fill_8 FILLER_0_41_929 ();
 sg13g2_fill_8 FILLER_0_41_937 ();
 sg13g2_fill_8 FILLER_0_41_945 ();
 sg13g2_fill_8 FILLER_0_41_953 ();
 sg13g2_fill_8 FILLER_0_41_961 ();
 sg13g2_fill_8 FILLER_0_41_969 ();
 sg13g2_fill_8 FILLER_0_41_977 ();
 sg13g2_fill_8 FILLER_0_41_985 ();
 sg13g2_fill_8 FILLER_0_41_993 ();
 sg13g2_fill_8 FILLER_0_41_1001 ();
 sg13g2_fill_8 FILLER_0_41_1009 ();
 sg13g2_fill_8 FILLER_0_41_1017 ();
 sg13g2_fill_8 FILLER_0_41_1025 ();
 sg13g2_fill_8 FILLER_0_41_1033 ();
 sg13g2_fill_8 FILLER_0_41_1041 ();
 sg13g2_fill_8 FILLER_0_41_1049 ();
 sg13g2_fill_8 FILLER_0_41_1057 ();
 sg13g2_fill_8 FILLER_0_41_1065 ();
 sg13g2_fill_8 FILLER_0_41_1073 ();
 sg13g2_fill_8 FILLER_0_41_1081 ();
 sg13g2_fill_8 FILLER_0_41_1089 ();
 sg13g2_fill_8 FILLER_0_41_1097 ();
 sg13g2_fill_8 FILLER_0_41_1105 ();
 sg13g2_fill_8 FILLER_0_41_1113 ();
 sg13g2_fill_8 FILLER_0_41_1121 ();
 sg13g2_fill_8 FILLER_0_41_1129 ();
 sg13g2_fill_8 FILLER_0_41_1137 ();
 sg13g2_fill_8 FILLER_0_41_1145 ();
 sg13g2_fill_8 FILLER_0_41_1153 ();
 sg13g2_fill_8 FILLER_0_41_1161 ();
 sg13g2_fill_8 FILLER_0_41_1169 ();
 sg13g2_fill_8 FILLER_0_41_1177 ();
 sg13g2_fill_8 FILLER_0_41_1185 ();
 sg13g2_fill_8 FILLER_0_41_1193 ();
 sg13g2_fill_8 FILLER_0_41_1201 ();
 sg13g2_fill_8 FILLER_0_41_1209 ();
 sg13g2_fill_8 FILLER_0_41_1217 ();
 sg13g2_fill_2 FILLER_0_41_1225 ();
 sg13g2_fill_1 FILLER_0_41_1227 ();
 sg13g2_decap_8 FILLER_0_42_0 ();
 sg13g2_fill_2 FILLER_0_42_20 ();
 sg13g2_fill_2 FILLER_0_42_48 ();
 sg13g2_fill_8 FILLER_0_42_72 ();
 sg13g2_fill_4 FILLER_0_42_80 ();
 sg13g2_fill_2 FILLER_0_42_84 ();
 sg13g2_fill_2 FILLER_0_42_136 ();
 sg13g2_fill_4 FILLER_0_42_142 ();
 sg13g2_decap_8 FILLER_0_42_176 ();
 sg13g2_decap_8 FILLER_0_42_193 ();
 sg13g2_fill_8 FILLER_0_42_212 ();
 sg13g2_fill_8 FILLER_0_42_220 ();
 sg13g2_fill_2 FILLER_0_42_228 ();
 sg13g2_fill_1 FILLER_0_42_230 ();
 sg13g2_fill_1 FILLER_0_42_255 ();
 sg13g2_fill_1 FILLER_0_42_271 ();
 sg13g2_fill_1 FILLER_0_42_282 ();
 sg13g2_fill_1 FILLER_0_42_288 ();
 sg13g2_fill_1 FILLER_0_42_297 ();
 sg13g2_fill_1 FILLER_0_42_308 ();
 sg13g2_fill_1 FILLER_0_42_335 ();
 sg13g2_fill_2 FILLER_0_42_340 ();
 sg13g2_fill_1 FILLER_0_42_342 ();
 sg13g2_fill_2 FILLER_0_42_405 ();
 sg13g2_fill_8 FILLER_0_42_445 ();
 sg13g2_fill_8 FILLER_0_42_453 ();
 sg13g2_fill_8 FILLER_0_42_461 ();
 sg13g2_fill_2 FILLER_0_42_469 ();
 sg13g2_fill_1 FILLER_0_42_471 ();
 sg13g2_fill_1 FILLER_0_42_476 ();
 sg13g2_fill_2 FILLER_0_42_522 ();
 sg13g2_fill_1 FILLER_0_42_524 ();
 sg13g2_fill_2 FILLER_0_42_589 ();
 sg13g2_fill_2 FILLER_0_42_601 ();
 sg13g2_fill_1 FILLER_0_42_603 ();
 sg13g2_fill_8 FILLER_0_42_618 ();
 sg13g2_fill_8 FILLER_0_42_626 ();
 sg13g2_fill_2 FILLER_0_42_634 ();
 sg13g2_fill_1 FILLER_0_42_636 ();
 sg13g2_fill_8 FILLER_0_42_641 ();
 sg13g2_fill_8 FILLER_0_42_649 ();
 sg13g2_fill_8 FILLER_0_42_657 ();
 sg13g2_fill_8 FILLER_0_42_665 ();
 sg13g2_fill_8 FILLER_0_42_673 ();
 sg13g2_fill_8 FILLER_0_42_681 ();
 sg13g2_decap_8 FILLER_0_42_689 ();
 sg13g2_fill_1 FILLER_0_42_722 ();
 sg13g2_fill_2 FILLER_0_42_727 ();
 sg13g2_fill_1 FILLER_0_42_755 ();
 sg13g2_fill_4 FILLER_0_42_786 ();
 sg13g2_fill_8 FILLER_0_42_795 ();
 sg13g2_fill_4 FILLER_0_42_803 ();
 sg13g2_fill_8 FILLER_0_42_843 ();
 sg13g2_fill_8 FILLER_0_42_851 ();
 sg13g2_fill_8 FILLER_0_42_859 ();
 sg13g2_fill_8 FILLER_0_42_867 ();
 sg13g2_fill_8 FILLER_0_42_875 ();
 sg13g2_fill_8 FILLER_0_42_883 ();
 sg13g2_fill_8 FILLER_0_42_891 ();
 sg13g2_fill_8 FILLER_0_42_899 ();
 sg13g2_fill_8 FILLER_0_42_907 ();
 sg13g2_fill_8 FILLER_0_42_915 ();
 sg13g2_fill_8 FILLER_0_42_923 ();
 sg13g2_fill_8 FILLER_0_42_931 ();
 sg13g2_fill_8 FILLER_0_42_939 ();
 sg13g2_fill_8 FILLER_0_42_947 ();
 sg13g2_fill_8 FILLER_0_42_955 ();
 sg13g2_fill_8 FILLER_0_42_963 ();
 sg13g2_fill_8 FILLER_0_42_971 ();
 sg13g2_fill_8 FILLER_0_42_979 ();
 sg13g2_fill_8 FILLER_0_42_987 ();
 sg13g2_fill_8 FILLER_0_42_995 ();
 sg13g2_fill_8 FILLER_0_42_1003 ();
 sg13g2_fill_8 FILLER_0_42_1011 ();
 sg13g2_fill_8 FILLER_0_42_1019 ();
 sg13g2_fill_8 FILLER_0_42_1027 ();
 sg13g2_fill_8 FILLER_0_42_1035 ();
 sg13g2_fill_8 FILLER_0_42_1043 ();
 sg13g2_fill_8 FILLER_0_42_1051 ();
 sg13g2_fill_8 FILLER_0_42_1059 ();
 sg13g2_fill_8 FILLER_0_42_1067 ();
 sg13g2_fill_8 FILLER_0_42_1075 ();
 sg13g2_fill_8 FILLER_0_42_1083 ();
 sg13g2_fill_8 FILLER_0_42_1091 ();
 sg13g2_fill_8 FILLER_0_42_1099 ();
 sg13g2_fill_8 FILLER_0_42_1107 ();
 sg13g2_fill_8 FILLER_0_42_1115 ();
 sg13g2_fill_8 FILLER_0_42_1123 ();
 sg13g2_fill_8 FILLER_0_42_1131 ();
 sg13g2_fill_8 FILLER_0_42_1139 ();
 sg13g2_fill_8 FILLER_0_42_1147 ();
 sg13g2_fill_8 FILLER_0_42_1155 ();
 sg13g2_fill_8 FILLER_0_42_1163 ();
 sg13g2_fill_8 FILLER_0_42_1171 ();
 sg13g2_fill_8 FILLER_0_42_1179 ();
 sg13g2_fill_8 FILLER_0_42_1187 ();
 sg13g2_fill_8 FILLER_0_42_1195 ();
 sg13g2_fill_8 FILLER_0_42_1203 ();
 sg13g2_fill_8 FILLER_0_42_1211 ();
 sg13g2_fill_8 FILLER_0_42_1219 ();
 sg13g2_fill_1 FILLER_0_42_1227 ();
 sg13g2_fill_2 FILLER_0_43_0 ();
 sg13g2_fill_1 FILLER_0_43_2 ();
 sg13g2_fill_2 FILLER_0_43_29 ();
 sg13g2_fill_8 FILLER_0_43_83 ();
 sg13g2_fill_1 FILLER_0_43_91 ();
 sg13g2_fill_1 FILLER_0_43_96 ();
 sg13g2_fill_1 FILLER_0_43_102 ();
 sg13g2_fill_1 FILLER_0_43_129 ();
 sg13g2_fill_1 FILLER_0_43_164 ();
 sg13g2_fill_1 FILLER_0_43_169 ();
 sg13g2_fill_8 FILLER_0_43_201 ();
 sg13g2_decap_8 FILLER_0_43_209 ();
 sg13g2_fill_8 FILLER_0_43_221 ();
 sg13g2_fill_8 FILLER_0_43_229 ();
 sg13g2_fill_8 FILLER_0_43_237 ();
 sg13g2_fill_4 FILLER_0_43_245 ();
 sg13g2_fill_1 FILLER_0_43_249 ();
 sg13g2_fill_4 FILLER_0_43_259 ();
 sg13g2_fill_2 FILLER_0_43_263 ();
 sg13g2_fill_4 FILLER_0_43_269 ();
 sg13g2_fill_2 FILLER_0_43_278 ();
 sg13g2_fill_8 FILLER_0_43_284 ();
 sg13g2_fill_2 FILLER_0_43_292 ();
 sg13g2_fill_8 FILLER_0_43_298 ();
 sg13g2_fill_4 FILLER_0_43_311 ();
 sg13g2_fill_1 FILLER_0_43_319 ();
 sg13g2_fill_1 FILLER_0_43_362 ();
 sg13g2_fill_1 FILLER_0_43_367 ();
 sg13g2_fill_2 FILLER_0_43_378 ();
 sg13g2_fill_1 FILLER_0_43_380 ();
 sg13g2_fill_8 FILLER_0_43_435 ();
 sg13g2_fill_8 FILLER_0_43_443 ();
 sg13g2_fill_8 FILLER_0_43_455 ();
 sg13g2_fill_4 FILLER_0_43_463 ();
 sg13g2_fill_2 FILLER_0_43_467 ();
 sg13g2_fill_2 FILLER_0_43_481 ();
 sg13g2_fill_1 FILLER_0_43_483 ();
 sg13g2_fill_1 FILLER_0_43_489 ();
 sg13g2_fill_2 FILLER_0_43_494 ();
 sg13g2_fill_1 FILLER_0_43_506 ();
 sg13g2_fill_8 FILLER_0_43_540 ();
 sg13g2_decap_8 FILLER_0_43_548 ();
 sg13g2_fill_2 FILLER_0_43_602 ();
 sg13g2_fill_8 FILLER_0_43_656 ();
 sg13g2_fill_8 FILLER_0_43_664 ();
 sg13g2_fill_8 FILLER_0_43_672 ();
 sg13g2_fill_8 FILLER_0_43_680 ();
 sg13g2_fill_8 FILLER_0_43_688 ();
 sg13g2_fill_4 FILLER_0_43_700 ();
 sg13g2_fill_4 FILLER_0_43_708 ();
 sg13g2_fill_1 FILLER_0_43_712 ();
 sg13g2_fill_2 FILLER_0_43_723 ();
 sg13g2_fill_1 FILLER_0_43_725 ();
 sg13g2_fill_2 FILLER_0_43_755 ();
 sg13g2_fill_1 FILLER_0_43_757 ();
 sg13g2_fill_4 FILLER_0_43_780 ();
 sg13g2_fill_2 FILLER_0_43_818 ();
 sg13g2_fill_1 FILLER_0_43_820 ();
 sg13g2_fill_8 FILLER_0_43_866 ();
 sg13g2_fill_8 FILLER_0_43_874 ();
 sg13g2_fill_8 FILLER_0_43_882 ();
 sg13g2_fill_8 FILLER_0_43_890 ();
 sg13g2_fill_8 FILLER_0_43_898 ();
 sg13g2_fill_8 FILLER_0_43_906 ();
 sg13g2_fill_8 FILLER_0_43_914 ();
 sg13g2_fill_8 FILLER_0_43_922 ();
 sg13g2_fill_8 FILLER_0_43_930 ();
 sg13g2_fill_8 FILLER_0_43_938 ();
 sg13g2_fill_8 FILLER_0_43_946 ();
 sg13g2_fill_8 FILLER_0_43_954 ();
 sg13g2_fill_8 FILLER_0_43_962 ();
 sg13g2_fill_8 FILLER_0_43_970 ();
 sg13g2_fill_8 FILLER_0_43_978 ();
 sg13g2_fill_8 FILLER_0_43_986 ();
 sg13g2_fill_8 FILLER_0_43_994 ();
 sg13g2_fill_8 FILLER_0_43_1002 ();
 sg13g2_fill_8 FILLER_0_43_1010 ();
 sg13g2_fill_8 FILLER_0_43_1018 ();
 sg13g2_fill_8 FILLER_0_43_1026 ();
 sg13g2_fill_8 FILLER_0_43_1034 ();
 sg13g2_fill_8 FILLER_0_43_1042 ();
 sg13g2_fill_8 FILLER_0_43_1050 ();
 sg13g2_fill_8 FILLER_0_43_1058 ();
 sg13g2_fill_8 FILLER_0_43_1066 ();
 sg13g2_fill_8 FILLER_0_43_1074 ();
 sg13g2_fill_8 FILLER_0_43_1082 ();
 sg13g2_fill_8 FILLER_0_43_1090 ();
 sg13g2_fill_8 FILLER_0_43_1098 ();
 sg13g2_fill_8 FILLER_0_43_1106 ();
 sg13g2_fill_8 FILLER_0_43_1114 ();
 sg13g2_fill_8 FILLER_0_43_1122 ();
 sg13g2_fill_8 FILLER_0_43_1130 ();
 sg13g2_fill_8 FILLER_0_43_1138 ();
 sg13g2_fill_8 FILLER_0_43_1146 ();
 sg13g2_fill_8 FILLER_0_43_1154 ();
 sg13g2_fill_8 FILLER_0_43_1162 ();
 sg13g2_fill_8 FILLER_0_43_1170 ();
 sg13g2_fill_8 FILLER_0_43_1178 ();
 sg13g2_fill_8 FILLER_0_43_1186 ();
 sg13g2_fill_8 FILLER_0_43_1194 ();
 sg13g2_fill_8 FILLER_0_43_1202 ();
 sg13g2_fill_8 FILLER_0_43_1210 ();
 sg13g2_fill_8 FILLER_0_43_1218 ();
 sg13g2_fill_2 FILLER_0_43_1226 ();
 sg13g2_fill_1 FILLER_0_44_0 ();
 sg13g2_fill_1 FILLER_0_44_37 ();
 sg13g2_fill_1 FILLER_0_44_48 ();
 sg13g2_fill_1 FILLER_0_44_67 ();
 sg13g2_fill_8 FILLER_0_44_82 ();
 sg13g2_fill_8 FILLER_0_44_90 ();
 sg13g2_fill_2 FILLER_0_44_98 ();
 sg13g2_fill_1 FILLER_0_44_100 ();
 sg13g2_fill_2 FILLER_0_44_105 ();
 sg13g2_fill_2 FILLER_0_44_117 ();
 sg13g2_fill_1 FILLER_0_44_129 ();
 sg13g2_fill_2 FILLER_0_44_135 ();
 sg13g2_fill_2 FILLER_0_44_141 ();
 sg13g2_fill_1 FILLER_0_44_143 ();
 sg13g2_fill_2 FILLER_0_44_153 ();
 sg13g2_fill_2 FILLER_0_44_193 ();
 sg13g2_fill_1 FILLER_0_44_195 ();
 sg13g2_fill_1 FILLER_0_44_204 ();
 sg13g2_fill_8 FILLER_0_44_236 ();
 sg13g2_fill_8 FILLER_0_44_244 ();
 sg13g2_fill_8 FILLER_0_44_252 ();
 sg13g2_fill_2 FILLER_0_44_260 ();
 sg13g2_fill_8 FILLER_0_44_276 ();
 sg13g2_fill_8 FILLER_0_44_284 ();
 sg13g2_fill_2 FILLER_0_44_292 ();
 sg13g2_fill_8 FILLER_0_44_317 ();
 sg13g2_fill_8 FILLER_0_44_325 ();
 sg13g2_fill_8 FILLER_0_44_333 ();
 sg13g2_fill_1 FILLER_0_44_350 ();
 sg13g2_fill_8 FILLER_0_44_361 ();
 sg13g2_fill_8 FILLER_0_44_369 ();
 sg13g2_fill_4 FILLER_0_44_385 ();
 sg13g2_fill_1 FILLER_0_44_389 ();
 sg13g2_fill_8 FILLER_0_44_433 ();
 sg13g2_fill_4 FILLER_0_44_441 ();
 sg13g2_fill_4 FILLER_0_44_481 ();
 sg13g2_fill_4 FILLER_0_44_516 ();
 sg13g2_fill_8 FILLER_0_44_550 ();
 sg13g2_fill_8 FILLER_0_44_558 ();
 sg13g2_fill_2 FILLER_0_44_566 ();
 sg13g2_fill_1 FILLER_0_44_588 ();
 sg13g2_fill_1 FILLER_0_44_609 ();
 sg13g2_fill_8 FILLER_0_44_619 ();
 sg13g2_fill_8 FILLER_0_44_627 ();
 sg13g2_fill_8 FILLER_0_44_635 ();
 sg13g2_fill_8 FILLER_0_44_643 ();
 sg13g2_fill_8 FILLER_0_44_651 ();
 sg13g2_fill_8 FILLER_0_44_659 ();
 sg13g2_fill_8 FILLER_0_44_667 ();
 sg13g2_fill_8 FILLER_0_44_675 ();
 sg13g2_fill_4 FILLER_0_44_683 ();
 sg13g2_fill_8 FILLER_0_44_728 ();
 sg13g2_fill_8 FILLER_0_44_736 ();
 sg13g2_fill_8 FILLER_0_44_744 ();
 sg13g2_fill_8 FILLER_0_44_771 ();
 sg13g2_fill_4 FILLER_0_44_779 ();
 sg13g2_fill_1 FILLER_0_44_788 ();
 sg13g2_fill_8 FILLER_0_44_803 ();
 sg13g2_fill_4 FILLER_0_44_811 ();
 sg13g2_fill_2 FILLER_0_44_815 ();
 sg13g2_fill_4 FILLER_0_44_821 ();
 sg13g2_fill_1 FILLER_0_44_825 ();
 sg13g2_fill_4 FILLER_0_44_831 ();
 sg13g2_fill_2 FILLER_0_44_835 ();
 sg13g2_fill_4 FILLER_0_44_841 ();
 sg13g2_fill_8 FILLER_0_44_881 ();
 sg13g2_fill_8 FILLER_0_44_889 ();
 sg13g2_fill_8 FILLER_0_44_897 ();
 sg13g2_fill_8 FILLER_0_44_905 ();
 sg13g2_fill_8 FILLER_0_44_913 ();
 sg13g2_fill_8 FILLER_0_44_921 ();
 sg13g2_fill_8 FILLER_0_44_929 ();
 sg13g2_fill_8 FILLER_0_44_937 ();
 sg13g2_fill_8 FILLER_0_44_945 ();
 sg13g2_fill_8 FILLER_0_44_953 ();
 sg13g2_fill_8 FILLER_0_44_961 ();
 sg13g2_fill_8 FILLER_0_44_969 ();
 sg13g2_fill_8 FILLER_0_44_977 ();
 sg13g2_fill_8 FILLER_0_44_985 ();
 sg13g2_fill_8 FILLER_0_44_993 ();
 sg13g2_fill_8 FILLER_0_44_1001 ();
 sg13g2_fill_8 FILLER_0_44_1009 ();
 sg13g2_fill_8 FILLER_0_44_1017 ();
 sg13g2_fill_8 FILLER_0_44_1025 ();
 sg13g2_fill_8 FILLER_0_44_1033 ();
 sg13g2_fill_8 FILLER_0_44_1041 ();
 sg13g2_fill_8 FILLER_0_44_1049 ();
 sg13g2_fill_8 FILLER_0_44_1057 ();
 sg13g2_fill_8 FILLER_0_44_1065 ();
 sg13g2_fill_8 FILLER_0_44_1073 ();
 sg13g2_fill_8 FILLER_0_44_1081 ();
 sg13g2_fill_8 FILLER_0_44_1089 ();
 sg13g2_fill_8 FILLER_0_44_1097 ();
 sg13g2_fill_8 FILLER_0_44_1105 ();
 sg13g2_fill_8 FILLER_0_44_1113 ();
 sg13g2_fill_8 FILLER_0_44_1121 ();
 sg13g2_fill_8 FILLER_0_44_1129 ();
 sg13g2_fill_8 FILLER_0_44_1137 ();
 sg13g2_fill_8 FILLER_0_44_1145 ();
 sg13g2_fill_8 FILLER_0_44_1153 ();
 sg13g2_fill_8 FILLER_0_44_1161 ();
 sg13g2_fill_8 FILLER_0_44_1169 ();
 sg13g2_fill_8 FILLER_0_44_1177 ();
 sg13g2_fill_8 FILLER_0_44_1185 ();
 sg13g2_fill_8 FILLER_0_44_1193 ();
 sg13g2_fill_8 FILLER_0_44_1201 ();
 sg13g2_fill_8 FILLER_0_44_1209 ();
 sg13g2_fill_8 FILLER_0_44_1217 ();
 sg13g2_fill_2 FILLER_0_44_1225 ();
 sg13g2_fill_1 FILLER_0_44_1227 ();
 sg13g2_fill_4 FILLER_0_45_0 ();
 sg13g2_fill_2 FILLER_0_45_4 ();
 sg13g2_fill_1 FILLER_0_45_10 ();
 sg13g2_fill_1 FILLER_0_45_15 ();
 sg13g2_fill_1 FILLER_0_45_21 ();
 sg13g2_fill_1 FILLER_0_45_32 ();
 sg13g2_fill_4 FILLER_0_45_37 ();
 sg13g2_fill_2 FILLER_0_45_41 ();
 sg13g2_fill_8 FILLER_0_45_47 ();
 sg13g2_fill_4 FILLER_0_45_55 ();
 sg13g2_fill_4 FILLER_0_45_63 ();
 sg13g2_fill_8 FILLER_0_45_71 ();
 sg13g2_fill_4 FILLER_0_45_79 ();
 sg13g2_fill_2 FILLER_0_45_83 ();
 sg13g2_fill_2 FILLER_0_45_127 ();
 sg13g2_fill_1 FILLER_0_45_155 ();
 sg13g2_fill_1 FILLER_0_45_178 ();
 sg13g2_fill_8 FILLER_0_45_245 ();
 sg13g2_fill_2 FILLER_0_45_287 ();
 sg13g2_fill_8 FILLER_0_45_320 ();
 sg13g2_fill_4 FILLER_0_45_328 ();
 sg13g2_fill_1 FILLER_0_45_332 ();
 sg13g2_fill_4 FILLER_0_45_337 ();
 sg13g2_fill_1 FILLER_0_45_341 ();
 sg13g2_fill_1 FILLER_0_45_351 ();
 sg13g2_fill_4 FILLER_0_45_362 ();
 sg13g2_fill_4 FILLER_0_45_388 ();
 sg13g2_fill_8 FILLER_0_45_422 ();
 sg13g2_decap_8 FILLER_0_45_430 ();
 sg13g2_fill_1 FILLER_0_45_441 ();
 sg13g2_fill_1 FILLER_0_45_468 ();
 sg13g2_fill_1 FILLER_0_45_484 ();
 sg13g2_fill_1 FILLER_0_45_521 ();
 sg13g2_fill_8 FILLER_0_45_537 ();
 sg13g2_decap_8 FILLER_0_45_545 ();
 sg13g2_fill_8 FILLER_0_45_583 ();
 sg13g2_fill_2 FILLER_0_45_591 ();
 sg13g2_fill_1 FILLER_0_45_593 ();
 sg13g2_fill_8 FILLER_0_45_609 ();
 sg13g2_fill_8 FILLER_0_45_617 ();
 sg13g2_fill_8 FILLER_0_45_625 ();
 sg13g2_fill_8 FILLER_0_45_633 ();
 sg13g2_fill_8 FILLER_0_45_641 ();
 sg13g2_fill_8 FILLER_0_45_649 ();
 sg13g2_fill_8 FILLER_0_45_657 ();
 sg13g2_fill_8 FILLER_0_45_665 ();
 sg13g2_fill_8 FILLER_0_45_673 ();
 sg13g2_fill_8 FILLER_0_45_681 ();
 sg13g2_fill_8 FILLER_0_45_689 ();
 sg13g2_fill_8 FILLER_0_45_697 ();
 sg13g2_fill_1 FILLER_0_45_709 ();
 sg13g2_fill_8 FILLER_0_45_718 ();
 sg13g2_fill_8 FILLER_0_45_726 ();
 sg13g2_fill_4 FILLER_0_45_734 ();
 sg13g2_fill_1 FILLER_0_45_738 ();
 sg13g2_fill_8 FILLER_0_45_773 ();
 sg13g2_fill_1 FILLER_0_45_781 ();
 sg13g2_fill_4 FILLER_0_45_787 ();
 sg13g2_fill_1 FILLER_0_45_791 ();
 sg13g2_fill_4 FILLER_0_45_796 ();
 sg13g2_fill_8 FILLER_0_45_810 ();
 sg13g2_fill_2 FILLER_0_45_818 ();
 sg13g2_fill_1 FILLER_0_45_820 ();
 sg13g2_fill_4 FILLER_0_45_826 ();
 sg13g2_fill_1 FILLER_0_45_830 ();
 sg13g2_fill_4 FILLER_0_45_841 ();
 sg13g2_fill_1 FILLER_0_45_845 ();
 sg13g2_fill_4 FILLER_0_45_856 ();
 sg13g2_fill_4 FILLER_0_45_865 ();
 sg13g2_fill_1 FILLER_0_45_869 ();
 sg13g2_fill_8 FILLER_0_45_874 ();
 sg13g2_fill_8 FILLER_0_45_882 ();
 sg13g2_fill_8 FILLER_0_45_890 ();
 sg13g2_fill_8 FILLER_0_45_898 ();
 sg13g2_fill_8 FILLER_0_45_906 ();
 sg13g2_fill_8 FILLER_0_45_914 ();
 sg13g2_fill_8 FILLER_0_45_922 ();
 sg13g2_fill_8 FILLER_0_45_930 ();
 sg13g2_fill_8 FILLER_0_45_938 ();
 sg13g2_fill_8 FILLER_0_45_946 ();
 sg13g2_fill_8 FILLER_0_45_954 ();
 sg13g2_fill_8 FILLER_0_45_962 ();
 sg13g2_fill_8 FILLER_0_45_970 ();
 sg13g2_fill_8 FILLER_0_45_978 ();
 sg13g2_fill_8 FILLER_0_45_986 ();
 sg13g2_fill_8 FILLER_0_45_994 ();
 sg13g2_fill_8 FILLER_0_45_1002 ();
 sg13g2_fill_8 FILLER_0_45_1010 ();
 sg13g2_fill_8 FILLER_0_45_1018 ();
 sg13g2_fill_8 FILLER_0_45_1026 ();
 sg13g2_fill_8 FILLER_0_45_1034 ();
 sg13g2_fill_8 FILLER_0_45_1042 ();
 sg13g2_fill_8 FILLER_0_45_1050 ();
 sg13g2_fill_8 FILLER_0_45_1058 ();
 sg13g2_fill_8 FILLER_0_45_1066 ();
 sg13g2_fill_8 FILLER_0_45_1074 ();
 sg13g2_fill_8 FILLER_0_45_1082 ();
 sg13g2_fill_8 FILLER_0_45_1090 ();
 sg13g2_fill_8 FILLER_0_45_1098 ();
 sg13g2_fill_8 FILLER_0_45_1106 ();
 sg13g2_fill_8 FILLER_0_45_1114 ();
 sg13g2_fill_8 FILLER_0_45_1122 ();
 sg13g2_fill_8 FILLER_0_45_1130 ();
 sg13g2_fill_8 FILLER_0_45_1138 ();
 sg13g2_fill_8 FILLER_0_45_1146 ();
 sg13g2_fill_8 FILLER_0_45_1154 ();
 sg13g2_fill_8 FILLER_0_45_1162 ();
 sg13g2_fill_8 FILLER_0_45_1170 ();
 sg13g2_fill_8 FILLER_0_45_1178 ();
 sg13g2_fill_8 FILLER_0_45_1186 ();
 sg13g2_fill_8 FILLER_0_45_1194 ();
 sg13g2_fill_8 FILLER_0_45_1202 ();
 sg13g2_fill_8 FILLER_0_45_1210 ();
 sg13g2_fill_8 FILLER_0_45_1218 ();
 sg13g2_fill_2 FILLER_0_45_1226 ();
 sg13g2_fill_8 FILLER_0_46_0 ();
 sg13g2_fill_4 FILLER_0_46_8 ();
 sg13g2_fill_4 FILLER_0_46_17 ();
 sg13g2_fill_1 FILLER_0_46_21 ();
 sg13g2_fill_8 FILLER_0_46_32 ();
 sg13g2_fill_8 FILLER_0_46_40 ();
 sg13g2_fill_4 FILLER_0_46_48 ();
 sg13g2_fill_2 FILLER_0_46_52 ();
 sg13g2_fill_2 FILLER_0_46_58 ();
 sg13g2_fill_2 FILLER_0_46_65 ();
 sg13g2_fill_1 FILLER_0_46_67 ();
 sg13g2_decap_8 FILLER_0_46_72 ();
 sg13g2_fill_2 FILLER_0_46_119 ();
 sg13g2_fill_8 FILLER_0_46_126 ();
 sg13g2_fill_4 FILLER_0_46_134 ();
 sg13g2_fill_2 FILLER_0_46_138 ();
 sg13g2_fill_4 FILLER_0_46_150 ();
 sg13g2_fill_1 FILLER_0_46_154 ();
 sg13g2_fill_2 FILLER_0_46_175 ();
 sg13g2_fill_1 FILLER_0_46_177 ();
 sg13g2_fill_4 FILLER_0_46_192 ();
 sg13g2_fill_2 FILLER_0_46_206 ();
 sg13g2_fill_2 FILLER_0_46_218 ();
 sg13g2_fill_1 FILLER_0_46_220 ();
 sg13g2_fill_4 FILLER_0_46_278 ();
 sg13g2_fill_2 FILLER_0_46_386 ();
 sg13g2_fill_2 FILLER_0_46_398 ();
 sg13g2_fill_2 FILLER_0_46_405 ();
 sg13g2_fill_1 FILLER_0_46_407 ();
 sg13g2_fill_4 FILLER_0_46_434 ();
 sg13g2_fill_2 FILLER_0_46_438 ();
 sg13g2_fill_2 FILLER_0_46_481 ();
 sg13g2_fill_2 FILLER_0_46_513 ();
 sg13g2_fill_8 FILLER_0_46_546 ();
 sg13g2_fill_8 FILLER_0_46_554 ();
 sg13g2_fill_4 FILLER_0_46_562 ();
 sg13g2_fill_1 FILLER_0_46_570 ();
 sg13g2_fill_1 FILLER_0_46_597 ();
 sg13g2_fill_8 FILLER_0_46_624 ();
 sg13g2_fill_8 FILLER_0_46_632 ();
 sg13g2_fill_8 FILLER_0_46_640 ();
 sg13g2_fill_8 FILLER_0_46_648 ();
 sg13g2_fill_8 FILLER_0_46_656 ();
 sg13g2_fill_8 FILLER_0_46_664 ();
 sg13g2_fill_8 FILLER_0_46_672 ();
 sg13g2_fill_8 FILLER_0_46_680 ();
 sg13g2_fill_4 FILLER_0_46_688 ();
 sg13g2_fill_1 FILLER_0_46_692 ();
 sg13g2_fill_2 FILLER_0_46_734 ();
 sg13g2_fill_4 FILLER_0_46_812 ();
 sg13g2_fill_1 FILLER_0_46_816 ();
 sg13g2_fill_1 FILLER_0_46_843 ();
 sg13g2_fill_8 FILLER_0_46_880 ();
 sg13g2_fill_8 FILLER_0_46_888 ();
 sg13g2_fill_8 FILLER_0_46_896 ();
 sg13g2_fill_8 FILLER_0_46_904 ();
 sg13g2_fill_8 FILLER_0_46_912 ();
 sg13g2_fill_8 FILLER_0_46_920 ();
 sg13g2_fill_8 FILLER_0_46_928 ();
 sg13g2_fill_8 FILLER_0_46_936 ();
 sg13g2_fill_8 FILLER_0_46_944 ();
 sg13g2_fill_8 FILLER_0_46_952 ();
 sg13g2_fill_8 FILLER_0_46_960 ();
 sg13g2_fill_8 FILLER_0_46_968 ();
 sg13g2_fill_8 FILLER_0_46_976 ();
 sg13g2_fill_8 FILLER_0_46_984 ();
 sg13g2_fill_8 FILLER_0_46_992 ();
 sg13g2_fill_8 FILLER_0_46_1000 ();
 sg13g2_fill_8 FILLER_0_46_1008 ();
 sg13g2_fill_8 FILLER_0_46_1016 ();
 sg13g2_fill_8 FILLER_0_46_1024 ();
 sg13g2_fill_8 FILLER_0_46_1032 ();
 sg13g2_fill_8 FILLER_0_46_1040 ();
 sg13g2_fill_8 FILLER_0_46_1048 ();
 sg13g2_fill_8 FILLER_0_46_1056 ();
 sg13g2_fill_8 FILLER_0_46_1064 ();
 sg13g2_fill_8 FILLER_0_46_1072 ();
 sg13g2_fill_8 FILLER_0_46_1080 ();
 sg13g2_fill_8 FILLER_0_46_1088 ();
 sg13g2_fill_8 FILLER_0_46_1096 ();
 sg13g2_fill_8 FILLER_0_46_1104 ();
 sg13g2_fill_8 FILLER_0_46_1112 ();
 sg13g2_fill_8 FILLER_0_46_1120 ();
 sg13g2_fill_8 FILLER_0_46_1128 ();
 sg13g2_fill_8 FILLER_0_46_1136 ();
 sg13g2_fill_8 FILLER_0_46_1144 ();
 sg13g2_fill_8 FILLER_0_46_1152 ();
 sg13g2_fill_8 FILLER_0_46_1160 ();
 sg13g2_fill_8 FILLER_0_46_1168 ();
 sg13g2_fill_8 FILLER_0_46_1176 ();
 sg13g2_fill_8 FILLER_0_46_1184 ();
 sg13g2_fill_8 FILLER_0_46_1192 ();
 sg13g2_fill_8 FILLER_0_46_1200 ();
 sg13g2_fill_8 FILLER_0_46_1208 ();
 sg13g2_fill_8 FILLER_0_46_1216 ();
 sg13g2_fill_4 FILLER_0_46_1224 ();
 sg13g2_fill_1 FILLER_0_47_0 ();
 sg13g2_fill_2 FILLER_0_47_27 ();
 sg13g2_fill_2 FILLER_0_47_115 ();
 sg13g2_fill_8 FILLER_0_47_127 ();
 sg13g2_fill_1 FILLER_0_47_135 ();
 sg13g2_fill_4 FILLER_0_47_177 ();
 sg13g2_fill_1 FILLER_0_47_181 ();
 sg13g2_fill_8 FILLER_0_47_186 ();
 sg13g2_fill_8 FILLER_0_47_194 ();
 sg13g2_fill_4 FILLER_0_47_202 ();
 sg13g2_fill_2 FILLER_0_47_206 ();
 sg13g2_fill_2 FILLER_0_47_223 ();
 sg13g2_fill_1 FILLER_0_47_225 ();
 sg13g2_fill_2 FILLER_0_47_230 ();
 sg13g2_fill_4 FILLER_0_47_236 ();
 sg13g2_fill_2 FILLER_0_47_262 ();
 sg13g2_fill_1 FILLER_0_47_264 ();
 sg13g2_fill_1 FILLER_0_47_318 ();
 sg13g2_fill_2 FILLER_0_47_323 ();
 sg13g2_fill_8 FILLER_0_47_335 ();
 sg13g2_fill_2 FILLER_0_47_343 ();
 sg13g2_fill_1 FILLER_0_47_345 ();
 sg13g2_fill_8 FILLER_0_47_350 ();
 sg13g2_fill_2 FILLER_0_47_358 ();
 sg13g2_fill_2 FILLER_0_47_374 ();
 sg13g2_fill_1 FILLER_0_47_401 ();
 sg13g2_fill_8 FILLER_0_47_406 ();
 sg13g2_fill_2 FILLER_0_47_414 ();
 sg13g2_fill_8 FILLER_0_47_420 ();
 sg13g2_fill_8 FILLER_0_47_428 ();
 sg13g2_fill_2 FILLER_0_47_436 ();
 sg13g2_fill_1 FILLER_0_47_438 ();
 sg13g2_fill_1 FILLER_0_47_456 ();
 sg13g2_fill_2 FILLER_0_47_462 ();
 sg13g2_fill_8 FILLER_0_47_483 ();
 sg13g2_fill_1 FILLER_0_47_491 ();
 sg13g2_fill_1 FILLER_0_47_500 ();
 sg13g2_fill_8 FILLER_0_47_509 ();
 sg13g2_fill_2 FILLER_0_47_517 ();
 sg13g2_fill_1 FILLER_0_47_529 ();
 sg13g2_fill_4 FILLER_0_47_542 ();
 sg13g2_fill_2 FILLER_0_47_546 ();
 sg13g2_fill_4 FILLER_0_47_563 ();
 sg13g2_fill_1 FILLER_0_47_567 ();
 sg13g2_fill_1 FILLER_0_47_573 ();
 sg13g2_fill_4 FILLER_0_47_588 ();
 sg13g2_fill_2 FILLER_0_47_592 ();
 sg13g2_fill_8 FILLER_0_47_630 ();
 sg13g2_fill_8 FILLER_0_47_638 ();
 sg13g2_fill_8 FILLER_0_47_646 ();
 sg13g2_fill_8 FILLER_0_47_654 ();
 sg13g2_fill_8 FILLER_0_47_662 ();
 sg13g2_fill_8 FILLER_0_47_670 ();
 sg13g2_fill_8 FILLER_0_47_678 ();
 sg13g2_fill_4 FILLER_0_47_686 ();
 sg13g2_fill_2 FILLER_0_47_690 ();
 sg13g2_fill_1 FILLER_0_47_733 ();
 sg13g2_fill_2 FILLER_0_47_760 ();
 sg13g2_fill_2 FILLER_0_47_772 ();
 sg13g2_fill_1 FILLER_0_47_774 ();
 sg13g2_fill_2 FILLER_0_47_779 ();
 sg13g2_fill_1 FILLER_0_47_781 ();
 sg13g2_fill_1 FILLER_0_47_848 ();
 sg13g2_fill_8 FILLER_0_47_880 ();
 sg13g2_fill_8 FILLER_0_47_888 ();
 sg13g2_fill_8 FILLER_0_47_896 ();
 sg13g2_fill_8 FILLER_0_47_904 ();
 sg13g2_fill_8 FILLER_0_47_912 ();
 sg13g2_fill_8 FILLER_0_47_920 ();
 sg13g2_fill_8 FILLER_0_47_928 ();
 sg13g2_fill_8 FILLER_0_47_936 ();
 sg13g2_fill_8 FILLER_0_47_944 ();
 sg13g2_fill_8 FILLER_0_47_952 ();
 sg13g2_fill_8 FILLER_0_47_960 ();
 sg13g2_fill_8 FILLER_0_47_968 ();
 sg13g2_fill_8 FILLER_0_47_976 ();
 sg13g2_fill_8 FILLER_0_47_984 ();
 sg13g2_fill_8 FILLER_0_47_992 ();
 sg13g2_fill_8 FILLER_0_47_1000 ();
 sg13g2_fill_8 FILLER_0_47_1008 ();
 sg13g2_fill_8 FILLER_0_47_1016 ();
 sg13g2_fill_8 FILLER_0_47_1024 ();
 sg13g2_fill_8 FILLER_0_47_1032 ();
 sg13g2_fill_8 FILLER_0_47_1040 ();
 sg13g2_fill_8 FILLER_0_47_1048 ();
 sg13g2_fill_8 FILLER_0_47_1056 ();
 sg13g2_fill_8 FILLER_0_47_1064 ();
 sg13g2_fill_8 FILLER_0_47_1072 ();
 sg13g2_fill_8 FILLER_0_47_1080 ();
 sg13g2_fill_8 FILLER_0_47_1088 ();
 sg13g2_fill_8 FILLER_0_47_1096 ();
 sg13g2_fill_8 FILLER_0_47_1104 ();
 sg13g2_fill_8 FILLER_0_47_1112 ();
 sg13g2_fill_8 FILLER_0_47_1120 ();
 sg13g2_fill_8 FILLER_0_47_1128 ();
 sg13g2_fill_8 FILLER_0_47_1136 ();
 sg13g2_fill_8 FILLER_0_47_1144 ();
 sg13g2_fill_8 FILLER_0_47_1152 ();
 sg13g2_fill_8 FILLER_0_47_1160 ();
 sg13g2_fill_8 FILLER_0_47_1168 ();
 sg13g2_fill_8 FILLER_0_47_1176 ();
 sg13g2_fill_8 FILLER_0_47_1184 ();
 sg13g2_fill_8 FILLER_0_47_1192 ();
 sg13g2_fill_8 FILLER_0_47_1200 ();
 sg13g2_fill_8 FILLER_0_47_1208 ();
 sg13g2_fill_8 FILLER_0_47_1216 ();
 sg13g2_fill_4 FILLER_0_47_1224 ();
 sg13g2_decap_8 FILLER_0_48_0 ();
 sg13g2_fill_8 FILLER_0_48_11 ();
 sg13g2_fill_2 FILLER_0_48_19 ();
 sg13g2_fill_4 FILLER_0_48_47 ();
 sg13g2_decap_8 FILLER_0_48_81 ();
 sg13g2_fill_1 FILLER_0_48_123 ();
 sg13g2_fill_2 FILLER_0_48_129 ();
 sg13g2_fill_2 FILLER_0_48_157 ();
 sg13g2_fill_2 FILLER_0_48_185 ();
 sg13g2_fill_8 FILLER_0_48_197 ();
 sg13g2_fill_4 FILLER_0_48_205 ();
 sg13g2_fill_4 FILLER_0_48_224 ();
 sg13g2_fill_2 FILLER_0_48_228 ();
 sg13g2_fill_8 FILLER_0_48_234 ();
 sg13g2_fill_4 FILLER_0_48_242 ();
 sg13g2_fill_2 FILLER_0_48_250 ();
 sg13g2_fill_4 FILLER_0_48_278 ();
 sg13g2_fill_8 FILLER_0_48_286 ();
 sg13g2_fill_2 FILLER_0_48_294 ();
 sg13g2_fill_1 FILLER_0_48_296 ();
 sg13g2_fill_8 FILLER_0_48_301 ();
 sg13g2_fill_1 FILLER_0_48_309 ();
 sg13g2_fill_2 FILLER_0_48_330 ();
 sg13g2_fill_1 FILLER_0_48_332 ();
 sg13g2_fill_1 FILLER_0_48_338 ();
 sg13g2_fill_8 FILLER_0_48_395 ();
 sg13g2_fill_8 FILLER_0_48_403 ();
 sg13g2_fill_8 FILLER_0_48_411 ();
 sg13g2_fill_2 FILLER_0_48_419 ();
 sg13g2_fill_1 FILLER_0_48_421 ();
 sg13g2_fill_4 FILLER_0_48_432 ();
 sg13g2_fill_8 FILLER_0_48_487 ();
 sg13g2_fill_8 FILLER_0_48_495 ();
 sg13g2_fill_1 FILLER_0_48_548 ();
 sg13g2_fill_4 FILLER_0_48_575 ();
 sg13g2_fill_2 FILLER_0_48_579 ();
 sg13g2_fill_2 FILLER_0_48_599 ();
 sg13g2_fill_8 FILLER_0_48_619 ();
 sg13g2_fill_8 FILLER_0_48_627 ();
 sg13g2_fill_8 FILLER_0_48_635 ();
 sg13g2_fill_8 FILLER_0_48_643 ();
 sg13g2_fill_8 FILLER_0_48_651 ();
 sg13g2_fill_8 FILLER_0_48_659 ();
 sg13g2_fill_8 FILLER_0_48_667 ();
 sg13g2_fill_8 FILLER_0_48_675 ();
 sg13g2_fill_8 FILLER_0_48_683 ();
 sg13g2_fill_8 FILLER_0_48_691 ();
 sg13g2_fill_1 FILLER_0_48_703 ();
 sg13g2_fill_2 FILLER_0_48_708 ();
 sg13g2_fill_8 FILLER_0_48_766 ();
 sg13g2_fill_2 FILLER_0_48_774 ();
 sg13g2_fill_4 FILLER_0_48_800 ();
 sg13g2_fill_4 FILLER_0_48_812 ();
 sg13g2_fill_2 FILLER_0_48_816 ();
 sg13g2_fill_4 FILLER_0_48_827 ();
 sg13g2_fill_2 FILLER_0_48_835 ();
 sg13g2_fill_1 FILLER_0_48_837 ();
 sg13g2_fill_8 FILLER_0_48_848 ();
 sg13g2_fill_4 FILLER_0_48_856 ();
 sg13g2_fill_8 FILLER_0_48_872 ();
 sg13g2_fill_8 FILLER_0_48_880 ();
 sg13g2_fill_8 FILLER_0_48_888 ();
 sg13g2_fill_8 FILLER_0_48_896 ();
 sg13g2_fill_8 FILLER_0_48_904 ();
 sg13g2_fill_8 FILLER_0_48_912 ();
 sg13g2_fill_8 FILLER_0_48_920 ();
 sg13g2_fill_8 FILLER_0_48_928 ();
 sg13g2_fill_8 FILLER_0_48_936 ();
 sg13g2_fill_8 FILLER_0_48_944 ();
 sg13g2_fill_8 FILLER_0_48_952 ();
 sg13g2_fill_8 FILLER_0_48_960 ();
 sg13g2_fill_8 FILLER_0_48_968 ();
 sg13g2_fill_8 FILLER_0_48_976 ();
 sg13g2_fill_8 FILLER_0_48_984 ();
 sg13g2_fill_8 FILLER_0_48_992 ();
 sg13g2_fill_8 FILLER_0_48_1000 ();
 sg13g2_fill_8 FILLER_0_48_1008 ();
 sg13g2_fill_8 FILLER_0_48_1016 ();
 sg13g2_fill_8 FILLER_0_48_1024 ();
 sg13g2_fill_8 FILLER_0_48_1032 ();
 sg13g2_fill_8 FILLER_0_48_1040 ();
 sg13g2_fill_8 FILLER_0_48_1048 ();
 sg13g2_fill_8 FILLER_0_48_1056 ();
 sg13g2_fill_8 FILLER_0_48_1064 ();
 sg13g2_fill_8 FILLER_0_48_1072 ();
 sg13g2_fill_8 FILLER_0_48_1080 ();
 sg13g2_fill_8 FILLER_0_48_1088 ();
 sg13g2_fill_8 FILLER_0_48_1096 ();
 sg13g2_fill_8 FILLER_0_48_1104 ();
 sg13g2_fill_8 FILLER_0_48_1112 ();
 sg13g2_fill_8 FILLER_0_48_1120 ();
 sg13g2_fill_8 FILLER_0_48_1128 ();
 sg13g2_fill_8 FILLER_0_48_1136 ();
 sg13g2_fill_8 FILLER_0_48_1144 ();
 sg13g2_fill_8 FILLER_0_48_1152 ();
 sg13g2_fill_8 FILLER_0_48_1160 ();
 sg13g2_fill_8 FILLER_0_48_1168 ();
 sg13g2_fill_8 FILLER_0_48_1176 ();
 sg13g2_fill_8 FILLER_0_48_1184 ();
 sg13g2_fill_8 FILLER_0_48_1192 ();
 sg13g2_fill_8 FILLER_0_48_1200 ();
 sg13g2_fill_8 FILLER_0_48_1208 ();
 sg13g2_fill_8 FILLER_0_48_1216 ();
 sg13g2_fill_4 FILLER_0_48_1224 ();
 sg13g2_fill_8 FILLER_0_49_0 ();
 sg13g2_fill_8 FILLER_0_49_8 ();
 sg13g2_fill_1 FILLER_0_49_16 ();
 sg13g2_fill_2 FILLER_0_49_31 ();
 sg13g2_fill_8 FILLER_0_49_41 ();
 sg13g2_fill_1 FILLER_0_49_49 ();
 sg13g2_fill_2 FILLER_0_49_55 ();
 sg13g2_fill_1 FILLER_0_49_71 ();
 sg13g2_fill_8 FILLER_0_49_82 ();
 sg13g2_fill_8 FILLER_0_49_90 ();
 sg13g2_fill_2 FILLER_0_49_98 ();
 sg13g2_fill_1 FILLER_0_49_100 ();
 sg13g2_fill_2 FILLER_0_49_115 ();
 sg13g2_fill_1 FILLER_0_49_117 ();
 sg13g2_fill_2 FILLER_0_49_158 ();
 sg13g2_fill_2 FILLER_0_49_201 ();
 sg13g2_fill_2 FILLER_0_49_213 ();
 sg13g2_fill_2 FILLER_0_49_220 ();
 sg13g2_fill_2 FILLER_0_49_248 ();
 sg13g2_fill_4 FILLER_0_49_276 ();
 sg13g2_fill_2 FILLER_0_49_285 ();
 sg13g2_fill_8 FILLER_0_49_306 ();
 sg13g2_fill_2 FILLER_0_49_314 ();
 sg13g2_fill_8 FILLER_0_49_332 ();
 sg13g2_fill_4 FILLER_0_49_344 ();
 sg13g2_fill_8 FILLER_0_49_393 ();
 sg13g2_fill_2 FILLER_0_49_401 ();
 sg13g2_fill_8 FILLER_0_49_438 ();
 sg13g2_fill_8 FILLER_0_49_446 ();
 sg13g2_fill_2 FILLER_0_49_510 ();
 sg13g2_fill_1 FILLER_0_49_512 ();
 sg13g2_fill_4 FILLER_0_49_518 ();
 sg13g2_fill_1 FILLER_0_49_522 ();
 sg13g2_fill_4 FILLER_0_49_532 ();
 sg13g2_fill_1 FILLER_0_49_536 ();
 sg13g2_fill_8 FILLER_0_49_541 ();
 sg13g2_fill_8 FILLER_0_49_549 ();
 sg13g2_fill_1 FILLER_0_49_557 ();
 sg13g2_fill_1 FILLER_0_49_562 ();
 sg13g2_fill_8 FILLER_0_49_567 ();
 sg13g2_fill_8 FILLER_0_49_575 ();
 sg13g2_fill_1 FILLER_0_49_591 ();
 sg13g2_fill_8 FILLER_0_49_618 ();
 sg13g2_fill_8 FILLER_0_49_626 ();
 sg13g2_fill_8 FILLER_0_49_634 ();
 sg13g2_fill_8 FILLER_0_49_642 ();
 sg13g2_fill_4 FILLER_0_49_650 ();
 sg13g2_fill_2 FILLER_0_49_654 ();
 sg13g2_fill_8 FILLER_0_49_682 ();
 sg13g2_fill_8 FILLER_0_49_690 ();
 sg13g2_fill_4 FILLER_0_49_698 ();
 sg13g2_fill_1 FILLER_0_49_702 ();
 sg13g2_fill_1 FILLER_0_49_716 ();
 sg13g2_fill_2 FILLER_0_49_735 ();
 sg13g2_fill_1 FILLER_0_49_737 ();
 sg13g2_fill_2 FILLER_0_49_743 ();
 sg13g2_fill_8 FILLER_0_49_759 ();
 sg13g2_fill_2 FILLER_0_49_767 ();
 sg13g2_fill_1 FILLER_0_49_769 ();
 sg13g2_fill_2 FILLER_0_49_778 ();
 sg13g2_fill_8 FILLER_0_49_785 ();
 sg13g2_fill_4 FILLER_0_49_793 ();
 sg13g2_fill_8 FILLER_0_49_801 ();
 sg13g2_fill_4 FILLER_0_49_809 ();
 sg13g2_fill_2 FILLER_0_49_822 ();
 sg13g2_fill_1 FILLER_0_49_855 ();
 sg13g2_fill_2 FILLER_0_49_861 ();
 sg13g2_fill_2 FILLER_0_49_867 ();
 sg13g2_fill_8 FILLER_0_49_873 ();
 sg13g2_fill_8 FILLER_0_49_886 ();
 sg13g2_fill_8 FILLER_0_49_894 ();
 sg13g2_fill_8 FILLER_0_49_902 ();
 sg13g2_fill_8 FILLER_0_49_910 ();
 sg13g2_fill_8 FILLER_0_49_918 ();
 sg13g2_fill_8 FILLER_0_49_926 ();
 sg13g2_fill_8 FILLER_0_49_934 ();
 sg13g2_fill_8 FILLER_0_49_942 ();
 sg13g2_fill_8 FILLER_0_49_950 ();
 sg13g2_fill_8 FILLER_0_49_958 ();
 sg13g2_fill_8 FILLER_0_49_966 ();
 sg13g2_fill_8 FILLER_0_49_974 ();
 sg13g2_fill_8 FILLER_0_49_982 ();
 sg13g2_fill_8 FILLER_0_49_990 ();
 sg13g2_fill_8 FILLER_0_49_998 ();
 sg13g2_fill_8 FILLER_0_49_1006 ();
 sg13g2_fill_8 FILLER_0_49_1014 ();
 sg13g2_fill_8 FILLER_0_49_1022 ();
 sg13g2_fill_8 FILLER_0_49_1030 ();
 sg13g2_fill_8 FILLER_0_49_1038 ();
 sg13g2_fill_8 FILLER_0_49_1046 ();
 sg13g2_fill_8 FILLER_0_49_1054 ();
 sg13g2_fill_8 FILLER_0_49_1062 ();
 sg13g2_fill_8 FILLER_0_49_1070 ();
 sg13g2_fill_8 FILLER_0_49_1078 ();
 sg13g2_fill_8 FILLER_0_49_1086 ();
 sg13g2_fill_8 FILLER_0_49_1094 ();
 sg13g2_fill_8 FILLER_0_49_1102 ();
 sg13g2_fill_8 FILLER_0_49_1110 ();
 sg13g2_fill_8 FILLER_0_49_1118 ();
 sg13g2_fill_8 FILLER_0_49_1126 ();
 sg13g2_fill_8 FILLER_0_49_1134 ();
 sg13g2_fill_8 FILLER_0_49_1142 ();
 sg13g2_fill_8 FILLER_0_49_1150 ();
 sg13g2_fill_8 FILLER_0_49_1158 ();
 sg13g2_fill_8 FILLER_0_49_1166 ();
 sg13g2_fill_8 FILLER_0_49_1174 ();
 sg13g2_fill_8 FILLER_0_49_1182 ();
 sg13g2_fill_8 FILLER_0_49_1190 ();
 sg13g2_fill_8 FILLER_0_49_1198 ();
 sg13g2_fill_8 FILLER_0_49_1206 ();
 sg13g2_fill_8 FILLER_0_49_1214 ();
 sg13g2_fill_4 FILLER_0_49_1222 ();
 sg13g2_fill_2 FILLER_0_49_1226 ();
 sg13g2_fill_1 FILLER_0_50_0 ();
 sg13g2_fill_8 FILLER_0_50_32 ();
 sg13g2_fill_2 FILLER_0_50_40 ();
 sg13g2_fill_8 FILLER_0_50_81 ();
 sg13g2_fill_8 FILLER_0_50_89 ();
 sg13g2_fill_4 FILLER_0_50_97 ();
 sg13g2_fill_1 FILLER_0_50_101 ();
 sg13g2_fill_1 FILLER_0_50_128 ();
 sg13g2_fill_4 FILLER_0_50_133 ();
 sg13g2_fill_1 FILLER_0_50_137 ();
 sg13g2_fill_8 FILLER_0_50_142 ();
 sg13g2_fill_2 FILLER_0_50_150 ();
 sg13g2_fill_8 FILLER_0_50_157 ();
 sg13g2_fill_2 FILLER_0_50_165 ();
 sg13g2_fill_1 FILLER_0_50_176 ();
 sg13g2_fill_1 FILLER_0_50_182 ();
 sg13g2_fill_1 FILLER_0_50_219 ();
 sg13g2_fill_8 FILLER_0_50_246 ();
 sg13g2_fill_2 FILLER_0_50_254 ();
 sg13g2_fill_1 FILLER_0_50_256 ();
 sg13g2_fill_2 FILLER_0_50_261 ();
 sg13g2_fill_2 FILLER_0_50_319 ();
 sg13g2_fill_2 FILLER_0_50_347 ();
 sg13g2_fill_1 FILLER_0_50_349 ();
 sg13g2_fill_2 FILLER_0_50_368 ();
 sg13g2_fill_8 FILLER_0_50_440 ();
 sg13g2_fill_4 FILLER_0_50_448 ();
 sg13g2_fill_8 FILLER_0_50_456 ();
 sg13g2_fill_2 FILLER_0_50_464 ();
 sg13g2_fill_2 FILLER_0_50_480 ();
 sg13g2_fill_2 FILLER_0_50_522 ();
 sg13g2_fill_1 FILLER_0_50_558 ();
 sg13g2_fill_2 FILLER_0_50_564 ();
 sg13g2_fill_1 FILLER_0_50_566 ();
 sg13g2_fill_4 FILLER_0_50_577 ();
 sg13g2_fill_1 FILLER_0_50_622 ();
 sg13g2_fill_1 FILLER_0_50_685 ();
 sg13g2_fill_8 FILLER_0_50_690 ();
 sg13g2_fill_2 FILLER_0_50_698 ();
 sg13g2_fill_4 FILLER_0_50_731 ();
 sg13g2_fill_2 FILLER_0_50_735 ();
 sg13g2_fill_4 FILLER_0_50_768 ();
 sg13g2_fill_1 FILLER_0_50_808 ();
 sg13g2_fill_2 FILLER_0_50_814 ();
 sg13g2_fill_1 FILLER_0_50_914 ();
 sg13g2_fill_8 FILLER_0_50_919 ();
 sg13g2_fill_8 FILLER_0_50_927 ();
 sg13g2_fill_8 FILLER_0_50_935 ();
 sg13g2_fill_8 FILLER_0_50_943 ();
 sg13g2_fill_8 FILLER_0_50_951 ();
 sg13g2_fill_8 FILLER_0_50_959 ();
 sg13g2_fill_8 FILLER_0_50_967 ();
 sg13g2_fill_8 FILLER_0_50_975 ();
 sg13g2_fill_8 FILLER_0_50_983 ();
 sg13g2_fill_8 FILLER_0_50_991 ();
 sg13g2_fill_8 FILLER_0_50_999 ();
 sg13g2_fill_8 FILLER_0_50_1007 ();
 sg13g2_fill_8 FILLER_0_50_1015 ();
 sg13g2_fill_8 FILLER_0_50_1023 ();
 sg13g2_fill_8 FILLER_0_50_1031 ();
 sg13g2_fill_8 FILLER_0_50_1039 ();
 sg13g2_fill_8 FILLER_0_50_1047 ();
 sg13g2_fill_8 FILLER_0_50_1055 ();
 sg13g2_fill_8 FILLER_0_50_1063 ();
 sg13g2_fill_8 FILLER_0_50_1071 ();
 sg13g2_fill_8 FILLER_0_50_1079 ();
 sg13g2_fill_8 FILLER_0_50_1087 ();
 sg13g2_fill_8 FILLER_0_50_1095 ();
 sg13g2_fill_8 FILLER_0_50_1103 ();
 sg13g2_fill_8 FILLER_0_50_1111 ();
 sg13g2_fill_8 FILLER_0_50_1119 ();
 sg13g2_fill_8 FILLER_0_50_1127 ();
 sg13g2_fill_8 FILLER_0_50_1135 ();
 sg13g2_fill_8 FILLER_0_50_1143 ();
 sg13g2_fill_8 FILLER_0_50_1151 ();
 sg13g2_fill_8 FILLER_0_50_1159 ();
 sg13g2_fill_8 FILLER_0_50_1167 ();
 sg13g2_fill_8 FILLER_0_50_1175 ();
 sg13g2_fill_8 FILLER_0_50_1183 ();
 sg13g2_fill_8 FILLER_0_50_1191 ();
 sg13g2_fill_8 FILLER_0_50_1199 ();
 sg13g2_fill_8 FILLER_0_50_1207 ();
 sg13g2_fill_8 FILLER_0_50_1215 ();
 sg13g2_fill_4 FILLER_0_50_1223 ();
 sg13g2_fill_1 FILLER_0_50_1227 ();
 sg13g2_fill_1 FILLER_0_51_0 ();
 sg13g2_fill_8 FILLER_0_51_63 ();
 sg13g2_fill_8 FILLER_0_51_71 ();
 sg13g2_fill_1 FILLER_0_51_79 ();
 sg13g2_fill_8 FILLER_0_51_84 ();
 sg13g2_fill_8 FILLER_0_51_92 ();
 sg13g2_fill_1 FILLER_0_51_100 ();
 sg13g2_fill_4 FILLER_0_51_111 ();
 sg13g2_fill_2 FILLER_0_51_115 ();
 sg13g2_fill_2 FILLER_0_51_121 ();
 sg13g2_fill_1 FILLER_0_51_123 ();
 sg13g2_fill_2 FILLER_0_51_132 ();
 sg13g2_fill_1 FILLER_0_51_134 ();
 sg13g2_fill_8 FILLER_0_51_161 ();
 sg13g2_fill_8 FILLER_0_51_169 ();
 sg13g2_fill_1 FILLER_0_51_177 ();
 sg13g2_fill_4 FILLER_0_51_186 ();
 sg13g2_fill_2 FILLER_0_51_190 ();
 sg13g2_fill_2 FILLER_0_51_196 ();
 sg13g2_fill_1 FILLER_0_51_198 ();
 sg13g2_fill_8 FILLER_0_51_239 ();
 sg13g2_fill_4 FILLER_0_51_247 ();
 sg13g2_fill_2 FILLER_0_51_251 ();
 sg13g2_fill_4 FILLER_0_51_258 ();
 sg13g2_fill_1 FILLER_0_51_262 ();
 sg13g2_fill_1 FILLER_0_51_293 ();
 sg13g2_fill_4 FILLER_0_51_320 ();
 sg13g2_fill_1 FILLER_0_51_324 ();
 sg13g2_fill_2 FILLER_0_51_361 ();
 sg13g2_fill_2 FILLER_0_51_373 ();
 sg13g2_fill_1 FILLER_0_51_375 ();
 sg13g2_fill_2 FILLER_0_51_402 ();
 sg13g2_decap_8 FILLER_0_51_471 ();
 sg13g2_fill_8 FILLER_0_51_493 ();
 sg13g2_fill_4 FILLER_0_51_501 ();
 sg13g2_fill_2 FILLER_0_51_509 ();
 sg13g2_fill_4 FILLER_0_51_515 ();
 sg13g2_fill_1 FILLER_0_51_519 ();
 sg13g2_fill_1 FILLER_0_51_530 ();
 sg13g2_fill_1 FILLER_0_51_535 ();
 sg13g2_fill_2 FILLER_0_51_546 ();
 sg13g2_fill_2 FILLER_0_51_552 ();
 sg13g2_fill_1 FILLER_0_51_554 ();
 sg13g2_fill_2 FILLER_0_51_581 ();
 sg13g2_fill_4 FILLER_0_51_619 ();
 sg13g2_fill_1 FILLER_0_51_623 ();
 sg13g2_fill_1 FILLER_0_51_655 ();
 sg13g2_fill_2 FILLER_0_51_706 ();
 sg13g2_fill_1 FILLER_0_51_708 ();
 sg13g2_fill_8 FILLER_0_51_717 ();
 sg13g2_fill_2 FILLER_0_51_725 ();
 sg13g2_fill_1 FILLER_0_51_766 ();
 sg13g2_fill_1 FILLER_0_51_797 ();
 sg13g2_fill_1 FILLER_0_51_802 ();
 sg13g2_fill_1 FILLER_0_51_855 ();
 sg13g2_fill_8 FILLER_0_51_918 ();
 sg13g2_fill_8 FILLER_0_51_926 ();
 sg13g2_fill_8 FILLER_0_51_934 ();
 sg13g2_fill_8 FILLER_0_51_942 ();
 sg13g2_fill_8 FILLER_0_51_950 ();
 sg13g2_fill_8 FILLER_0_51_958 ();
 sg13g2_fill_8 FILLER_0_51_966 ();
 sg13g2_fill_8 FILLER_0_51_974 ();
 sg13g2_fill_8 FILLER_0_51_982 ();
 sg13g2_fill_8 FILLER_0_51_990 ();
 sg13g2_fill_8 FILLER_0_51_998 ();
 sg13g2_fill_8 FILLER_0_51_1006 ();
 sg13g2_fill_8 FILLER_0_51_1014 ();
 sg13g2_fill_8 FILLER_0_51_1022 ();
 sg13g2_fill_8 FILLER_0_51_1030 ();
 sg13g2_fill_8 FILLER_0_51_1038 ();
 sg13g2_fill_8 FILLER_0_51_1046 ();
 sg13g2_fill_8 FILLER_0_51_1054 ();
 sg13g2_fill_8 FILLER_0_51_1062 ();
 sg13g2_fill_8 FILLER_0_51_1070 ();
 sg13g2_fill_8 FILLER_0_51_1078 ();
 sg13g2_fill_8 FILLER_0_51_1086 ();
 sg13g2_fill_8 FILLER_0_51_1094 ();
 sg13g2_fill_8 FILLER_0_51_1102 ();
 sg13g2_fill_8 FILLER_0_51_1110 ();
 sg13g2_fill_8 FILLER_0_51_1118 ();
 sg13g2_fill_8 FILLER_0_51_1126 ();
 sg13g2_fill_8 FILLER_0_51_1134 ();
 sg13g2_fill_8 FILLER_0_51_1142 ();
 sg13g2_fill_8 FILLER_0_51_1150 ();
 sg13g2_fill_8 FILLER_0_51_1158 ();
 sg13g2_fill_8 FILLER_0_51_1166 ();
 sg13g2_fill_8 FILLER_0_51_1174 ();
 sg13g2_fill_8 FILLER_0_51_1182 ();
 sg13g2_fill_8 FILLER_0_51_1190 ();
 sg13g2_fill_8 FILLER_0_51_1198 ();
 sg13g2_fill_8 FILLER_0_51_1206 ();
 sg13g2_fill_8 FILLER_0_51_1214 ();
 sg13g2_fill_4 FILLER_0_51_1222 ();
 sg13g2_fill_2 FILLER_0_51_1226 ();
 sg13g2_decap_8 FILLER_0_52_0 ();
 sg13g2_fill_1 FILLER_0_52_20 ();
 sg13g2_fill_1 FILLER_0_52_73 ();
 sg13g2_fill_1 FILLER_0_52_100 ();
 sg13g2_fill_1 FILLER_0_52_106 ();
 sg13g2_fill_2 FILLER_0_52_133 ();
 sg13g2_fill_1 FILLER_0_52_140 ();
 sg13g2_fill_2 FILLER_0_52_167 ();
 sg13g2_fill_8 FILLER_0_52_195 ();
 sg13g2_fill_8 FILLER_0_52_203 ();
 sg13g2_fill_8 FILLER_0_52_215 ();
 sg13g2_fill_1 FILLER_0_52_223 ();
 sg13g2_fill_4 FILLER_0_52_260 ();
 sg13g2_fill_1 FILLER_0_52_264 ();
 sg13g2_fill_8 FILLER_0_52_275 ();
 sg13g2_decap_8 FILLER_0_52_283 ();
 sg13g2_fill_2 FILLER_0_52_295 ();
 sg13g2_fill_1 FILLER_0_52_297 ();
 sg13g2_fill_8 FILLER_0_52_306 ();
 sg13g2_fill_8 FILLER_0_52_314 ();
 sg13g2_fill_1 FILLER_0_52_336 ();
 sg13g2_fill_1 FILLER_0_52_389 ();
 sg13g2_fill_4 FILLER_0_52_406 ();
 sg13g2_fill_4 FILLER_0_52_414 ();
 sg13g2_fill_1 FILLER_0_52_418 ();
 sg13g2_fill_2 FILLER_0_52_442 ();
 sg13g2_fill_1 FILLER_0_52_444 ();
 sg13g2_fill_1 FILLER_0_52_449 ();
 sg13g2_fill_2 FILLER_0_52_462 ();
 sg13g2_fill_1 FILLER_0_52_473 ();
 sg13g2_fill_4 FILLER_0_52_504 ();
 sg13g2_fill_1 FILLER_0_52_538 ();
 sg13g2_fill_1 FILLER_0_52_549 ();
 sg13g2_fill_1 FILLER_0_52_554 ();
 sg13g2_fill_4 FILLER_0_52_586 ();
 sg13g2_fill_1 FILLER_0_52_590 ();
 sg13g2_fill_2 FILLER_0_52_596 ();
 sg13g2_fill_1 FILLER_0_52_602 ();
 sg13g2_fill_8 FILLER_0_52_615 ();
 sg13g2_fill_4 FILLER_0_52_623 ();
 sg13g2_fill_1 FILLER_0_52_627 ();
 sg13g2_fill_1 FILLER_0_52_632 ();
 sg13g2_fill_1 FILLER_0_52_638 ();
 sg13g2_fill_2 FILLER_0_52_690 ();
 sg13g2_fill_2 FILLER_0_52_702 ();
 sg13g2_fill_8 FILLER_0_52_714 ();
 sg13g2_fill_2 FILLER_0_52_722 ();
 sg13g2_fill_1 FILLER_0_52_732 ();
 sg13g2_fill_2 FILLER_0_52_743 ();
 sg13g2_fill_1 FILLER_0_52_749 ();
 sg13g2_fill_2 FILLER_0_52_760 ();
 sg13g2_fill_2 FILLER_0_52_772 ();
 sg13g2_fill_1 FILLER_0_52_774 ();
 sg13g2_fill_8 FILLER_0_52_788 ();
 sg13g2_fill_2 FILLER_0_52_796 ();
 sg13g2_fill_4 FILLER_0_52_808 ();
 sg13g2_fill_8 FILLER_0_52_816 ();
 sg13g2_fill_1 FILLER_0_52_824 ();
 sg13g2_fill_1 FILLER_0_52_835 ();
 sg13g2_fill_1 FILLER_0_52_846 ();
 sg13g2_fill_1 FILLER_0_52_873 ();
 sg13g2_fill_1 FILLER_0_52_884 ();
 sg13g2_fill_8 FILLER_0_52_917 ();
 sg13g2_fill_8 FILLER_0_52_925 ();
 sg13g2_fill_8 FILLER_0_52_933 ();
 sg13g2_fill_8 FILLER_0_52_941 ();
 sg13g2_fill_8 FILLER_0_52_949 ();
 sg13g2_fill_8 FILLER_0_52_957 ();
 sg13g2_fill_8 FILLER_0_52_965 ();
 sg13g2_fill_8 FILLER_0_52_973 ();
 sg13g2_fill_8 FILLER_0_52_981 ();
 sg13g2_fill_8 FILLER_0_52_989 ();
 sg13g2_fill_8 FILLER_0_52_997 ();
 sg13g2_fill_8 FILLER_0_52_1005 ();
 sg13g2_fill_8 FILLER_0_52_1013 ();
 sg13g2_fill_8 FILLER_0_52_1021 ();
 sg13g2_fill_8 FILLER_0_52_1029 ();
 sg13g2_fill_8 FILLER_0_52_1037 ();
 sg13g2_fill_8 FILLER_0_52_1045 ();
 sg13g2_fill_8 FILLER_0_52_1053 ();
 sg13g2_fill_8 FILLER_0_52_1061 ();
 sg13g2_fill_8 FILLER_0_52_1069 ();
 sg13g2_fill_8 FILLER_0_52_1077 ();
 sg13g2_fill_8 FILLER_0_52_1085 ();
 sg13g2_fill_8 FILLER_0_52_1093 ();
 sg13g2_fill_8 FILLER_0_52_1101 ();
 sg13g2_fill_8 FILLER_0_52_1109 ();
 sg13g2_fill_8 FILLER_0_52_1117 ();
 sg13g2_fill_8 FILLER_0_52_1125 ();
 sg13g2_fill_8 FILLER_0_52_1133 ();
 sg13g2_fill_8 FILLER_0_52_1141 ();
 sg13g2_fill_8 FILLER_0_52_1149 ();
 sg13g2_fill_8 FILLER_0_52_1157 ();
 sg13g2_fill_8 FILLER_0_52_1165 ();
 sg13g2_fill_8 FILLER_0_52_1173 ();
 sg13g2_fill_8 FILLER_0_52_1181 ();
 sg13g2_fill_8 FILLER_0_52_1189 ();
 sg13g2_fill_8 FILLER_0_52_1197 ();
 sg13g2_fill_8 FILLER_0_52_1205 ();
 sg13g2_fill_8 FILLER_0_52_1213 ();
 sg13g2_decap_8 FILLER_0_52_1221 ();
 sg13g2_fill_8 FILLER_0_53_0 ();
 sg13g2_fill_4 FILLER_0_53_8 ();
 sg13g2_fill_1 FILLER_0_53_17 ();
 sg13g2_fill_2 FILLER_0_53_32 ();
 sg13g2_fill_1 FILLER_0_53_39 ();
 sg13g2_fill_1 FILLER_0_53_50 ();
 sg13g2_fill_1 FILLER_0_53_56 ();
 sg13g2_fill_2 FILLER_0_53_67 ();
 sg13g2_fill_8 FILLER_0_53_73 ();
 sg13g2_decap_8 FILLER_0_53_81 ();
 sg13g2_fill_1 FILLER_0_53_93 ();
 sg13g2_fill_1 FILLER_0_53_104 ();
 sg13g2_fill_1 FILLER_0_53_114 ();
 sg13g2_fill_2 FILLER_0_53_125 ();
 sg13g2_fill_1 FILLER_0_53_168 ();
 sg13g2_fill_2 FILLER_0_53_195 ();
 sg13g2_fill_2 FILLER_0_53_207 ();
 sg13g2_fill_8 FILLER_0_53_223 ();
 sg13g2_fill_8 FILLER_0_53_231 ();
 sg13g2_fill_8 FILLER_0_53_274 ();
 sg13g2_fill_8 FILLER_0_53_282 ();
 sg13g2_fill_4 FILLER_0_53_290 ();
 sg13g2_fill_4 FILLER_0_53_298 ();
 sg13g2_fill_1 FILLER_0_53_302 ();
 sg13g2_fill_8 FILLER_0_53_308 ();
 sg13g2_decap_8 FILLER_0_53_316 ();
 sg13g2_fill_4 FILLER_0_53_336 ();
 sg13g2_fill_2 FILLER_0_53_340 ();
 sg13g2_fill_1 FILLER_0_53_346 ();
 sg13g2_fill_8 FILLER_0_53_352 ();
 sg13g2_fill_2 FILLER_0_53_360 ();
 sg13g2_fill_2 FILLER_0_53_367 ();
 sg13g2_fill_1 FILLER_0_53_369 ();
 sg13g2_fill_8 FILLER_0_53_374 ();
 sg13g2_fill_8 FILLER_0_53_382 ();
 sg13g2_fill_8 FILLER_0_53_390 ();
 sg13g2_fill_8 FILLER_0_53_398 ();
 sg13g2_fill_8 FILLER_0_53_406 ();
 sg13g2_fill_2 FILLER_0_53_414 ();
 sg13g2_fill_1 FILLER_0_53_416 ();
 sg13g2_fill_4 FILLER_0_53_427 ();
 sg13g2_fill_4 FILLER_0_53_486 ();
 sg13g2_fill_1 FILLER_0_53_490 ();
 sg13g2_fill_8 FILLER_0_53_501 ();
 sg13g2_fill_1 FILLER_0_53_509 ();
 sg13g2_fill_1 FILLER_0_53_523 ();
 sg13g2_fill_1 FILLER_0_53_560 ();
 sg13g2_fill_8 FILLER_0_53_571 ();
 sg13g2_fill_8 FILLER_0_53_579 ();
 sg13g2_fill_8 FILLER_0_53_587 ();
 sg13g2_fill_8 FILLER_0_53_595 ();
 sg13g2_fill_8 FILLER_0_53_603 ();
 sg13g2_fill_8 FILLER_0_53_611 ();
 sg13g2_fill_8 FILLER_0_53_619 ();
 sg13g2_fill_2 FILLER_0_53_627 ();
 sg13g2_fill_2 FILLER_0_53_634 ();
 sg13g2_fill_4 FILLER_0_53_640 ();
 sg13g2_fill_8 FILLER_0_53_654 ();
 sg13g2_fill_4 FILLER_0_53_662 ();
 sg13g2_fill_2 FILLER_0_53_674 ();
 sg13g2_fill_2 FILLER_0_53_685 ();
 sg13g2_fill_1 FILLER_0_53_687 ();
 sg13g2_fill_4 FILLER_0_53_724 ();
 sg13g2_fill_1 FILLER_0_53_728 ();
 sg13g2_fill_8 FILLER_0_53_748 ();
 sg13g2_fill_4 FILLER_0_53_756 ();
 sg13g2_fill_1 FILLER_0_53_760 ();
 sg13g2_fill_8 FILLER_0_53_765 ();
 sg13g2_fill_8 FILLER_0_53_814 ();
 sg13g2_fill_8 FILLER_0_53_822 ();
 sg13g2_fill_2 FILLER_0_53_835 ();
 sg13g2_fill_2 FILLER_0_53_841 ();
 sg13g2_fill_1 FILLER_0_53_843 ();
 sg13g2_decap_8 FILLER_0_53_848 ();
 sg13g2_fill_8 FILLER_0_53_859 ();
 sg13g2_decap_8 FILLER_0_53_867 ();
 sg13g2_fill_8 FILLER_0_53_878 ();
 sg13g2_fill_4 FILLER_0_53_886 ();
 sg13g2_fill_1 FILLER_0_53_895 ();
 sg13g2_fill_8 FILLER_0_53_906 ();
 sg13g2_fill_8 FILLER_0_53_914 ();
 sg13g2_fill_8 FILLER_0_53_922 ();
 sg13g2_fill_8 FILLER_0_53_930 ();
 sg13g2_fill_8 FILLER_0_53_938 ();
 sg13g2_fill_8 FILLER_0_53_946 ();
 sg13g2_fill_8 FILLER_0_53_954 ();
 sg13g2_fill_8 FILLER_0_53_962 ();
 sg13g2_fill_8 FILLER_0_53_970 ();
 sg13g2_fill_8 FILLER_0_53_978 ();
 sg13g2_fill_8 FILLER_0_53_986 ();
 sg13g2_fill_8 FILLER_0_53_994 ();
 sg13g2_fill_8 FILLER_0_53_1002 ();
 sg13g2_fill_8 FILLER_0_53_1010 ();
 sg13g2_fill_8 FILLER_0_53_1018 ();
 sg13g2_fill_8 FILLER_0_53_1026 ();
 sg13g2_fill_8 FILLER_0_53_1034 ();
 sg13g2_fill_8 FILLER_0_53_1042 ();
 sg13g2_fill_8 FILLER_0_53_1050 ();
 sg13g2_fill_8 FILLER_0_53_1058 ();
 sg13g2_fill_8 FILLER_0_53_1066 ();
 sg13g2_fill_8 FILLER_0_53_1074 ();
 sg13g2_fill_8 FILLER_0_53_1082 ();
 sg13g2_fill_8 FILLER_0_53_1090 ();
 sg13g2_fill_8 FILLER_0_53_1098 ();
 sg13g2_fill_8 FILLER_0_53_1106 ();
 sg13g2_fill_8 FILLER_0_53_1114 ();
 sg13g2_fill_8 FILLER_0_53_1122 ();
 sg13g2_fill_8 FILLER_0_53_1130 ();
 sg13g2_fill_8 FILLER_0_53_1138 ();
 sg13g2_fill_8 FILLER_0_53_1146 ();
 sg13g2_fill_8 FILLER_0_53_1154 ();
 sg13g2_fill_8 FILLER_0_53_1162 ();
 sg13g2_fill_8 FILLER_0_53_1170 ();
 sg13g2_fill_8 FILLER_0_53_1178 ();
 sg13g2_fill_8 FILLER_0_53_1186 ();
 sg13g2_fill_8 FILLER_0_53_1194 ();
 sg13g2_fill_8 FILLER_0_53_1202 ();
 sg13g2_fill_8 FILLER_0_53_1210 ();
 sg13g2_fill_8 FILLER_0_53_1218 ();
 sg13g2_fill_2 FILLER_0_53_1226 ();
 sg13g2_decap_8 FILLER_0_54_0 ();
 sg13g2_fill_8 FILLER_0_54_26 ();
 sg13g2_fill_8 FILLER_0_54_34 ();
 sg13g2_fill_1 FILLER_0_54_42 ();
 sg13g2_fill_4 FILLER_0_54_47 ();
 sg13g2_fill_2 FILLER_0_54_51 ();
 sg13g2_fill_8 FILLER_0_54_61 ();
 sg13g2_fill_8 FILLER_0_54_69 ();
 sg13g2_fill_8 FILLER_0_54_113 ();
 sg13g2_fill_8 FILLER_0_54_121 ();
 sg13g2_fill_4 FILLER_0_54_129 ();
 sg13g2_fill_1 FILLER_0_54_137 ();
 sg13g2_fill_1 FILLER_0_54_143 ();
 sg13g2_fill_1 FILLER_0_54_148 ();
 sg13g2_fill_1 FILLER_0_54_153 ();
 sg13g2_fill_2 FILLER_0_54_164 ();
 sg13g2_fill_1 FILLER_0_54_166 ();
 sg13g2_fill_1 FILLER_0_54_176 ();
 sg13g2_fill_2 FILLER_0_54_181 ();
 sg13g2_fill_1 FILLER_0_54_198 ();
 sg13g2_decap_8 FILLER_0_54_230 ();
 sg13g2_fill_2 FILLER_0_54_290 ();
 sg13g2_fill_1 FILLER_0_54_292 ();
 sg13g2_fill_4 FILLER_0_54_319 ();
 sg13g2_fill_8 FILLER_0_54_349 ();
 sg13g2_fill_8 FILLER_0_54_357 ();
 sg13g2_fill_2 FILLER_0_54_365 ();
 sg13g2_fill_1 FILLER_0_54_393 ();
 sg13g2_fill_1 FILLER_0_54_404 ();
 sg13g2_fill_1 FILLER_0_54_410 ();
 sg13g2_fill_1 FILLER_0_54_473 ();
 sg13g2_fill_2 FILLER_0_54_479 ();
 sg13g2_fill_1 FILLER_0_54_481 ();
 sg13g2_fill_4 FILLER_0_54_508 ();
 sg13g2_fill_2 FILLER_0_54_512 ();
 sg13g2_fill_2 FILLER_0_54_523 ();
 sg13g2_fill_1 FILLER_0_54_525 ();
 sg13g2_fill_8 FILLER_0_54_557 ();
 sg13g2_fill_8 FILLER_0_54_565 ();
 sg13g2_fill_8 FILLER_0_54_573 ();
 sg13g2_fill_2 FILLER_0_54_591 ();
 sg13g2_fill_2 FILLER_0_54_624 ();
 sg13g2_fill_1 FILLER_0_54_626 ();
 sg13g2_fill_8 FILLER_0_54_653 ();
 sg13g2_fill_8 FILLER_0_54_661 ();
 sg13g2_fill_8 FILLER_0_54_669 ();
 sg13g2_fill_1 FILLER_0_54_677 ();
 sg13g2_fill_2 FILLER_0_54_683 ();
 sg13g2_fill_1 FILLER_0_54_699 ();
 sg13g2_fill_1 FILLER_0_54_710 ();
 sg13g2_fill_1 FILLER_0_54_719 ();
 sg13g2_fill_2 FILLER_0_54_724 ();
 sg13g2_fill_8 FILLER_0_54_752 ();
 sg13g2_fill_1 FILLER_0_54_760 ();
 sg13g2_decap_8 FILLER_0_54_770 ();
 sg13g2_fill_1 FILLER_0_54_781 ();
 sg13g2_fill_8 FILLER_0_54_813 ();
 sg13g2_fill_1 FILLER_0_54_821 ();
 sg13g2_fill_4 FILLER_0_54_826 ();
 sg13g2_fill_1 FILLER_0_54_830 ();
 sg13g2_fill_8 FILLER_0_54_857 ();
 sg13g2_fill_1 FILLER_0_54_865 ();
 sg13g2_fill_8 FILLER_0_54_870 ();
 sg13g2_fill_8 FILLER_0_54_878 ();
 sg13g2_fill_2 FILLER_0_54_886 ();
 sg13g2_fill_1 FILLER_0_54_888 ();
 sg13g2_fill_8 FILLER_0_54_919 ();
 sg13g2_fill_8 FILLER_0_54_927 ();
 sg13g2_fill_8 FILLER_0_54_935 ();
 sg13g2_fill_8 FILLER_0_54_943 ();
 sg13g2_fill_8 FILLER_0_54_951 ();
 sg13g2_fill_8 FILLER_0_54_959 ();
 sg13g2_fill_8 FILLER_0_54_967 ();
 sg13g2_fill_8 FILLER_0_54_975 ();
 sg13g2_fill_8 FILLER_0_54_983 ();
 sg13g2_fill_8 FILLER_0_54_991 ();
 sg13g2_fill_8 FILLER_0_54_999 ();
 sg13g2_fill_8 FILLER_0_54_1007 ();
 sg13g2_fill_8 FILLER_0_54_1015 ();
 sg13g2_fill_8 FILLER_0_54_1023 ();
 sg13g2_fill_8 FILLER_0_54_1031 ();
 sg13g2_fill_8 FILLER_0_54_1039 ();
 sg13g2_fill_8 FILLER_0_54_1047 ();
 sg13g2_fill_8 FILLER_0_54_1055 ();
 sg13g2_fill_8 FILLER_0_54_1063 ();
 sg13g2_fill_8 FILLER_0_54_1071 ();
 sg13g2_fill_8 FILLER_0_54_1079 ();
 sg13g2_fill_8 FILLER_0_54_1087 ();
 sg13g2_fill_8 FILLER_0_54_1095 ();
 sg13g2_fill_8 FILLER_0_54_1103 ();
 sg13g2_fill_8 FILLER_0_54_1111 ();
 sg13g2_fill_8 FILLER_0_54_1119 ();
 sg13g2_fill_8 FILLER_0_54_1127 ();
 sg13g2_fill_8 FILLER_0_54_1135 ();
 sg13g2_fill_8 FILLER_0_54_1143 ();
 sg13g2_fill_8 FILLER_0_54_1151 ();
 sg13g2_fill_8 FILLER_0_54_1159 ();
 sg13g2_fill_8 FILLER_0_54_1167 ();
 sg13g2_fill_8 FILLER_0_54_1175 ();
 sg13g2_fill_8 FILLER_0_54_1183 ();
 sg13g2_fill_8 FILLER_0_54_1191 ();
 sg13g2_fill_8 FILLER_0_54_1199 ();
 sg13g2_fill_8 FILLER_0_54_1207 ();
 sg13g2_fill_8 FILLER_0_54_1215 ();
 sg13g2_fill_4 FILLER_0_54_1223 ();
 sg13g2_fill_1 FILLER_0_54_1227 ();
 sg13g2_fill_1 FILLER_0_55_0 ();
 sg13g2_fill_8 FILLER_0_55_42 ();
 sg13g2_fill_2 FILLER_0_55_50 ();
 sg13g2_fill_2 FILLER_0_55_83 ();
 sg13g2_fill_2 FILLER_0_55_89 ();
 sg13g2_fill_2 FILLER_0_55_96 ();
 sg13g2_fill_2 FILLER_0_55_102 ();
 sg13g2_fill_1 FILLER_0_55_104 ();
 sg13g2_decap_8 FILLER_0_55_120 ();
 sg13g2_fill_8 FILLER_0_55_131 ();
 sg13g2_decap_8 FILLER_0_55_139 ();
 sg13g2_fill_4 FILLER_0_55_164 ();
 sg13g2_fill_8 FILLER_0_55_176 ();
 sg13g2_fill_4 FILLER_0_55_184 ();
 sg13g2_fill_2 FILLER_0_55_198 ();
 sg13g2_fill_1 FILLER_0_55_200 ();
 sg13g2_decap_8 FILLER_0_55_236 ();
 sg13g2_fill_1 FILLER_0_55_269 ();
 sg13g2_fill_2 FILLER_0_55_337 ();
 sg13g2_fill_1 FILLER_0_55_339 ();
 sg13g2_fill_4 FILLER_0_55_366 ();
 sg13g2_fill_2 FILLER_0_55_370 ();
 sg13g2_fill_2 FILLER_0_55_376 ();
 sg13g2_fill_1 FILLER_0_55_378 ();
 sg13g2_fill_1 FILLER_0_55_410 ();
 sg13g2_fill_2 FILLER_0_55_415 ();
 sg13g2_fill_4 FILLER_0_55_421 ();
 sg13g2_fill_8 FILLER_0_55_435 ();
 sg13g2_fill_2 FILLER_0_55_479 ();
 sg13g2_fill_1 FILLER_0_55_481 ();
 sg13g2_fill_8 FILLER_0_55_508 ();
 sg13g2_fill_8 FILLER_0_55_516 ();
 sg13g2_fill_8 FILLER_0_55_524 ();
 sg13g2_fill_1 FILLER_0_55_532 ();
 sg13g2_fill_1 FILLER_0_55_537 ();
 sg13g2_fill_8 FILLER_0_55_542 ();
 sg13g2_fill_8 FILLER_0_55_550 ();
 sg13g2_fill_8 FILLER_0_55_558 ();
 sg13g2_fill_4 FILLER_0_55_566 ();
 sg13g2_fill_1 FILLER_0_55_570 ();
 sg13g2_fill_2 FILLER_0_55_576 ();
 sg13g2_fill_1 FILLER_0_55_604 ();
 sg13g2_fill_2 FILLER_0_55_631 ();
 sg13g2_fill_4 FILLER_0_55_659 ();
 sg13g2_fill_4 FILLER_0_55_689 ();
 sg13g2_fill_2 FILLER_0_55_724 ();
 sg13g2_fill_1 FILLER_0_55_726 ();
 sg13g2_fill_2 FILLER_0_55_793 ();
 sg13g2_fill_8 FILLER_0_55_809 ();
 sg13g2_fill_8 FILLER_0_55_817 ();
 sg13g2_fill_8 FILLER_0_55_825 ();
 sg13g2_fill_8 FILLER_0_55_833 ();
 sg13g2_fill_8 FILLER_0_55_841 ();
 sg13g2_fill_4 FILLER_0_55_849 ();
 sg13g2_fill_1 FILLER_0_55_853 ();
 sg13g2_fill_8 FILLER_0_55_921 ();
 sg13g2_fill_8 FILLER_0_55_929 ();
 sg13g2_fill_8 FILLER_0_55_937 ();
 sg13g2_fill_8 FILLER_0_55_945 ();
 sg13g2_fill_8 FILLER_0_55_953 ();
 sg13g2_fill_8 FILLER_0_55_961 ();
 sg13g2_fill_8 FILLER_0_55_969 ();
 sg13g2_fill_8 FILLER_0_55_977 ();
 sg13g2_fill_8 FILLER_0_55_985 ();
 sg13g2_fill_8 FILLER_0_55_993 ();
 sg13g2_fill_8 FILLER_0_55_1001 ();
 sg13g2_fill_8 FILLER_0_55_1009 ();
 sg13g2_fill_8 FILLER_0_55_1017 ();
 sg13g2_fill_8 FILLER_0_55_1025 ();
 sg13g2_fill_8 FILLER_0_55_1033 ();
 sg13g2_fill_8 FILLER_0_55_1041 ();
 sg13g2_fill_8 FILLER_0_55_1049 ();
 sg13g2_fill_8 FILLER_0_55_1057 ();
 sg13g2_fill_8 FILLER_0_55_1065 ();
 sg13g2_fill_8 FILLER_0_55_1073 ();
 sg13g2_fill_8 FILLER_0_55_1081 ();
 sg13g2_fill_8 FILLER_0_55_1089 ();
 sg13g2_fill_8 FILLER_0_55_1097 ();
 sg13g2_fill_8 FILLER_0_55_1105 ();
 sg13g2_fill_8 FILLER_0_55_1113 ();
 sg13g2_fill_8 FILLER_0_55_1121 ();
 sg13g2_fill_8 FILLER_0_55_1129 ();
 sg13g2_fill_8 FILLER_0_55_1137 ();
 sg13g2_fill_8 FILLER_0_55_1145 ();
 sg13g2_fill_8 FILLER_0_55_1153 ();
 sg13g2_fill_8 FILLER_0_55_1161 ();
 sg13g2_fill_8 FILLER_0_55_1169 ();
 sg13g2_fill_8 FILLER_0_55_1177 ();
 sg13g2_fill_8 FILLER_0_55_1185 ();
 sg13g2_fill_8 FILLER_0_55_1193 ();
 sg13g2_fill_8 FILLER_0_55_1201 ();
 sg13g2_fill_8 FILLER_0_55_1209 ();
 sg13g2_fill_8 FILLER_0_55_1217 ();
 sg13g2_fill_2 FILLER_0_55_1225 ();
 sg13g2_fill_1 FILLER_0_55_1227 ();
 sg13g2_fill_1 FILLER_0_56_0 ();
 sg13g2_fill_1 FILLER_0_56_27 ();
 sg13g2_fill_8 FILLER_0_56_58 ();
 sg13g2_fill_2 FILLER_0_56_70 ();
 sg13g2_fill_1 FILLER_0_56_86 ();
 sg13g2_fill_1 FILLER_0_56_97 ();
 sg13g2_fill_1 FILLER_0_56_124 ();
 sg13g2_fill_8 FILLER_0_56_129 ();
 sg13g2_fill_8 FILLER_0_56_137 ();
 sg13g2_decap_8 FILLER_0_56_145 ();
 sg13g2_fill_1 FILLER_0_56_167 ();
 sg13g2_fill_2 FILLER_0_56_178 ();
 sg13g2_fill_2 FILLER_0_56_185 ();
 sg13g2_fill_8 FILLER_0_56_197 ();
 sg13g2_fill_8 FILLER_0_56_235 ();
 sg13g2_fill_8 FILLER_0_56_243 ();
 sg13g2_fill_4 FILLER_0_56_255 ();
 sg13g2_fill_2 FILLER_0_56_259 ();
 sg13g2_fill_2 FILLER_0_56_276 ();
 sg13g2_fill_1 FILLER_0_56_278 ();
 sg13g2_fill_1 FILLER_0_56_289 ();
 sg13g2_fill_1 FILLER_0_56_295 ();
 sg13g2_fill_1 FILLER_0_56_306 ();
 sg13g2_fill_1 FILLER_0_56_311 ();
 sg13g2_fill_1 FILLER_0_56_322 ();
 sg13g2_fill_2 FILLER_0_56_337 ();
 sg13g2_fill_1 FILLER_0_56_339 ();
 sg13g2_fill_4 FILLER_0_56_345 ();
 sg13g2_fill_4 FILLER_0_56_353 ();
 sg13g2_fill_8 FILLER_0_56_437 ();
 sg13g2_fill_1 FILLER_0_56_445 ();
 sg13g2_fill_4 FILLER_0_56_451 ();
 sg13g2_fill_1 FILLER_0_56_455 ();
 sg13g2_fill_2 FILLER_0_56_464 ();
 sg13g2_fill_1 FILLER_0_56_466 ();
 sg13g2_fill_8 FILLER_0_56_472 ();
 sg13g2_fill_2 FILLER_0_56_480 ();
 sg13g2_fill_2 FILLER_0_56_487 ();
 sg13g2_fill_8 FILLER_0_56_497 ();
 sg13g2_fill_8 FILLER_0_56_505 ();
 sg13g2_fill_8 FILLER_0_56_513 ();
 sg13g2_fill_8 FILLER_0_56_521 ();
 sg13g2_fill_8 FILLER_0_56_529 ();
 sg13g2_fill_4 FILLER_0_56_537 ();
 sg13g2_decap_8 FILLER_0_56_546 ();
 sg13g2_fill_2 FILLER_0_56_644 ();
 sg13g2_fill_2 FILLER_0_56_650 ();
 sg13g2_fill_2 FILLER_0_56_747 ();
 sg13g2_fill_4 FILLER_0_56_784 ();
 sg13g2_fill_2 FILLER_0_56_788 ();
 sg13g2_fill_1 FILLER_0_56_800 ();
 sg13g2_fill_8 FILLER_0_56_832 ();
 sg13g2_fill_8 FILLER_0_56_840 ();
 sg13g2_fill_8 FILLER_0_56_848 ();
 sg13g2_fill_8 FILLER_0_56_856 ();
 sg13g2_fill_8 FILLER_0_56_864 ();
 sg13g2_fill_1 FILLER_0_56_872 ();
 sg13g2_fill_1 FILLER_0_56_877 ();
 sg13g2_fill_2 FILLER_0_56_888 ();
 sg13g2_fill_2 FILLER_0_56_895 ();
 sg13g2_fill_2 FILLER_0_56_907 ();
 sg13g2_fill_1 FILLER_0_56_909 ();
 sg13g2_fill_8 FILLER_0_56_914 ();
 sg13g2_fill_8 FILLER_0_56_922 ();
 sg13g2_fill_8 FILLER_0_56_930 ();
 sg13g2_fill_8 FILLER_0_56_938 ();
 sg13g2_fill_8 FILLER_0_56_946 ();
 sg13g2_fill_8 FILLER_0_56_954 ();
 sg13g2_fill_8 FILLER_0_56_962 ();
 sg13g2_fill_8 FILLER_0_56_970 ();
 sg13g2_fill_8 FILLER_0_56_978 ();
 sg13g2_fill_8 FILLER_0_56_986 ();
 sg13g2_fill_8 FILLER_0_56_994 ();
 sg13g2_fill_8 FILLER_0_56_1002 ();
 sg13g2_fill_8 FILLER_0_56_1010 ();
 sg13g2_fill_8 FILLER_0_56_1018 ();
 sg13g2_fill_8 FILLER_0_56_1026 ();
 sg13g2_fill_8 FILLER_0_56_1034 ();
 sg13g2_fill_8 FILLER_0_56_1042 ();
 sg13g2_fill_8 FILLER_0_56_1050 ();
 sg13g2_fill_8 FILLER_0_56_1058 ();
 sg13g2_fill_8 FILLER_0_56_1066 ();
 sg13g2_fill_8 FILLER_0_56_1074 ();
 sg13g2_fill_8 FILLER_0_56_1082 ();
 sg13g2_fill_8 FILLER_0_56_1090 ();
 sg13g2_fill_8 FILLER_0_56_1098 ();
 sg13g2_fill_8 FILLER_0_56_1106 ();
 sg13g2_fill_8 FILLER_0_56_1114 ();
 sg13g2_fill_8 FILLER_0_56_1122 ();
 sg13g2_fill_8 FILLER_0_56_1130 ();
 sg13g2_fill_8 FILLER_0_56_1138 ();
 sg13g2_fill_8 FILLER_0_56_1146 ();
 sg13g2_fill_8 FILLER_0_56_1154 ();
 sg13g2_fill_8 FILLER_0_56_1162 ();
 sg13g2_fill_8 FILLER_0_56_1170 ();
 sg13g2_fill_8 FILLER_0_56_1178 ();
 sg13g2_fill_8 FILLER_0_56_1186 ();
 sg13g2_fill_8 FILLER_0_56_1194 ();
 sg13g2_fill_8 FILLER_0_56_1202 ();
 sg13g2_fill_8 FILLER_0_56_1210 ();
 sg13g2_fill_8 FILLER_0_56_1218 ();
 sg13g2_fill_2 FILLER_0_56_1226 ();
 sg13g2_decap_8 FILLER_0_57_0 ();
 sg13g2_fill_8 FILLER_0_57_11 ();
 sg13g2_fill_4 FILLER_0_57_24 ();
 sg13g2_fill_1 FILLER_0_57_28 ();
 sg13g2_fill_8 FILLER_0_57_43 ();
 sg13g2_fill_4 FILLER_0_57_55 ();
 sg13g2_fill_2 FILLER_0_57_59 ();
 sg13g2_fill_1 FILLER_0_57_118 ();
 sg13g2_fill_1 FILLER_0_57_132 ();
 sg13g2_fill_4 FILLER_0_57_169 ();
 sg13g2_decap_8 FILLER_0_57_199 ();
 sg13g2_fill_8 FILLER_0_57_231 ();
 sg13g2_fill_8 FILLER_0_57_239 ();
 sg13g2_fill_8 FILLER_0_57_247 ();
 sg13g2_fill_8 FILLER_0_57_255 ();
 sg13g2_decap_8 FILLER_0_57_263 ();
 sg13g2_decap_8 FILLER_0_57_274 ();
 sg13g2_fill_8 FILLER_0_57_285 ();
 sg13g2_decap_8 FILLER_0_57_293 ();
 sg13g2_fill_8 FILLER_0_57_304 ();
 sg13g2_fill_8 FILLER_0_57_312 ();
 sg13g2_decap_8 FILLER_0_57_320 ();
 sg13g2_fill_8 FILLER_0_57_332 ();
 sg13g2_fill_8 FILLER_0_57_340 ();
 sg13g2_fill_2 FILLER_0_57_348 ();
 sg13g2_fill_8 FILLER_0_57_354 ();
 sg13g2_fill_8 FILLER_0_57_362 ();
 sg13g2_fill_4 FILLER_0_57_370 ();
 sg13g2_fill_2 FILLER_0_57_374 ();
 sg13g2_fill_8 FILLER_0_57_391 ();
 sg13g2_fill_8 FILLER_0_57_399 ();
 sg13g2_decap_8 FILLER_0_57_407 ();
 sg13g2_fill_2 FILLER_0_57_418 ();
 sg13g2_fill_1 FILLER_0_57_420 ();
 sg13g2_fill_8 FILLER_0_57_441 ();
 sg13g2_fill_4 FILLER_0_57_449 ();
 sg13g2_fill_1 FILLER_0_57_453 ();
 sg13g2_fill_8 FILLER_0_57_462 ();
 sg13g2_fill_8 FILLER_0_57_470 ();
 sg13g2_fill_8 FILLER_0_57_478 ();
 sg13g2_fill_8 FILLER_0_57_491 ();
 sg13g2_fill_8 FILLER_0_57_499 ();
 sg13g2_fill_8 FILLER_0_57_507 ();
 sg13g2_fill_2 FILLER_0_57_515 ();
 sg13g2_fill_1 FILLER_0_57_517 ();
 sg13g2_fill_2 FILLER_0_57_526 ();
 sg13g2_fill_1 FILLER_0_57_528 ();
 sg13g2_decap_8 FILLER_0_57_595 ();
 sg13g2_fill_1 FILLER_0_57_607 ();
 sg13g2_fill_4 FILLER_0_57_634 ();
 sg13g2_fill_2 FILLER_0_57_638 ();
 sg13g2_fill_1 FILLER_0_57_666 ();
 sg13g2_fill_1 FILLER_0_57_671 ();
 sg13g2_fill_1 FILLER_0_57_698 ();
 sg13g2_fill_2 FILLER_0_57_704 ();
 sg13g2_fill_8 FILLER_0_57_711 ();
 sg13g2_fill_8 FILLER_0_57_719 ();
 sg13g2_fill_1 FILLER_0_57_727 ();
 sg13g2_fill_2 FILLER_0_57_732 ();
 sg13g2_fill_1 FILLER_0_57_734 ();
 sg13g2_fill_1 FILLER_0_57_754 ();
 sg13g2_fill_8 FILLER_0_57_760 ();
 sg13g2_fill_1 FILLER_0_57_768 ();
 sg13g2_fill_2 FILLER_0_57_791 ();
 sg13g2_fill_8 FILLER_0_57_829 ();
 sg13g2_fill_8 FILLER_0_57_837 ();
 sg13g2_fill_2 FILLER_0_57_845 ();
 sg13g2_fill_1 FILLER_0_57_847 ();
 sg13g2_fill_2 FILLER_0_57_852 ();
 sg13g2_fill_1 FILLER_0_57_895 ();
 sg13g2_fill_8 FILLER_0_57_901 ();
 sg13g2_fill_8 FILLER_0_57_909 ();
 sg13g2_fill_8 FILLER_0_57_917 ();
 sg13g2_fill_8 FILLER_0_57_925 ();
 sg13g2_fill_1 FILLER_0_57_933 ();
 sg13g2_fill_8 FILLER_0_57_938 ();
 sg13g2_fill_2 FILLER_0_57_946 ();
 sg13g2_fill_8 FILLER_0_57_952 ();
 sg13g2_fill_8 FILLER_0_57_960 ();
 sg13g2_fill_4 FILLER_0_57_968 ();
 sg13g2_fill_1 FILLER_0_57_972 ();
 sg13g2_fill_8 FILLER_0_57_977 ();
 sg13g2_fill_8 FILLER_0_57_985 ();
 sg13g2_fill_8 FILLER_0_57_993 ();
 sg13g2_fill_8 FILLER_0_57_1001 ();
 sg13g2_fill_8 FILLER_0_57_1009 ();
 sg13g2_fill_8 FILLER_0_57_1017 ();
 sg13g2_fill_8 FILLER_0_57_1025 ();
 sg13g2_fill_8 FILLER_0_57_1033 ();
 sg13g2_fill_8 FILLER_0_57_1041 ();
 sg13g2_fill_8 FILLER_0_57_1049 ();
 sg13g2_fill_8 FILLER_0_57_1057 ();
 sg13g2_fill_8 FILLER_0_57_1065 ();
 sg13g2_fill_8 FILLER_0_57_1073 ();
 sg13g2_fill_8 FILLER_0_57_1081 ();
 sg13g2_fill_8 FILLER_0_57_1089 ();
 sg13g2_fill_8 FILLER_0_57_1097 ();
 sg13g2_fill_8 FILLER_0_57_1105 ();
 sg13g2_fill_8 FILLER_0_57_1113 ();
 sg13g2_fill_8 FILLER_0_57_1121 ();
 sg13g2_fill_8 FILLER_0_57_1129 ();
 sg13g2_fill_8 FILLER_0_57_1137 ();
 sg13g2_fill_8 FILLER_0_57_1145 ();
 sg13g2_fill_8 FILLER_0_57_1153 ();
 sg13g2_fill_8 FILLER_0_57_1161 ();
 sg13g2_fill_8 FILLER_0_57_1169 ();
 sg13g2_fill_8 FILLER_0_57_1177 ();
 sg13g2_fill_8 FILLER_0_57_1185 ();
 sg13g2_fill_8 FILLER_0_57_1193 ();
 sg13g2_fill_8 FILLER_0_57_1201 ();
 sg13g2_fill_8 FILLER_0_57_1209 ();
 sg13g2_fill_8 FILLER_0_57_1217 ();
 sg13g2_fill_2 FILLER_0_57_1225 ();
 sg13g2_fill_1 FILLER_0_57_1227 ();
 sg13g2_decap_8 FILLER_0_58_0 ();
 sg13g2_fill_4 FILLER_0_58_41 ();
 sg13g2_fill_8 FILLER_0_58_84 ();
 sg13g2_fill_4 FILLER_0_58_92 ();
 sg13g2_fill_1 FILLER_0_58_96 ();
 sg13g2_fill_1 FILLER_0_58_109 ();
 sg13g2_fill_1 FILLER_0_58_120 ();
 sg13g2_fill_1 FILLER_0_58_147 ();
 sg13g2_fill_1 FILLER_0_58_174 ();
 sg13g2_fill_2 FILLER_0_58_201 ();
 sg13g2_fill_1 FILLER_0_58_208 ();
 sg13g2_fill_2 FILLER_0_58_235 ();
 sg13g2_fill_1 FILLER_0_58_237 ();
 sg13g2_fill_8 FILLER_0_58_264 ();
 sg13g2_fill_4 FILLER_0_58_272 ();
 sg13g2_fill_1 FILLER_0_58_276 ();
 sg13g2_fill_2 FILLER_0_58_282 ();
 sg13g2_fill_8 FILLER_0_58_293 ();
 sg13g2_fill_2 FILLER_0_58_301 ();
 sg13g2_fill_1 FILLER_0_58_313 ();
 sg13g2_fill_2 FILLER_0_58_340 ();
 sg13g2_fill_1 FILLER_0_58_342 ();
 sg13g2_fill_8 FILLER_0_58_369 ();
 sg13g2_fill_2 FILLER_0_58_377 ();
 sg13g2_fill_8 FILLER_0_58_394 ();
 sg13g2_fill_8 FILLER_0_58_402 ();
 sg13g2_fill_8 FILLER_0_58_410 ();
 sg13g2_fill_1 FILLER_0_58_418 ();
 sg13g2_fill_1 FILLER_0_58_455 ();
 sg13g2_fill_1 FILLER_0_58_460 ();
 sg13g2_fill_1 FILLER_0_58_513 ();
 sg13g2_fill_1 FILLER_0_58_540 ();
 sg13g2_fill_1 FILLER_0_58_567 ();
 sg13g2_fill_1 FILLER_0_58_573 ();
 sg13g2_fill_8 FILLER_0_58_584 ();
 sg13g2_fill_8 FILLER_0_58_592 ();
 sg13g2_fill_8 FILLER_0_58_600 ();
 sg13g2_fill_2 FILLER_0_58_608 ();
 sg13g2_fill_1 FILLER_0_58_610 ();
 sg13g2_fill_8 FILLER_0_58_625 ();
 sg13g2_fill_2 FILLER_0_58_633 ();
 sg13g2_fill_1 FILLER_0_58_635 ();
 sg13g2_fill_4 FILLER_0_58_641 ();
 sg13g2_fill_1 FILLER_0_58_645 ();
 sg13g2_fill_8 FILLER_0_58_656 ();
 sg13g2_fill_1 FILLER_0_58_664 ();
 sg13g2_fill_4 FILLER_0_58_673 ();
 sg13g2_fill_1 FILLER_0_58_677 ();
 sg13g2_fill_8 FILLER_0_58_682 ();
 sg13g2_fill_4 FILLER_0_58_690 ();
 sg13g2_fill_4 FILLER_0_58_704 ();
 sg13g2_fill_1 FILLER_0_58_708 ();
 sg13g2_fill_8 FILLER_0_58_728 ();
 sg13g2_fill_8 FILLER_0_58_736 ();
 sg13g2_fill_8 FILLER_0_58_744 ();
 sg13g2_decap_8 FILLER_0_58_752 ();
 sg13g2_fill_8 FILLER_0_58_767 ();
 sg13g2_fill_2 FILLER_0_58_775 ();
 sg13g2_fill_1 FILLER_0_58_777 ();
 sg13g2_fill_2 FILLER_0_58_812 ();
 sg13g2_fill_1 FILLER_0_58_818 ();
 sg13g2_fill_8 FILLER_0_58_823 ();
 sg13g2_fill_8 FILLER_0_58_831 ();
 sg13g2_fill_2 FILLER_0_58_904 ();
 sg13g2_fill_1 FILLER_0_58_906 ();
 sg13g2_fill_1 FILLER_0_58_933 ();
 sg13g2_fill_2 FILLER_0_58_950 ();
 sg13g2_fill_1 FILLER_0_58_952 ();
 sg13g2_decap_8 FILLER_0_58_958 ();
 sg13g2_fill_8 FILLER_0_58_991 ();
 sg13g2_fill_8 FILLER_0_58_999 ();
 sg13g2_fill_8 FILLER_0_58_1007 ();
 sg13g2_fill_8 FILLER_0_58_1015 ();
 sg13g2_fill_8 FILLER_0_58_1023 ();
 sg13g2_fill_8 FILLER_0_58_1031 ();
 sg13g2_fill_8 FILLER_0_58_1039 ();
 sg13g2_fill_8 FILLER_0_58_1047 ();
 sg13g2_fill_8 FILLER_0_58_1055 ();
 sg13g2_fill_8 FILLER_0_58_1063 ();
 sg13g2_fill_8 FILLER_0_58_1071 ();
 sg13g2_fill_8 FILLER_0_58_1079 ();
 sg13g2_fill_8 FILLER_0_58_1087 ();
 sg13g2_fill_8 FILLER_0_58_1095 ();
 sg13g2_fill_8 FILLER_0_58_1103 ();
 sg13g2_fill_8 FILLER_0_58_1111 ();
 sg13g2_fill_8 FILLER_0_58_1119 ();
 sg13g2_fill_8 FILLER_0_58_1127 ();
 sg13g2_fill_8 FILLER_0_58_1135 ();
 sg13g2_fill_8 FILLER_0_58_1143 ();
 sg13g2_fill_8 FILLER_0_58_1151 ();
 sg13g2_fill_8 FILLER_0_58_1159 ();
 sg13g2_fill_8 FILLER_0_58_1167 ();
 sg13g2_fill_8 FILLER_0_58_1175 ();
 sg13g2_fill_8 FILLER_0_58_1183 ();
 sg13g2_fill_8 FILLER_0_58_1191 ();
 sg13g2_fill_8 FILLER_0_58_1199 ();
 sg13g2_fill_8 FILLER_0_58_1207 ();
 sg13g2_fill_8 FILLER_0_58_1215 ();
 sg13g2_fill_4 FILLER_0_58_1223 ();
 sg13g2_fill_1 FILLER_0_58_1227 ();
 sg13g2_fill_1 FILLER_0_59_0 ();
 sg13g2_fill_8 FILLER_0_59_27 ();
 sg13g2_fill_8 FILLER_0_59_35 ();
 sg13g2_fill_4 FILLER_0_59_43 ();
 sg13g2_fill_2 FILLER_0_59_47 ();
 sg13g2_fill_4 FILLER_0_59_53 ();
 sg13g2_fill_1 FILLER_0_59_57 ();
 sg13g2_fill_1 FILLER_0_59_75 ();
 sg13g2_fill_4 FILLER_0_59_117 ();
 sg13g2_fill_2 FILLER_0_59_121 ();
 sg13g2_fill_2 FILLER_0_59_131 ();
 sg13g2_fill_2 FILLER_0_59_152 ();
 sg13g2_fill_1 FILLER_0_59_154 ();
 sg13g2_fill_1 FILLER_0_59_168 ();
 sg13g2_fill_2 FILLER_0_59_173 ();
 sg13g2_fill_2 FILLER_0_59_180 ();
 sg13g2_fill_8 FILLER_0_59_195 ();
 sg13g2_fill_8 FILLER_0_59_203 ();
 sg13g2_fill_4 FILLER_0_59_211 ();
 sg13g2_fill_8 FILLER_0_59_227 ();
 sg13g2_fill_4 FILLER_0_59_235 ();
 sg13g2_fill_2 FILLER_0_59_239 ();
 sg13g2_fill_1 FILLER_0_59_256 ();
 sg13g2_fill_2 FILLER_0_59_340 ();
 sg13g2_fill_2 FILLER_0_59_347 ();
 sg13g2_fill_1 FILLER_0_59_349 ();
 sg13g2_fill_1 FILLER_0_59_376 ();
 sg13g2_fill_1 FILLER_0_59_403 ();
 sg13g2_fill_2 FILLER_0_59_414 ();
 sg13g2_fill_1 FILLER_0_59_420 ();
 sg13g2_fill_1 FILLER_0_59_447 ();
 sg13g2_fill_4 FILLER_0_59_452 ();
 sg13g2_fill_1 FILLER_0_59_492 ();
 sg13g2_fill_1 FILLER_0_59_528 ();
 sg13g2_fill_1 FILLER_0_59_533 ();
 sg13g2_fill_1 FILLER_0_59_549 ();
 sg13g2_fill_2 FILLER_0_59_598 ();
 sg13g2_fill_1 FILLER_0_59_639 ();
 sg13g2_fill_8 FILLER_0_59_666 ();
 sg13g2_fill_4 FILLER_0_59_674 ();
 sg13g2_fill_1 FILLER_0_59_678 ();
 sg13g2_fill_2 FILLER_0_59_710 ();
 sg13g2_fill_1 FILLER_0_59_712 ();
 sg13g2_fill_2 FILLER_0_59_739 ();
 sg13g2_fill_8 FILLER_0_59_802 ();
 sg13g2_fill_8 FILLER_0_59_810 ();
 sg13g2_fill_8 FILLER_0_59_818 ();
 sg13g2_fill_8 FILLER_0_59_826 ();
 sg13g2_fill_4 FILLER_0_59_834 ();
 sg13g2_fill_4 FILLER_0_59_842 ();
 sg13g2_fill_8 FILLER_0_59_859 ();
 sg13g2_fill_1 FILLER_0_59_884 ();
 sg13g2_fill_2 FILLER_0_59_895 ();
 sg13g2_fill_2 FILLER_0_59_923 ();
 sg13g2_fill_2 FILLER_0_59_951 ();
 sg13g2_fill_1 FILLER_0_59_953 ();
 sg13g2_fill_8 FILLER_0_59_964 ();
 sg13g2_fill_8 FILLER_0_59_976 ();
 sg13g2_fill_8 FILLER_0_59_984 ();
 sg13g2_fill_8 FILLER_0_59_992 ();
 sg13g2_fill_8 FILLER_0_59_1000 ();
 sg13g2_fill_8 FILLER_0_59_1008 ();
 sg13g2_fill_8 FILLER_0_59_1016 ();
 sg13g2_fill_8 FILLER_0_59_1024 ();
 sg13g2_fill_8 FILLER_0_59_1032 ();
 sg13g2_fill_8 FILLER_0_59_1040 ();
 sg13g2_fill_8 FILLER_0_59_1048 ();
 sg13g2_fill_8 FILLER_0_59_1056 ();
 sg13g2_fill_8 FILLER_0_59_1064 ();
 sg13g2_fill_8 FILLER_0_59_1072 ();
 sg13g2_fill_8 FILLER_0_59_1080 ();
 sg13g2_fill_8 FILLER_0_59_1088 ();
 sg13g2_fill_8 FILLER_0_59_1096 ();
 sg13g2_fill_8 FILLER_0_59_1104 ();
 sg13g2_fill_8 FILLER_0_59_1112 ();
 sg13g2_fill_8 FILLER_0_59_1120 ();
 sg13g2_fill_8 FILLER_0_59_1128 ();
 sg13g2_fill_8 FILLER_0_59_1136 ();
 sg13g2_fill_8 FILLER_0_59_1144 ();
 sg13g2_fill_8 FILLER_0_59_1152 ();
 sg13g2_fill_8 FILLER_0_59_1160 ();
 sg13g2_fill_8 FILLER_0_59_1168 ();
 sg13g2_fill_8 FILLER_0_59_1176 ();
 sg13g2_fill_8 FILLER_0_59_1184 ();
 sg13g2_fill_8 FILLER_0_59_1192 ();
 sg13g2_fill_8 FILLER_0_59_1200 ();
 sg13g2_fill_8 FILLER_0_59_1208 ();
 sg13g2_fill_8 FILLER_0_59_1216 ();
 sg13g2_fill_4 FILLER_0_59_1224 ();
 sg13g2_fill_2 FILLER_0_60_32 ();
 sg13g2_fill_1 FILLER_0_60_44 ();
 sg13g2_fill_2 FILLER_0_60_50 ();
 sg13g2_fill_2 FILLER_0_60_78 ();
 sg13g2_fill_1 FILLER_0_60_80 ();
 sg13g2_fill_4 FILLER_0_60_91 ();
 sg13g2_fill_1 FILLER_0_60_95 ();
 sg13g2_fill_8 FILLER_0_60_127 ();
 sg13g2_fill_1 FILLER_0_60_135 ();
 sg13g2_fill_4 FILLER_0_60_141 ();
 sg13g2_fill_2 FILLER_0_60_154 ();
 sg13g2_fill_1 FILLER_0_60_156 ();
 sg13g2_fill_8 FILLER_0_60_161 ();
 sg13g2_fill_8 FILLER_0_60_169 ();
 sg13g2_fill_2 FILLER_0_60_177 ();
 sg13g2_fill_1 FILLER_0_60_179 ();
 sg13g2_fill_2 FILLER_0_60_188 ();
 sg13g2_fill_1 FILLER_0_60_190 ();
 sg13g2_fill_2 FILLER_0_60_199 ();
 sg13g2_fill_1 FILLER_0_60_201 ();
 sg13g2_fill_2 FILLER_0_60_232 ();
 sg13g2_fill_1 FILLER_0_60_234 ();
 sg13g2_fill_1 FILLER_0_60_315 ();
 sg13g2_fill_2 FILLER_0_60_320 ();
 sg13g2_fill_2 FILLER_0_60_326 ();
 sg13g2_fill_8 FILLER_0_60_436 ();
 sg13g2_fill_8 FILLER_0_60_444 ();
 sg13g2_fill_8 FILLER_0_60_452 ();
 sg13g2_fill_2 FILLER_0_60_460 ();
 sg13g2_fill_1 FILLER_0_60_462 ();
 sg13g2_fill_2 FILLER_0_60_501 ();
 sg13g2_fill_4 FILLER_0_60_528 ();
 sg13g2_fill_1 FILLER_0_60_532 ();
 sg13g2_fill_2 FILLER_0_60_537 ();
 sg13g2_fill_4 FILLER_0_60_559 ();
 sg13g2_fill_2 FILLER_0_60_563 ();
 sg13g2_fill_1 FILLER_0_60_601 ();
 sg13g2_fill_1 FILLER_0_60_610 ();
 sg13g2_fill_1 FILLER_0_60_637 ();
 sg13g2_fill_2 FILLER_0_60_664 ();
 sg13g2_fill_1 FILLER_0_60_697 ();
 sg13g2_fill_2 FILLER_0_60_702 ();
 sg13g2_fill_1 FILLER_0_60_704 ();
 sg13g2_fill_1 FILLER_0_60_715 ();
 sg13g2_fill_4 FILLER_0_60_747 ();
 sg13g2_fill_2 FILLER_0_60_751 ();
 sg13g2_fill_4 FILLER_0_60_757 ();
 sg13g2_fill_2 FILLER_0_60_761 ();
 sg13g2_fill_8 FILLER_0_60_773 ();
 sg13g2_fill_1 FILLER_0_60_781 ();
 sg13g2_fill_4 FILLER_0_60_786 ();
 sg13g2_fill_2 FILLER_0_60_790 ();
 sg13g2_fill_4 FILLER_0_60_823 ();
 sg13g2_fill_4 FILLER_0_60_861 ();
 sg13g2_fill_2 FILLER_0_60_865 ();
 sg13g2_fill_2 FILLER_0_60_877 ();
 sg13g2_fill_8 FILLER_0_60_883 ();
 sg13g2_fill_1 FILLER_0_60_891 ();
 sg13g2_fill_2 FILLER_0_60_931 ();
 sg13g2_fill_1 FILLER_0_60_933 ();
 sg13g2_fill_8 FILLER_0_60_991 ();
 sg13g2_fill_8 FILLER_0_60_999 ();
 sg13g2_fill_8 FILLER_0_60_1007 ();
 sg13g2_fill_8 FILLER_0_60_1015 ();
 sg13g2_fill_8 FILLER_0_60_1023 ();
 sg13g2_fill_8 FILLER_0_60_1031 ();
 sg13g2_fill_8 FILLER_0_60_1039 ();
 sg13g2_fill_8 FILLER_0_60_1047 ();
 sg13g2_fill_8 FILLER_0_60_1055 ();
 sg13g2_fill_8 FILLER_0_60_1063 ();
 sg13g2_fill_8 FILLER_0_60_1071 ();
 sg13g2_fill_8 FILLER_0_60_1079 ();
 sg13g2_fill_8 FILLER_0_60_1087 ();
 sg13g2_fill_8 FILLER_0_60_1095 ();
 sg13g2_fill_8 FILLER_0_60_1103 ();
 sg13g2_fill_8 FILLER_0_60_1111 ();
 sg13g2_fill_8 FILLER_0_60_1119 ();
 sg13g2_fill_8 FILLER_0_60_1127 ();
 sg13g2_fill_8 FILLER_0_60_1135 ();
 sg13g2_fill_8 FILLER_0_60_1143 ();
 sg13g2_fill_8 FILLER_0_60_1151 ();
 sg13g2_fill_8 FILLER_0_60_1159 ();
 sg13g2_fill_8 FILLER_0_60_1167 ();
 sg13g2_fill_8 FILLER_0_60_1175 ();
 sg13g2_fill_8 FILLER_0_60_1183 ();
 sg13g2_fill_8 FILLER_0_60_1191 ();
 sg13g2_fill_8 FILLER_0_60_1199 ();
 sg13g2_fill_8 FILLER_0_60_1207 ();
 sg13g2_fill_8 FILLER_0_60_1215 ();
 sg13g2_fill_4 FILLER_0_60_1223 ();
 sg13g2_fill_1 FILLER_0_60_1227 ();
 sg13g2_fill_1 FILLER_0_61_0 ();
 sg13g2_decap_8 FILLER_0_61_27 ();
 sg13g2_fill_1 FILLER_0_61_60 ();
 sg13g2_fill_2 FILLER_0_61_106 ();
 sg13g2_fill_8 FILLER_0_61_112 ();
 sg13g2_fill_8 FILLER_0_61_120 ();
 sg13g2_decap_8 FILLER_0_61_128 ();
 sg13g2_fill_2 FILLER_0_61_165 ();
 sg13g2_fill_8 FILLER_0_61_228 ();
 sg13g2_decap_8 FILLER_0_61_236 ();
 sg13g2_fill_1 FILLER_0_61_252 ();
 sg13g2_fill_1 FILLER_0_61_263 ();
 sg13g2_fill_1 FILLER_0_61_268 ();
 sg13g2_fill_1 FILLER_0_61_274 ();
 sg13g2_fill_2 FILLER_0_61_301 ();
 sg13g2_fill_8 FILLER_0_61_313 ();
 sg13g2_fill_8 FILLER_0_61_321 ();
 sg13g2_fill_8 FILLER_0_61_358 ();
 sg13g2_fill_8 FILLER_0_61_366 ();
 sg13g2_fill_2 FILLER_0_61_374 ();
 sg13g2_fill_1 FILLER_0_61_376 ();
 sg13g2_fill_1 FILLER_0_61_399 ();
 sg13g2_fill_2 FILLER_0_61_410 ();
 sg13g2_fill_1 FILLER_0_61_412 ();
 sg13g2_fill_2 FILLER_0_61_418 ();
 sg13g2_fill_1 FILLER_0_61_420 ();
 sg13g2_fill_8 FILLER_0_61_425 ();
 sg13g2_fill_8 FILLER_0_61_433 ();
 sg13g2_fill_8 FILLER_0_61_441 ();
 sg13g2_fill_8 FILLER_0_61_449 ();
 sg13g2_fill_4 FILLER_0_61_457 ();
 sg13g2_fill_8 FILLER_0_61_465 ();
 sg13g2_fill_8 FILLER_0_61_483 ();
 sg13g2_fill_8 FILLER_0_61_491 ();
 sg13g2_fill_8 FILLER_0_61_499 ();
 sg13g2_fill_8 FILLER_0_61_507 ();
 sg13g2_fill_2 FILLER_0_61_515 ();
 sg13g2_fill_8 FILLER_0_61_525 ();
 sg13g2_fill_4 FILLER_0_61_533 ();
 sg13g2_fill_2 FILLER_0_61_537 ();
 sg13g2_fill_2 FILLER_0_61_555 ();
 sg13g2_fill_2 FILLER_0_61_562 ();
 sg13g2_fill_1 FILLER_0_61_564 ();
 sg13g2_fill_1 FILLER_0_61_591 ();
 sg13g2_fill_8 FILLER_0_61_596 ();
 sg13g2_fill_1 FILLER_0_61_604 ();
 sg13g2_fill_1 FILLER_0_61_632 ();
 sg13g2_fill_1 FILLER_0_61_643 ();
 sg13g2_fill_2 FILLER_0_61_658 ();
 sg13g2_fill_1 FILLER_0_61_660 ();
 sg13g2_fill_8 FILLER_0_61_671 ();
 sg13g2_fill_8 FILLER_0_61_683 ();
 sg13g2_fill_8 FILLER_0_61_691 ();
 sg13g2_fill_8 FILLER_0_61_699 ();
 sg13g2_fill_1 FILLER_0_61_707 ();
 sg13g2_fill_2 FILLER_0_61_735 ();
 sg13g2_fill_8 FILLER_0_61_777 ();
 sg13g2_fill_2 FILLER_0_61_785 ();
 sg13g2_fill_1 FILLER_0_61_787 ();
 sg13g2_fill_4 FILLER_0_61_843 ();
 sg13g2_fill_1 FILLER_0_61_847 ();
 sg13g2_fill_1 FILLER_0_61_874 ();
 sg13g2_fill_8 FILLER_0_61_894 ();
 sg13g2_fill_8 FILLER_0_61_902 ();
 sg13g2_fill_2 FILLER_0_61_910 ();
 sg13g2_fill_1 FILLER_0_61_912 ();
 sg13g2_decap_8 FILLER_0_61_917 ();
 sg13g2_fill_2 FILLER_0_61_929 ();
 sg13g2_fill_8 FILLER_0_61_992 ();
 sg13g2_fill_8 FILLER_0_61_1000 ();
 sg13g2_fill_8 FILLER_0_61_1008 ();
 sg13g2_fill_8 FILLER_0_61_1016 ();
 sg13g2_fill_8 FILLER_0_61_1024 ();
 sg13g2_fill_8 FILLER_0_61_1032 ();
 sg13g2_fill_8 FILLER_0_61_1040 ();
 sg13g2_fill_8 FILLER_0_61_1048 ();
 sg13g2_fill_8 FILLER_0_61_1056 ();
 sg13g2_fill_8 FILLER_0_61_1064 ();
 sg13g2_fill_8 FILLER_0_61_1072 ();
 sg13g2_fill_8 FILLER_0_61_1080 ();
 sg13g2_fill_8 FILLER_0_61_1088 ();
 sg13g2_fill_8 FILLER_0_61_1096 ();
 sg13g2_fill_8 FILLER_0_61_1104 ();
 sg13g2_fill_8 FILLER_0_61_1112 ();
 sg13g2_fill_8 FILLER_0_61_1120 ();
 sg13g2_fill_8 FILLER_0_61_1128 ();
 sg13g2_fill_8 FILLER_0_61_1136 ();
 sg13g2_fill_8 FILLER_0_61_1144 ();
 sg13g2_fill_8 FILLER_0_61_1152 ();
 sg13g2_fill_8 FILLER_0_61_1160 ();
 sg13g2_fill_8 FILLER_0_61_1168 ();
 sg13g2_fill_8 FILLER_0_61_1176 ();
 sg13g2_fill_8 FILLER_0_61_1184 ();
 sg13g2_fill_8 FILLER_0_61_1192 ();
 sg13g2_fill_8 FILLER_0_61_1200 ();
 sg13g2_fill_8 FILLER_0_61_1208 ();
 sg13g2_fill_8 FILLER_0_61_1216 ();
 sg13g2_fill_4 FILLER_0_61_1224 ();
 sg13g2_fill_8 FILLER_0_62_0 ();
 sg13g2_fill_8 FILLER_0_62_8 ();
 sg13g2_fill_4 FILLER_0_62_16 ();
 sg13g2_fill_1 FILLER_0_62_20 ();
 sg13g2_fill_8 FILLER_0_62_87 ();
 sg13g2_decap_8 FILLER_0_62_95 ();
 sg13g2_fill_4 FILLER_0_62_133 ();
 sg13g2_fill_1 FILLER_0_62_145 ();
 sg13g2_fill_1 FILLER_0_62_150 ();
 sg13g2_fill_1 FILLER_0_62_177 ();
 sg13g2_fill_2 FILLER_0_62_204 ();
 sg13g2_fill_2 FILLER_0_62_216 ();
 sg13g2_fill_2 FILLER_0_62_244 ();
 sg13g2_fill_1 FILLER_0_62_246 ();
 sg13g2_fill_8 FILLER_0_62_251 ();
 sg13g2_fill_2 FILLER_0_62_259 ();
 sg13g2_fill_1 FILLER_0_62_271 ();
 sg13g2_fill_1 FILLER_0_62_285 ();
 sg13g2_fill_2 FILLER_0_62_291 ();
 sg13g2_fill_1 FILLER_0_62_293 ();
 sg13g2_fill_8 FILLER_0_62_312 ();
 sg13g2_fill_4 FILLER_0_62_320 ();
 sg13g2_fill_1 FILLER_0_62_324 ();
 sg13g2_fill_4 FILLER_0_62_335 ();
 sg13g2_fill_2 FILLER_0_62_339 ();
 sg13g2_fill_2 FILLER_0_62_398 ();
 sg13g2_fill_8 FILLER_0_62_425 ();
 sg13g2_fill_8 FILLER_0_62_433 ();
 sg13g2_fill_8 FILLER_0_62_441 ();
 sg13g2_fill_4 FILLER_0_62_449 ();
 sg13g2_fill_1 FILLER_0_62_453 ();
 sg13g2_fill_1 FILLER_0_62_485 ();
 sg13g2_fill_8 FILLER_0_62_500 ();
 sg13g2_fill_2 FILLER_0_62_508 ();
 sg13g2_fill_1 FILLER_0_62_540 ();
 sg13g2_fill_8 FILLER_0_62_555 ();
 sg13g2_fill_1 FILLER_0_62_563 ();
 sg13g2_fill_4 FILLER_0_62_568 ();
 sg13g2_fill_4 FILLER_0_62_576 ();
 sg13g2_fill_2 FILLER_0_62_580 ();
 sg13g2_fill_8 FILLER_0_62_586 ();
 sg13g2_fill_8 FILLER_0_62_594 ();
 sg13g2_fill_4 FILLER_0_62_602 ();
 sg13g2_fill_2 FILLER_0_62_606 ();
 sg13g2_fill_2 FILLER_0_62_612 ();
 sg13g2_fill_8 FILLER_0_62_618 ();
 sg13g2_fill_8 FILLER_0_62_636 ();
 sg13g2_fill_2 FILLER_0_62_644 ();
 sg13g2_fill_8 FILLER_0_62_650 ();
 sg13g2_fill_8 FILLER_0_62_658 ();
 sg13g2_fill_1 FILLER_0_62_692 ();
 sg13g2_fill_4 FILLER_0_62_703 ();
 sg13g2_fill_8 FILLER_0_62_737 ();
 sg13g2_fill_2 FILLER_0_62_745 ();
 sg13g2_fill_4 FILLER_0_62_782 ();
 sg13g2_fill_2 FILLER_0_62_786 ();
 sg13g2_fill_1 FILLER_0_62_822 ();
 sg13g2_fill_2 FILLER_0_62_847 ();
 sg13g2_fill_2 FILLER_0_62_864 ();
 sg13g2_fill_1 FILLER_0_62_866 ();
 sg13g2_fill_2 FILLER_0_62_903 ();
 sg13g2_fill_8 FILLER_0_62_909 ();
 sg13g2_fill_8 FILLER_0_62_917 ();
 sg13g2_fill_2 FILLER_0_62_934 ();
 sg13g2_fill_1 FILLER_0_62_936 ();
 sg13g2_fill_1 FILLER_0_62_941 ();
 sg13g2_fill_4 FILLER_0_62_946 ();
 sg13g2_fill_2 FILLER_0_62_954 ();
 sg13g2_fill_1 FILLER_0_62_956 ();
 sg13g2_fill_1 FILLER_0_62_972 ();
 sg13g2_fill_8 FILLER_0_62_977 ();
 sg13g2_fill_8 FILLER_0_62_985 ();
 sg13g2_fill_8 FILLER_0_62_993 ();
 sg13g2_fill_8 FILLER_0_62_1001 ();
 sg13g2_fill_8 FILLER_0_62_1009 ();
 sg13g2_fill_8 FILLER_0_62_1017 ();
 sg13g2_fill_8 FILLER_0_62_1025 ();
 sg13g2_fill_8 FILLER_0_62_1033 ();
 sg13g2_fill_8 FILLER_0_62_1041 ();
 sg13g2_fill_8 FILLER_0_62_1049 ();
 sg13g2_fill_8 FILLER_0_62_1057 ();
 sg13g2_fill_8 FILLER_0_62_1065 ();
 sg13g2_fill_8 FILLER_0_62_1073 ();
 sg13g2_fill_8 FILLER_0_62_1081 ();
 sg13g2_fill_8 FILLER_0_62_1089 ();
 sg13g2_fill_8 FILLER_0_62_1097 ();
 sg13g2_fill_8 FILLER_0_62_1105 ();
 sg13g2_fill_8 FILLER_0_62_1113 ();
 sg13g2_fill_8 FILLER_0_62_1121 ();
 sg13g2_fill_8 FILLER_0_62_1129 ();
 sg13g2_fill_8 FILLER_0_62_1137 ();
 sg13g2_fill_8 FILLER_0_62_1145 ();
 sg13g2_fill_8 FILLER_0_62_1153 ();
 sg13g2_fill_8 FILLER_0_62_1161 ();
 sg13g2_fill_8 FILLER_0_62_1169 ();
 sg13g2_fill_8 FILLER_0_62_1177 ();
 sg13g2_fill_8 FILLER_0_62_1185 ();
 sg13g2_fill_8 FILLER_0_62_1193 ();
 sg13g2_fill_8 FILLER_0_62_1201 ();
 sg13g2_fill_8 FILLER_0_62_1209 ();
 sg13g2_fill_8 FILLER_0_62_1217 ();
 sg13g2_fill_2 FILLER_0_62_1225 ();
 sg13g2_fill_1 FILLER_0_62_1227 ();
 sg13g2_fill_8 FILLER_0_63_0 ();
 sg13g2_fill_8 FILLER_0_63_8 ();
 sg13g2_fill_8 FILLER_0_63_16 ();
 sg13g2_fill_2 FILLER_0_63_24 ();
 sg13g2_fill_8 FILLER_0_63_30 ();
 sg13g2_fill_2 FILLER_0_63_38 ();
 sg13g2_fill_1 FILLER_0_63_40 ();
 sg13g2_fill_8 FILLER_0_63_45 ();
 sg13g2_fill_8 FILLER_0_63_53 ();
 sg13g2_fill_8 FILLER_0_63_61 ();
 sg13g2_fill_8 FILLER_0_63_69 ();
 sg13g2_fill_8 FILLER_0_63_77 ();
 sg13g2_fill_2 FILLER_0_63_90 ();
 sg13g2_fill_1 FILLER_0_63_96 ();
 sg13g2_fill_2 FILLER_0_63_117 ();
 sg13g2_fill_1 FILLER_0_63_119 ();
 sg13g2_fill_1 FILLER_0_63_150 ();
 sg13g2_fill_1 FILLER_0_63_161 ();
 sg13g2_fill_1 FILLER_0_63_177 ();
 sg13g2_fill_2 FILLER_0_63_183 ();
 sg13g2_fill_1 FILLER_0_63_185 ();
 sg13g2_fill_4 FILLER_0_63_190 ();
 sg13g2_fill_2 FILLER_0_63_194 ();
 sg13g2_fill_8 FILLER_0_63_200 ();
 sg13g2_decap_8 FILLER_0_63_208 ();
 sg13g2_decap_8 FILLER_0_63_220 ();
 sg13g2_decap_8 FILLER_0_63_231 ();
 sg13g2_fill_4 FILLER_0_63_264 ();
 sg13g2_fill_1 FILLER_0_63_277 ();
 sg13g2_fill_1 FILLER_0_63_282 ();
 sg13g2_fill_4 FILLER_0_63_309 ();
 sg13g2_decap_8 FILLER_0_63_317 ();
 sg13g2_fill_8 FILLER_0_63_336 ();
 sg13g2_fill_4 FILLER_0_63_344 ();
 sg13g2_fill_1 FILLER_0_63_374 ();
 sg13g2_fill_2 FILLER_0_63_383 ();
 sg13g2_fill_1 FILLER_0_63_385 ();
 sg13g2_fill_4 FILLER_0_63_394 ();
 sg13g2_fill_1 FILLER_0_63_398 ();
 sg13g2_fill_4 FILLER_0_63_456 ();
 sg13g2_fill_1 FILLER_0_63_486 ();
 sg13g2_fill_1 FILLER_0_63_513 ();
 sg13g2_fill_4 FILLER_0_63_523 ();
 sg13g2_fill_2 FILLER_0_63_527 ();
 sg13g2_fill_8 FILLER_0_63_555 ();
 sg13g2_fill_4 FILLER_0_63_563 ();
 sg13g2_fill_8 FILLER_0_63_577 ();
 sg13g2_fill_4 FILLER_0_63_585 ();
 sg13g2_fill_2 FILLER_0_63_599 ();
 sg13g2_fill_2 FILLER_0_63_605 ();
 sg13g2_fill_4 FILLER_0_63_612 ();
 sg13g2_fill_4 FILLER_0_63_626 ();
 sg13g2_fill_1 FILLER_0_63_630 ();
 sg13g2_fill_2 FILLER_0_63_636 ();
 sg13g2_fill_1 FILLER_0_63_638 ();
 sg13g2_fill_8 FILLER_0_63_643 ();
 sg13g2_fill_8 FILLER_0_63_651 ();
 sg13g2_fill_8 FILLER_0_63_659 ();
 sg13g2_fill_2 FILLER_0_63_667 ();
 sg13g2_fill_1 FILLER_0_63_669 ();
 sg13g2_fill_1 FILLER_0_63_674 ();
 sg13g2_fill_2 FILLER_0_63_705 ();
 sg13g2_fill_1 FILLER_0_63_707 ();
 sg13g2_fill_8 FILLER_0_63_723 ();
 sg13g2_decap_8 FILLER_0_63_731 ();
 sg13g2_fill_1 FILLER_0_63_774 ();
 sg13g2_fill_8 FILLER_0_63_806 ();
 sg13g2_fill_8 FILLER_0_63_818 ();
 sg13g2_fill_2 FILLER_0_63_826 ();
 sg13g2_fill_8 FILLER_0_63_847 ();
 sg13g2_fill_8 FILLER_0_63_855 ();
 sg13g2_fill_2 FILLER_0_63_889 ();
 sg13g2_decap_8 FILLER_0_63_917 ();
 sg13g2_fill_4 FILLER_0_63_955 ();
 sg13g2_fill_2 FILLER_0_63_959 ();
 sg13g2_fill_2 FILLER_0_63_966 ();
 sg13g2_fill_1 FILLER_0_63_968 ();
 sg13g2_fill_8 FILLER_0_63_995 ();
 sg13g2_fill_8 FILLER_0_63_1003 ();
 sg13g2_fill_8 FILLER_0_63_1011 ();
 sg13g2_fill_8 FILLER_0_63_1019 ();
 sg13g2_fill_8 FILLER_0_63_1027 ();
 sg13g2_fill_8 FILLER_0_63_1035 ();
 sg13g2_fill_8 FILLER_0_63_1043 ();
 sg13g2_fill_8 FILLER_0_63_1051 ();
 sg13g2_fill_8 FILLER_0_63_1059 ();
 sg13g2_fill_8 FILLER_0_63_1067 ();
 sg13g2_fill_8 FILLER_0_63_1075 ();
 sg13g2_fill_8 FILLER_0_63_1083 ();
 sg13g2_fill_8 FILLER_0_63_1091 ();
 sg13g2_fill_8 FILLER_0_63_1099 ();
 sg13g2_fill_8 FILLER_0_63_1107 ();
 sg13g2_fill_8 FILLER_0_63_1115 ();
 sg13g2_fill_8 FILLER_0_63_1123 ();
 sg13g2_fill_8 FILLER_0_63_1131 ();
 sg13g2_fill_8 FILLER_0_63_1139 ();
 sg13g2_fill_8 FILLER_0_63_1147 ();
 sg13g2_fill_8 FILLER_0_63_1155 ();
 sg13g2_fill_8 FILLER_0_63_1163 ();
 sg13g2_fill_8 FILLER_0_63_1171 ();
 sg13g2_fill_8 FILLER_0_63_1179 ();
 sg13g2_fill_8 FILLER_0_63_1187 ();
 sg13g2_fill_8 FILLER_0_63_1195 ();
 sg13g2_fill_8 FILLER_0_63_1203 ();
 sg13g2_fill_8 FILLER_0_63_1211 ();
 sg13g2_fill_8 FILLER_0_63_1219 ();
 sg13g2_fill_1 FILLER_0_63_1227 ();
 sg13g2_fill_8 FILLER_0_64_0 ();
 sg13g2_fill_8 FILLER_0_64_8 ();
 sg13g2_fill_8 FILLER_0_64_16 ();
 sg13g2_fill_8 FILLER_0_64_24 ();
 sg13g2_fill_8 FILLER_0_64_32 ();
 sg13g2_fill_8 FILLER_0_64_40 ();
 sg13g2_fill_8 FILLER_0_64_48 ();
 sg13g2_fill_1 FILLER_0_64_56 ();
 sg13g2_fill_4 FILLER_0_64_67 ();
 sg13g2_fill_1 FILLER_0_64_71 ();
 sg13g2_fill_2 FILLER_0_64_80 ();
 sg13g2_fill_1 FILLER_0_64_82 ();
 sg13g2_fill_2 FILLER_0_64_109 ();
 sg13g2_fill_2 FILLER_0_64_119 ();
 sg13g2_fill_8 FILLER_0_64_141 ();
 sg13g2_fill_1 FILLER_0_64_149 ();
 sg13g2_fill_2 FILLER_0_64_180 ();
 sg13g2_decap_8 FILLER_0_64_187 ();
 sg13g2_fill_1 FILLER_0_64_225 ();
 sg13g2_fill_2 FILLER_0_64_252 ();
 sg13g2_fill_2 FILLER_0_64_264 ();
 sg13g2_fill_2 FILLER_0_64_276 ();
 sg13g2_fill_2 FILLER_0_64_292 ();
 sg13g2_fill_1 FILLER_0_64_294 ();
 sg13g2_fill_1 FILLER_0_64_351 ();
 sg13g2_fill_8 FILLER_0_64_356 ();
 sg13g2_fill_8 FILLER_0_64_364 ();
 sg13g2_fill_8 FILLER_0_64_372 ();
 sg13g2_fill_2 FILLER_0_64_380 ();
 sg13g2_fill_1 FILLER_0_64_382 ();
 sg13g2_fill_8 FILLER_0_64_387 ();
 sg13g2_fill_8 FILLER_0_64_395 ();
 sg13g2_fill_4 FILLER_0_64_403 ();
 sg13g2_fill_1 FILLER_0_64_407 ();
 sg13g2_fill_4 FILLER_0_64_464 ();
 sg13g2_fill_1 FILLER_0_64_468 ();
 sg13g2_fill_2 FILLER_0_64_478 ();
 sg13g2_fill_2 FILLER_0_64_490 ();
 sg13g2_fill_1 FILLER_0_64_492 ();
 sg13g2_fill_2 FILLER_0_64_498 ();
 sg13g2_fill_1 FILLER_0_64_500 ();
 sg13g2_fill_2 FILLER_0_64_509 ();
 sg13g2_fill_4 FILLER_0_64_521 ();
 sg13g2_fill_2 FILLER_0_64_530 ();
 sg13g2_fill_2 FILLER_0_64_550 ();
 sg13g2_fill_1 FILLER_0_64_578 ();
 sg13g2_fill_1 FILLER_0_64_584 ();
 sg13g2_fill_1 FILLER_0_64_599 ();
 sg13g2_fill_1 FILLER_0_64_626 ();
 sg13g2_fill_4 FILLER_0_64_658 ();
 sg13g2_fill_2 FILLER_0_64_662 ();
 sg13g2_fill_2 FILLER_0_64_672 ();
 sg13g2_fill_1 FILLER_0_64_679 ();
 sg13g2_fill_1 FILLER_0_64_685 ();
 sg13g2_fill_2 FILLER_0_64_709 ();
 sg13g2_fill_1 FILLER_0_64_745 ();
 sg13g2_fill_4 FILLER_0_64_750 ();
 sg13g2_fill_2 FILLER_0_64_754 ();
 sg13g2_fill_4 FILLER_0_64_761 ();
 sg13g2_fill_2 FILLER_0_64_765 ();
 sg13g2_fill_8 FILLER_0_64_802 ();
 sg13g2_fill_8 FILLER_0_64_810 ();
 sg13g2_fill_2 FILLER_0_64_818 ();
 sg13g2_fill_1 FILLER_0_64_820 ();
 sg13g2_fill_2 FILLER_0_64_861 ();
 sg13g2_fill_1 FILLER_0_64_863 ();
 sg13g2_fill_1 FILLER_0_64_926 ();
 sg13g2_fill_8 FILLER_0_64_994 ();
 sg13g2_fill_8 FILLER_0_64_1002 ();
 sg13g2_fill_8 FILLER_0_64_1010 ();
 sg13g2_fill_8 FILLER_0_64_1018 ();
 sg13g2_fill_8 FILLER_0_64_1026 ();
 sg13g2_fill_8 FILLER_0_64_1034 ();
 sg13g2_fill_8 FILLER_0_64_1042 ();
 sg13g2_fill_8 FILLER_0_64_1050 ();
 sg13g2_fill_8 FILLER_0_64_1058 ();
 sg13g2_fill_8 FILLER_0_64_1066 ();
 sg13g2_fill_8 FILLER_0_64_1074 ();
 sg13g2_fill_8 FILLER_0_64_1082 ();
 sg13g2_fill_8 FILLER_0_64_1090 ();
 sg13g2_fill_8 FILLER_0_64_1098 ();
 sg13g2_fill_8 FILLER_0_64_1106 ();
 sg13g2_fill_8 FILLER_0_64_1114 ();
 sg13g2_fill_8 FILLER_0_64_1122 ();
 sg13g2_fill_8 FILLER_0_64_1130 ();
 sg13g2_fill_8 FILLER_0_64_1138 ();
 sg13g2_fill_8 FILLER_0_64_1146 ();
 sg13g2_fill_8 FILLER_0_64_1154 ();
 sg13g2_fill_8 FILLER_0_64_1162 ();
 sg13g2_fill_8 FILLER_0_64_1170 ();
 sg13g2_fill_8 FILLER_0_64_1178 ();
 sg13g2_fill_8 FILLER_0_64_1186 ();
 sg13g2_fill_8 FILLER_0_64_1194 ();
 sg13g2_fill_8 FILLER_0_64_1202 ();
 sg13g2_fill_8 FILLER_0_64_1210 ();
 sg13g2_fill_8 FILLER_0_64_1218 ();
 sg13g2_fill_2 FILLER_0_64_1226 ();
 sg13g2_fill_8 FILLER_0_65_0 ();
 sg13g2_fill_8 FILLER_0_65_8 ();
 sg13g2_fill_4 FILLER_0_65_16 ();
 sg13g2_fill_8 FILLER_0_65_30 ();
 sg13g2_fill_2 FILLER_0_65_38 ();
 sg13g2_fill_4 FILLER_0_65_44 ();
 sg13g2_fill_2 FILLER_0_65_48 ();
 sg13g2_fill_1 FILLER_0_65_147 ();
 sg13g2_fill_4 FILLER_0_65_158 ();
 sg13g2_fill_1 FILLER_0_65_172 ();
 sg13g2_fill_1 FILLER_0_65_183 ();
 sg13g2_fill_1 FILLER_0_65_199 ();
 sg13g2_fill_2 FILLER_0_65_226 ();
 sg13g2_fill_1 FILLER_0_65_292 ();
 sg13g2_fill_1 FILLER_0_65_319 ();
 sg13g2_fill_1 FILLER_0_65_346 ();
 sg13g2_fill_8 FILLER_0_65_365 ();
 sg13g2_fill_4 FILLER_0_65_373 ();
 sg13g2_fill_8 FILLER_0_65_403 ();
 sg13g2_fill_2 FILLER_0_65_411 ();
 sg13g2_fill_8 FILLER_0_65_441 ();
 sg13g2_fill_4 FILLER_0_65_449 ();
 sg13g2_fill_1 FILLER_0_65_453 ();
 sg13g2_fill_1 FILLER_0_65_480 ();
 sg13g2_fill_2 FILLER_0_65_491 ();
 sg13g2_fill_1 FILLER_0_65_493 ();
 sg13g2_fill_8 FILLER_0_65_502 ();
 sg13g2_fill_2 FILLER_0_65_510 ();
 sg13g2_fill_1 FILLER_0_65_512 ();
 sg13g2_fill_8 FILLER_0_65_528 ();
 sg13g2_fill_8 FILLER_0_65_536 ();
 sg13g2_fill_2 FILLER_0_65_544 ();
 sg13g2_fill_1 FILLER_0_65_546 ();
 sg13g2_fill_2 FILLER_0_65_660 ();
 sg13g2_fill_1 FILLER_0_65_662 ();
 sg13g2_fill_2 FILLER_0_65_699 ();
 sg13g2_decap_8 FILLER_0_65_710 ();
 sg13g2_fill_8 FILLER_0_65_721 ();
 sg13g2_fill_4 FILLER_0_65_729 ();
 sg13g2_fill_1 FILLER_0_65_737 ();
 sg13g2_fill_8 FILLER_0_65_774 ();
 sg13g2_fill_8 FILLER_0_65_786 ();
 sg13g2_fill_8 FILLER_0_65_794 ();
 sg13g2_fill_4 FILLER_0_65_802 ();
 sg13g2_fill_1 FILLER_0_65_806 ();
 sg13g2_fill_4 FILLER_0_65_811 ();
 sg13g2_fill_1 FILLER_0_65_815 ();
 sg13g2_fill_4 FILLER_0_65_857 ();
 sg13g2_fill_2 FILLER_0_65_861 ();
 sg13g2_fill_1 FILLER_0_65_881 ();
 sg13g2_fill_1 FILLER_0_65_892 ();
 sg13g2_fill_2 FILLER_0_65_903 ();
 sg13g2_fill_1 FILLER_0_65_931 ();
 sg13g2_fill_2 FILLER_0_65_942 ();
 sg13g2_fill_2 FILLER_0_65_948 ();
 sg13g2_fill_2 FILLER_0_65_960 ();
 sg13g2_fill_1 FILLER_0_65_962 ();
 sg13g2_fill_8 FILLER_0_65_984 ();
 sg13g2_fill_8 FILLER_0_65_992 ();
 sg13g2_fill_8 FILLER_0_65_1000 ();
 sg13g2_fill_8 FILLER_0_65_1008 ();
 sg13g2_fill_8 FILLER_0_65_1016 ();
 sg13g2_fill_8 FILLER_0_65_1024 ();
 sg13g2_fill_8 FILLER_0_65_1032 ();
 sg13g2_fill_8 FILLER_0_65_1040 ();
 sg13g2_fill_8 FILLER_0_65_1048 ();
 sg13g2_fill_8 FILLER_0_65_1056 ();
 sg13g2_fill_8 FILLER_0_65_1064 ();
 sg13g2_fill_8 FILLER_0_65_1072 ();
 sg13g2_fill_8 FILLER_0_65_1080 ();
 sg13g2_fill_8 FILLER_0_65_1088 ();
 sg13g2_fill_8 FILLER_0_65_1096 ();
 sg13g2_fill_8 FILLER_0_65_1104 ();
 sg13g2_fill_8 FILLER_0_65_1112 ();
 sg13g2_fill_8 FILLER_0_65_1120 ();
 sg13g2_fill_8 FILLER_0_65_1128 ();
 sg13g2_fill_8 FILLER_0_65_1136 ();
 sg13g2_fill_8 FILLER_0_65_1144 ();
 sg13g2_fill_8 FILLER_0_65_1152 ();
 sg13g2_fill_8 FILLER_0_65_1160 ();
 sg13g2_fill_8 FILLER_0_65_1168 ();
 sg13g2_fill_8 FILLER_0_65_1176 ();
 sg13g2_fill_8 FILLER_0_65_1184 ();
 sg13g2_fill_8 FILLER_0_65_1192 ();
 sg13g2_fill_8 FILLER_0_65_1200 ();
 sg13g2_fill_8 FILLER_0_65_1208 ();
 sg13g2_fill_8 FILLER_0_65_1216 ();
 sg13g2_fill_4 FILLER_0_65_1224 ();
 sg13g2_decap_8 FILLER_0_66_0 ();
 sg13g2_fill_2 FILLER_0_66_37 ();
 sg13g2_fill_2 FILLER_0_66_91 ();
 sg13g2_fill_1 FILLER_0_66_93 ();
 sg13g2_fill_4 FILLER_0_66_104 ();
 sg13g2_fill_2 FILLER_0_66_108 ();
 sg13g2_fill_1 FILLER_0_66_115 ();
 sg13g2_fill_2 FILLER_0_66_125 ();
 sg13g2_fill_1 FILLER_0_66_127 ();
 sg13g2_fill_4 FILLER_0_66_132 ();
 sg13g2_fill_2 FILLER_0_66_146 ();
 sg13g2_fill_2 FILLER_0_66_156 ();
 sg13g2_fill_8 FILLER_0_66_194 ();
 sg13g2_fill_2 FILLER_0_66_202 ();
 sg13g2_fill_2 FILLER_0_66_208 ();
 sg13g2_fill_1 FILLER_0_66_210 ();
 sg13g2_fill_8 FILLER_0_66_215 ();
 sg13g2_fill_8 FILLER_0_66_223 ();
 sg13g2_fill_2 FILLER_0_66_231 ();
 sg13g2_fill_1 FILLER_0_66_233 ();
 sg13g2_fill_2 FILLER_0_66_257 ();
 sg13g2_fill_1 FILLER_0_66_259 ();
 sg13g2_fill_1 FILLER_0_66_265 ();
 sg13g2_fill_2 FILLER_0_66_270 ();
 sg13g2_fill_1 FILLER_0_66_272 ();
 sg13g2_fill_4 FILLER_0_66_313 ();
 sg13g2_fill_1 FILLER_0_66_357 ();
 sg13g2_fill_2 FILLER_0_66_387 ();
 sg13g2_fill_2 FILLER_0_66_415 ();
 sg13g2_fill_1 FILLER_0_66_417 ();
 sg13g2_fill_2 FILLER_0_66_444 ();
 sg13g2_fill_1 FILLER_0_66_446 ();
 sg13g2_fill_4 FILLER_0_66_478 ();
 sg13g2_fill_2 FILLER_0_66_518 ();
 sg13g2_fill_4 FILLER_0_66_546 ();
 sg13g2_fill_1 FILLER_0_66_550 ();
 sg13g2_fill_1 FILLER_0_66_559 ();
 sg13g2_fill_1 FILLER_0_66_574 ();
 sg13g2_fill_1 FILLER_0_66_585 ();
 sg13g2_fill_1 FILLER_0_66_591 ();
 sg13g2_fill_1 FILLER_0_66_648 ();
 sg13g2_fill_8 FILLER_0_66_653 ();
 sg13g2_fill_8 FILLER_0_66_661 ();
 sg13g2_fill_4 FILLER_0_66_669 ();
 sg13g2_fill_1 FILLER_0_66_673 ();
 sg13g2_fill_2 FILLER_0_66_689 ();
 sg13g2_fill_1 FILLER_0_66_691 ();
 sg13g2_fill_1 FILLER_0_66_736 ();
 sg13g2_fill_1 FILLER_0_66_768 ();
 sg13g2_fill_1 FILLER_0_66_799 ();
 sg13g2_fill_2 FILLER_0_66_831 ();
 sg13g2_fill_2 FILLER_0_66_837 ();
 sg13g2_decap_8 FILLER_0_66_865 ();
 sg13g2_fill_8 FILLER_0_66_886 ();
 sg13g2_fill_4 FILLER_0_66_894 ();
 sg13g2_fill_1 FILLER_0_66_898 ();
 sg13g2_fill_4 FILLER_0_66_908 ();
 sg13g2_fill_2 FILLER_0_66_912 ();
 sg13g2_fill_8 FILLER_0_66_923 ();
 sg13g2_fill_4 FILLER_0_66_931 ();
 sg13g2_fill_1 FILLER_0_66_935 ();
 sg13g2_fill_8 FILLER_0_66_940 ();
 sg13g2_fill_4 FILLER_0_66_948 ();
 sg13g2_fill_2 FILLER_0_66_952 ();
 sg13g2_fill_8 FILLER_0_66_980 ();
 sg13g2_fill_8 FILLER_0_66_988 ();
 sg13g2_fill_8 FILLER_0_66_996 ();
 sg13g2_fill_8 FILLER_0_66_1004 ();
 sg13g2_fill_8 FILLER_0_66_1012 ();
 sg13g2_fill_8 FILLER_0_66_1020 ();
 sg13g2_fill_8 FILLER_0_66_1028 ();
 sg13g2_fill_8 FILLER_0_66_1036 ();
 sg13g2_fill_8 FILLER_0_66_1044 ();
 sg13g2_fill_8 FILLER_0_66_1052 ();
 sg13g2_fill_8 FILLER_0_66_1060 ();
 sg13g2_fill_8 FILLER_0_66_1068 ();
 sg13g2_fill_8 FILLER_0_66_1076 ();
 sg13g2_fill_8 FILLER_0_66_1084 ();
 sg13g2_fill_8 FILLER_0_66_1092 ();
 sg13g2_fill_8 FILLER_0_66_1100 ();
 sg13g2_fill_8 FILLER_0_66_1108 ();
 sg13g2_fill_8 FILLER_0_66_1116 ();
 sg13g2_fill_8 FILLER_0_66_1124 ();
 sg13g2_fill_8 FILLER_0_66_1132 ();
 sg13g2_fill_8 FILLER_0_66_1140 ();
 sg13g2_fill_8 FILLER_0_66_1148 ();
 sg13g2_fill_8 FILLER_0_66_1156 ();
 sg13g2_fill_8 FILLER_0_66_1164 ();
 sg13g2_fill_8 FILLER_0_66_1172 ();
 sg13g2_fill_8 FILLER_0_66_1180 ();
 sg13g2_fill_8 FILLER_0_66_1188 ();
 sg13g2_fill_8 FILLER_0_66_1196 ();
 sg13g2_fill_8 FILLER_0_66_1204 ();
 sg13g2_fill_8 FILLER_0_66_1212 ();
 sg13g2_fill_8 FILLER_0_66_1220 ();
 sg13g2_fill_1 FILLER_0_67_0 ();
 sg13g2_fill_2 FILLER_0_67_31 ();
 sg13g2_fill_2 FILLER_0_67_68 ();
 sg13g2_fill_1 FILLER_0_67_80 ();
 sg13g2_fill_2 FILLER_0_67_91 ();
 sg13g2_fill_8 FILLER_0_67_97 ();
 sg13g2_fill_8 FILLER_0_67_105 ();
 sg13g2_fill_8 FILLER_0_67_113 ();
 sg13g2_fill_1 FILLER_0_67_121 ();
 sg13g2_fill_4 FILLER_0_67_131 ();
 sg13g2_fill_1 FILLER_0_67_135 ();
 sg13g2_fill_4 FILLER_0_67_146 ();
 sg13g2_fill_1 FILLER_0_67_160 ();
 sg13g2_fill_8 FILLER_0_67_169 ();
 sg13g2_fill_8 FILLER_0_67_207 ();
 sg13g2_fill_8 FILLER_0_67_215 ();
 sg13g2_fill_8 FILLER_0_67_223 ();
 sg13g2_fill_8 FILLER_0_67_231 ();
 sg13g2_fill_1 FILLER_0_67_239 ();
 sg13g2_fill_8 FILLER_0_67_244 ();
 sg13g2_fill_8 FILLER_0_67_252 ();
 sg13g2_fill_8 FILLER_0_67_260 ();
 sg13g2_decap_8 FILLER_0_67_268 ();
 sg13g2_fill_8 FILLER_0_67_294 ();
 sg13g2_fill_8 FILLER_0_67_302 ();
 sg13g2_fill_2 FILLER_0_67_310 ();
 sg13g2_fill_1 FILLER_0_67_312 ();
 sg13g2_fill_2 FILLER_0_67_321 ();
 sg13g2_fill_1 FILLER_0_67_323 ();
 sg13g2_fill_1 FILLER_0_67_328 ();
 sg13g2_fill_1 FILLER_0_67_393 ();
 sg13g2_fill_2 FILLER_0_67_433 ();
 sg13g2_fill_8 FILLER_0_67_439 ();
 sg13g2_decap_8 FILLER_0_67_447 ();
 sg13g2_fill_4 FILLER_0_67_458 ();
 sg13g2_fill_1 FILLER_0_67_462 ();
 sg13g2_fill_2 FILLER_0_67_482 ();
 sg13g2_fill_4 FILLER_0_67_499 ();
 sg13g2_fill_8 FILLER_0_67_541 ();
 sg13g2_fill_1 FILLER_0_67_549 ();
 sg13g2_fill_2 FILLER_0_67_576 ();
 sg13g2_fill_8 FILLER_0_67_586 ();
 sg13g2_fill_2 FILLER_0_67_594 ();
 sg13g2_fill_2 FILLER_0_67_605 ();
 sg13g2_fill_8 FILLER_0_67_620 ();
 sg13g2_fill_8 FILLER_0_67_628 ();
 sg13g2_fill_8 FILLER_0_67_636 ();
 sg13g2_fill_8 FILLER_0_67_644 ();
 sg13g2_fill_8 FILLER_0_67_652 ();
 sg13g2_fill_4 FILLER_0_67_660 ();
 sg13g2_fill_8 FILLER_0_67_690 ();
 sg13g2_fill_4 FILLER_0_67_698 ();
 sg13g2_fill_1 FILLER_0_67_702 ();
 sg13g2_fill_2 FILLER_0_67_707 ();
 sg13g2_fill_1 FILLER_0_67_744 ();
 sg13g2_fill_8 FILLER_0_67_759 ();
 sg13g2_fill_2 FILLER_0_67_767 ();
 sg13g2_fill_8 FILLER_0_67_784 ();
 sg13g2_fill_1 FILLER_0_67_792 ();
 sg13g2_fill_1 FILLER_0_67_819 ();
 sg13g2_fill_2 FILLER_0_67_830 ();
 sg13g2_fill_1 FILLER_0_67_842 ();
 sg13g2_fill_2 FILLER_0_67_848 ();
 sg13g2_fill_8 FILLER_0_67_854 ();
 sg13g2_fill_8 FILLER_0_67_862 ();
 sg13g2_fill_4 FILLER_0_67_870 ();
 sg13g2_fill_1 FILLER_0_67_874 ();
 sg13g2_fill_4 FILLER_0_67_901 ();
 sg13g2_fill_2 FILLER_0_67_905 ();
 sg13g2_fill_8 FILLER_0_67_933 ();
 sg13g2_fill_2 FILLER_0_67_941 ();
 sg13g2_fill_2 FILLER_0_67_963 ();
 sg13g2_fill_1 FILLER_0_67_965 ();
 sg13g2_fill_4 FILLER_0_67_976 ();
 sg13g2_fill_1 FILLER_0_67_980 ();
 sg13g2_fill_2 FILLER_0_67_986 ();
 sg13g2_fill_1 FILLER_0_67_988 ();
 sg13g2_fill_2 FILLER_0_67_993 ();
 sg13g2_fill_8 FILLER_0_67_1000 ();
 sg13g2_fill_8 FILLER_0_67_1008 ();
 sg13g2_fill_8 FILLER_0_67_1016 ();
 sg13g2_fill_8 FILLER_0_67_1024 ();
 sg13g2_fill_8 FILLER_0_67_1032 ();
 sg13g2_fill_8 FILLER_0_67_1040 ();
 sg13g2_fill_8 FILLER_0_67_1048 ();
 sg13g2_fill_8 FILLER_0_67_1056 ();
 sg13g2_fill_8 FILLER_0_67_1064 ();
 sg13g2_fill_8 FILLER_0_67_1072 ();
 sg13g2_fill_8 FILLER_0_67_1080 ();
 sg13g2_fill_8 FILLER_0_67_1088 ();
 sg13g2_fill_8 FILLER_0_67_1096 ();
 sg13g2_fill_8 FILLER_0_67_1104 ();
 sg13g2_fill_8 FILLER_0_67_1112 ();
 sg13g2_fill_8 FILLER_0_67_1120 ();
 sg13g2_fill_8 FILLER_0_67_1128 ();
 sg13g2_fill_8 FILLER_0_67_1136 ();
 sg13g2_fill_8 FILLER_0_67_1144 ();
 sg13g2_fill_8 FILLER_0_67_1152 ();
 sg13g2_fill_8 FILLER_0_67_1160 ();
 sg13g2_fill_8 FILLER_0_67_1168 ();
 sg13g2_fill_8 FILLER_0_67_1176 ();
 sg13g2_fill_8 FILLER_0_67_1184 ();
 sg13g2_fill_8 FILLER_0_67_1192 ();
 sg13g2_fill_8 FILLER_0_67_1200 ();
 sg13g2_fill_8 FILLER_0_67_1208 ();
 sg13g2_fill_8 FILLER_0_67_1216 ();
 sg13g2_fill_4 FILLER_0_67_1224 ();
 sg13g2_fill_8 FILLER_0_68_0 ();
 sg13g2_fill_1 FILLER_0_68_18 ();
 sg13g2_fill_1 FILLER_0_68_29 ();
 sg13g2_fill_2 FILLER_0_68_48 ();
 sg13g2_fill_4 FILLER_0_68_65 ();
 sg13g2_fill_2 FILLER_0_68_69 ();
 sg13g2_fill_1 FILLER_0_68_84 ();
 sg13g2_decap_8 FILLER_0_68_111 ();
 sg13g2_fill_1 FILLER_0_68_149 ();
 sg13g2_fill_8 FILLER_0_68_176 ();
 sg13g2_fill_1 FILLER_0_68_184 ();
 sg13g2_fill_8 FILLER_0_68_200 ();
 sg13g2_fill_8 FILLER_0_68_208 ();
 sg13g2_fill_4 FILLER_0_68_216 ();
 sg13g2_fill_1 FILLER_0_68_220 ();
 sg13g2_fill_1 FILLER_0_68_251 ();
 sg13g2_fill_8 FILLER_0_68_281 ();
 sg13g2_fill_8 FILLER_0_68_289 ();
 sg13g2_fill_8 FILLER_0_68_327 ();
 sg13g2_fill_4 FILLER_0_68_340 ();
 sg13g2_fill_2 FILLER_0_68_344 ();
 sg13g2_fill_2 FILLER_0_68_354 ();
 sg13g2_fill_1 FILLER_0_68_368 ();
 sg13g2_fill_2 FILLER_0_68_377 ();
 sg13g2_fill_2 FILLER_0_68_383 ();
 sg13g2_fill_2 FILLER_0_68_411 ();
 sg13g2_fill_8 FILLER_0_68_439 ();
 sg13g2_fill_8 FILLER_0_68_447 ();
 sg13g2_fill_8 FILLER_0_68_455 ();
 sg13g2_decap_8 FILLER_0_68_463 ();
 sg13g2_fill_2 FILLER_0_68_480 ();
 sg13g2_fill_1 FILLER_0_68_482 ();
 sg13g2_fill_2 FILLER_0_68_519 ();
 sg13g2_fill_1 FILLER_0_68_521 ();
 sg13g2_fill_4 FILLER_0_68_548 ();
 sg13g2_fill_2 FILLER_0_68_552 ();
 sg13g2_fill_4 FILLER_0_68_559 ();
 sg13g2_fill_2 FILLER_0_68_563 ();
 sg13g2_fill_1 FILLER_0_68_575 ();
 sg13g2_fill_8 FILLER_0_68_581 ();
 sg13g2_fill_8 FILLER_0_68_604 ();
 sg13g2_fill_2 FILLER_0_68_612 ();
 sg13g2_fill_4 FILLER_0_68_622 ();
 sg13g2_fill_1 FILLER_0_68_640 ();
 sg13g2_fill_4 FILLER_0_68_667 ();
 sg13g2_fill_2 FILLER_0_68_671 ();
 sg13g2_fill_2 FILLER_0_68_677 ();
 sg13g2_fill_2 FILLER_0_68_684 ();
 sg13g2_fill_1 FILLER_0_68_686 ();
 sg13g2_fill_4 FILLER_0_68_706 ();
 sg13g2_fill_2 FILLER_0_68_715 ();
 sg13g2_fill_2 FILLER_0_68_721 ();
 sg13g2_decap_8 FILLER_0_68_733 ();
 sg13g2_fill_8 FILLER_0_68_748 ();
 sg13g2_fill_4 FILLER_0_68_764 ();
 sg13g2_fill_2 FILLER_0_68_799 ();
 sg13g2_fill_1 FILLER_0_68_801 ();
 sg13g2_fill_4 FILLER_0_68_806 ();
 sg13g2_fill_8 FILLER_0_68_833 ();
 sg13g2_fill_4 FILLER_0_68_841 ();
 sg13g2_fill_8 FILLER_0_68_855 ();
 sg13g2_fill_4 FILLER_0_68_863 ();
 sg13g2_fill_8 FILLER_0_68_901 ();
 sg13g2_fill_8 FILLER_0_68_909 ();
 sg13g2_fill_2 FILLER_0_68_917 ();
 sg13g2_fill_1 FILLER_0_68_919 ();
 sg13g2_fill_1 FILLER_0_68_946 ();
 sg13g2_fill_1 FILLER_0_68_952 ();
 sg13g2_fill_1 FILLER_0_68_979 ();
 sg13g2_fill_8 FILLER_0_68_1006 ();
 sg13g2_fill_8 FILLER_0_68_1014 ();
 sg13g2_fill_8 FILLER_0_68_1022 ();
 sg13g2_fill_8 FILLER_0_68_1030 ();
 sg13g2_fill_8 FILLER_0_68_1038 ();
 sg13g2_fill_8 FILLER_0_68_1046 ();
 sg13g2_fill_8 FILLER_0_68_1054 ();
 sg13g2_fill_8 FILLER_0_68_1062 ();
 sg13g2_fill_8 FILLER_0_68_1070 ();
 sg13g2_fill_8 FILLER_0_68_1078 ();
 sg13g2_fill_8 FILLER_0_68_1086 ();
 sg13g2_fill_8 FILLER_0_68_1094 ();
 sg13g2_fill_8 FILLER_0_68_1102 ();
 sg13g2_fill_8 FILLER_0_68_1110 ();
 sg13g2_fill_8 FILLER_0_68_1118 ();
 sg13g2_fill_8 FILLER_0_68_1126 ();
 sg13g2_fill_8 FILLER_0_68_1134 ();
 sg13g2_fill_8 FILLER_0_68_1142 ();
 sg13g2_fill_8 FILLER_0_68_1150 ();
 sg13g2_fill_8 FILLER_0_68_1158 ();
 sg13g2_fill_8 FILLER_0_68_1166 ();
 sg13g2_fill_8 FILLER_0_68_1174 ();
 sg13g2_fill_8 FILLER_0_68_1182 ();
 sg13g2_fill_8 FILLER_0_68_1190 ();
 sg13g2_fill_8 FILLER_0_68_1198 ();
 sg13g2_fill_8 FILLER_0_68_1206 ();
 sg13g2_fill_8 FILLER_0_68_1214 ();
 sg13g2_fill_4 FILLER_0_68_1222 ();
 sg13g2_fill_2 FILLER_0_68_1226 ();
 sg13g2_fill_1 FILLER_0_69_31 ();
 sg13g2_fill_8 FILLER_0_69_51 ();
 sg13g2_fill_2 FILLER_0_69_59 ();
 sg13g2_fill_1 FILLER_0_69_61 ();
 sg13g2_fill_4 FILLER_0_69_67 ();
 sg13g2_fill_1 FILLER_0_69_71 ();
 sg13g2_fill_1 FILLER_0_69_89 ();
 sg13g2_fill_2 FILLER_0_69_116 ();
 sg13g2_fill_2 FILLER_0_69_122 ();
 sg13g2_fill_4 FILLER_0_69_150 ();
 sg13g2_fill_2 FILLER_0_69_154 ();
 sg13g2_fill_8 FILLER_0_69_161 ();
 sg13g2_fill_4 FILLER_0_69_169 ();
 sg13g2_fill_2 FILLER_0_69_173 ();
 sg13g2_fill_8 FILLER_0_69_185 ();
 sg13g2_fill_1 FILLER_0_69_193 ();
 sg13g2_fill_2 FILLER_0_69_224 ();
 sg13g2_fill_2 FILLER_0_69_265 ();
 sg13g2_fill_1 FILLER_0_69_267 ();
 sg13g2_fill_8 FILLER_0_69_294 ();
 sg13g2_fill_2 FILLER_0_69_306 ();
 sg13g2_fill_4 FILLER_0_69_313 ();
 sg13g2_fill_2 FILLER_0_69_343 ();
 sg13g2_fill_4 FILLER_0_69_355 ();
 sg13g2_fill_4 FILLER_0_69_385 ();
 sg13g2_fill_2 FILLER_0_69_389 ();
 sg13g2_fill_2 FILLER_0_69_395 ();
 sg13g2_fill_1 FILLER_0_69_397 ();
 sg13g2_fill_4 FILLER_0_69_403 ();
 sg13g2_fill_1 FILLER_0_69_407 ();
 sg13g2_fill_1 FILLER_0_69_412 ();
 sg13g2_fill_8 FILLER_0_69_430 ();
 sg13g2_fill_4 FILLER_0_69_438 ();
 sg13g2_fill_2 FILLER_0_69_442 ();
 sg13g2_fill_4 FILLER_0_69_489 ();
 sg13g2_fill_2 FILLER_0_69_515 ();
 sg13g2_fill_8 FILLER_0_69_521 ();
 sg13g2_fill_1 FILLER_0_69_529 ();
 sg13g2_fill_2 FILLER_0_69_539 ();
 sg13g2_fill_1 FILLER_0_69_551 ();
 sg13g2_decap_8 FILLER_0_69_582 ();
 sg13g2_fill_8 FILLER_0_69_629 ();
 sg13g2_fill_1 FILLER_0_69_637 ();
 sg13g2_fill_4 FILLER_0_69_643 ();
 sg13g2_fill_8 FILLER_0_69_657 ();
 sg13g2_fill_2 FILLER_0_69_665 ();
 sg13g2_fill_2 FILLER_0_69_693 ();
 sg13g2_fill_1 FILLER_0_69_721 ();
 sg13g2_fill_1 FILLER_0_69_730 ();
 sg13g2_fill_1 FILLER_0_69_757 ();
 sg13g2_fill_1 FILLER_0_69_763 ();
 sg13g2_fill_2 FILLER_0_69_795 ();
 sg13g2_fill_4 FILLER_0_69_833 ();
 sg13g2_fill_2 FILLER_0_69_841 ();
 sg13g2_fill_8 FILLER_0_69_851 ();
 sg13g2_fill_8 FILLER_0_69_859 ();
 sg13g2_fill_1 FILLER_0_69_867 ();
 sg13g2_fill_2 FILLER_0_69_873 ();
 sg13g2_fill_4 FILLER_0_69_905 ();
 sg13g2_fill_1 FILLER_0_69_909 ();
 sg13g2_fill_1 FILLER_0_69_914 ();
 sg13g2_fill_4 FILLER_0_69_924 ();
 sg13g2_fill_1 FILLER_0_69_942 ();
 sg13g2_fill_1 FILLER_0_69_969 ();
 sg13g2_fill_1 FILLER_0_69_985 ();
 sg13g2_fill_1 FILLER_0_69_1022 ();
 sg13g2_fill_8 FILLER_0_69_1027 ();
 sg13g2_fill_8 FILLER_0_69_1035 ();
 sg13g2_fill_8 FILLER_0_69_1043 ();
 sg13g2_fill_8 FILLER_0_69_1051 ();
 sg13g2_fill_8 FILLER_0_69_1059 ();
 sg13g2_fill_8 FILLER_0_69_1067 ();
 sg13g2_fill_8 FILLER_0_69_1075 ();
 sg13g2_fill_8 FILLER_0_69_1083 ();
 sg13g2_fill_8 FILLER_0_69_1091 ();
 sg13g2_fill_8 FILLER_0_69_1099 ();
 sg13g2_fill_8 FILLER_0_69_1107 ();
 sg13g2_fill_8 FILLER_0_69_1115 ();
 sg13g2_fill_8 FILLER_0_69_1123 ();
 sg13g2_fill_8 FILLER_0_69_1131 ();
 sg13g2_fill_8 FILLER_0_69_1139 ();
 sg13g2_fill_8 FILLER_0_69_1147 ();
 sg13g2_fill_8 FILLER_0_69_1155 ();
 sg13g2_fill_8 FILLER_0_69_1163 ();
 sg13g2_fill_8 FILLER_0_69_1171 ();
 sg13g2_fill_8 FILLER_0_69_1179 ();
 sg13g2_fill_8 FILLER_0_69_1187 ();
 sg13g2_fill_8 FILLER_0_69_1195 ();
 sg13g2_fill_8 FILLER_0_69_1203 ();
 sg13g2_fill_8 FILLER_0_69_1211 ();
 sg13g2_fill_8 FILLER_0_69_1219 ();
 sg13g2_fill_1 FILLER_0_69_1227 ();
 sg13g2_fill_4 FILLER_0_70_0 ();
 sg13g2_fill_2 FILLER_0_70_4 ();
 sg13g2_fill_4 FILLER_0_70_10 ();
 sg13g2_fill_2 FILLER_0_70_14 ();
 sg13g2_fill_4 FILLER_0_70_42 ();
 sg13g2_fill_1 FILLER_0_70_64 ();
 sg13g2_fill_2 FILLER_0_70_105 ();
 sg13g2_fill_4 FILLER_0_70_144 ();
 sg13g2_fill_1 FILLER_0_70_148 ();
 sg13g2_fill_2 FILLER_0_70_179 ();
 sg13g2_fill_1 FILLER_0_70_181 ();
 sg13g2_fill_4 FILLER_0_70_213 ();
 sg13g2_fill_1 FILLER_0_70_217 ();
 sg13g2_fill_1 FILLER_0_70_244 ();
 sg13g2_fill_1 FILLER_0_70_259 ();
 sg13g2_decap_8 FILLER_0_70_286 ();
 sg13g2_fill_2 FILLER_0_70_297 ();
 sg13g2_fill_1 FILLER_0_70_303 ();
 sg13g2_fill_2 FILLER_0_70_314 ();
 sg13g2_fill_1 FILLER_0_70_321 ();
 sg13g2_fill_2 FILLER_0_70_332 ();
 sg13g2_fill_1 FILLER_0_70_360 ();
 sg13g2_fill_2 FILLER_0_70_366 ();
 sg13g2_fill_1 FILLER_0_70_378 ();
 sg13g2_fill_2 FILLER_0_70_384 ();
 sg13g2_fill_8 FILLER_0_70_390 ();
 sg13g2_fill_2 FILLER_0_70_398 ();
 sg13g2_fill_1 FILLER_0_70_400 ();
 sg13g2_fill_8 FILLER_0_70_427 ();
 sg13g2_fill_8 FILLER_0_70_435 ();
 sg13g2_fill_2 FILLER_0_70_443 ();
 sg13g2_fill_1 FILLER_0_70_445 ();
 sg13g2_fill_2 FILLER_0_70_472 ();
 sg13g2_fill_2 FILLER_0_70_483 ();
 sg13g2_fill_1 FILLER_0_70_516 ();
 sg13g2_fill_8 FILLER_0_70_522 ();
 sg13g2_fill_2 FILLER_0_70_530 ();
 sg13g2_fill_8 FILLER_0_70_536 ();
 sg13g2_fill_8 FILLER_0_70_544 ();
 sg13g2_fill_4 FILLER_0_70_552 ();
 sg13g2_fill_4 FILLER_0_70_590 ();
 sg13g2_fill_1 FILLER_0_70_594 ();
 sg13g2_fill_8 FILLER_0_70_599 ();
 sg13g2_fill_1 FILLER_0_70_673 ();
 sg13g2_fill_1 FILLER_0_70_678 ();
 sg13g2_fill_1 FILLER_0_70_689 ();
 sg13g2_fill_1 FILLER_0_70_698 ();
 sg13g2_fill_4 FILLER_0_70_725 ();
 sg13g2_fill_2 FILLER_0_70_729 ();
 sg13g2_fill_2 FILLER_0_70_740 ();
 sg13g2_fill_8 FILLER_0_70_808 ();
 sg13g2_fill_2 FILLER_0_70_816 ();
 sg13g2_fill_2 FILLER_0_70_885 ();
 sg13g2_fill_2 FILLER_0_70_897 ();
 sg13g2_fill_8 FILLER_0_70_903 ();
 sg13g2_fill_4 FILLER_0_70_911 ();
 sg13g2_fill_1 FILLER_0_70_915 ();
 sg13g2_fill_2 FILLER_0_70_925 ();
 sg13g2_fill_8 FILLER_0_70_937 ();
 sg13g2_fill_2 FILLER_0_70_945 ();
 sg13g2_fill_2 FILLER_0_70_956 ();
 sg13g2_fill_8 FILLER_0_70_966 ();
 sg13g2_fill_8 FILLER_0_70_974 ();
 sg13g2_fill_8 FILLER_0_70_982 ();
 sg13g2_fill_4 FILLER_0_70_990 ();
 sg13g2_fill_2 FILLER_0_70_1009 ();
 sg13g2_fill_8 FILLER_0_70_1015 ();
 sg13g2_fill_8 FILLER_0_70_1023 ();
 sg13g2_fill_8 FILLER_0_70_1031 ();
 sg13g2_fill_8 FILLER_0_70_1039 ();
 sg13g2_fill_8 FILLER_0_70_1047 ();
 sg13g2_fill_8 FILLER_0_70_1055 ();
 sg13g2_fill_8 FILLER_0_70_1063 ();
 sg13g2_fill_8 FILLER_0_70_1071 ();
 sg13g2_fill_8 FILLER_0_70_1079 ();
 sg13g2_fill_8 FILLER_0_70_1087 ();
 sg13g2_fill_8 FILLER_0_70_1095 ();
 sg13g2_fill_8 FILLER_0_70_1103 ();
 sg13g2_fill_8 FILLER_0_70_1111 ();
 sg13g2_fill_8 FILLER_0_70_1119 ();
 sg13g2_fill_8 FILLER_0_70_1127 ();
 sg13g2_fill_8 FILLER_0_70_1135 ();
 sg13g2_fill_8 FILLER_0_70_1143 ();
 sg13g2_fill_8 FILLER_0_70_1151 ();
 sg13g2_fill_8 FILLER_0_70_1159 ();
 sg13g2_fill_8 FILLER_0_70_1167 ();
 sg13g2_fill_8 FILLER_0_70_1175 ();
 sg13g2_fill_8 FILLER_0_70_1183 ();
 sg13g2_fill_8 FILLER_0_70_1191 ();
 sg13g2_fill_8 FILLER_0_70_1199 ();
 sg13g2_fill_8 FILLER_0_70_1207 ();
 sg13g2_fill_8 FILLER_0_70_1215 ();
 sg13g2_fill_4 FILLER_0_70_1223 ();
 sg13g2_fill_1 FILLER_0_70_1227 ();
 sg13g2_fill_8 FILLER_0_71_0 ();
 sg13g2_decap_8 FILLER_0_71_8 ();
 sg13g2_fill_1 FILLER_0_71_20 ();
 sg13g2_fill_1 FILLER_0_71_25 ();
 sg13g2_fill_4 FILLER_0_71_41 ();
 sg13g2_fill_1 FILLER_0_71_45 ();
 sg13g2_fill_4 FILLER_0_71_51 ();
 sg13g2_fill_1 FILLER_0_71_55 ();
 sg13g2_fill_1 FILLER_0_71_60 ();
 sg13g2_fill_4 FILLER_0_71_95 ();
 sg13g2_fill_1 FILLER_0_71_99 ();
 sg13g2_fill_1 FILLER_0_71_104 ();
 sg13g2_fill_1 FILLER_0_71_131 ();
 sg13g2_fill_1 FILLER_0_71_158 ();
 sg13g2_fill_1 FILLER_0_71_167 ();
 sg13g2_fill_1 FILLER_0_71_204 ();
 sg13g2_fill_8 FILLER_0_71_209 ();
 sg13g2_fill_8 FILLER_0_71_217 ();
 sg13g2_fill_8 FILLER_0_71_254 ();
 sg13g2_fill_8 FILLER_0_71_270 ();
 sg13g2_fill_8 FILLER_0_71_278 ();
 sg13g2_fill_4 FILLER_0_71_286 ();
 sg13g2_fill_2 FILLER_0_71_290 ();
 sg13g2_fill_1 FILLER_0_71_332 ();
 sg13g2_fill_8 FILLER_0_71_403 ();
 sg13g2_fill_8 FILLER_0_71_411 ();
 sg13g2_fill_2 FILLER_0_71_419 ();
 sg13g2_fill_1 FILLER_0_71_421 ();
 sg13g2_fill_8 FILLER_0_71_427 ();
 sg13g2_fill_8 FILLER_0_71_435 ();
 sg13g2_fill_8 FILLER_0_71_443 ();
 sg13g2_fill_1 FILLER_0_71_460 ();
 sg13g2_fill_1 FILLER_0_71_471 ();
 sg13g2_fill_1 FILLER_0_71_503 ();
 sg13g2_fill_1 FILLER_0_71_514 ();
 sg13g2_fill_1 FILLER_0_71_545 ();
 sg13g2_fill_2 FILLER_0_71_550 ();
 sg13g2_fill_8 FILLER_0_71_590 ();
 sg13g2_fill_2 FILLER_0_71_598 ();
 sg13g2_fill_1 FILLER_0_71_630 ();
 sg13g2_fill_8 FILLER_0_71_679 ();
 sg13g2_fill_2 FILLER_0_71_687 ();
 sg13g2_fill_2 FILLER_0_71_714 ();
 sg13g2_fill_2 FILLER_0_71_720 ();
 sg13g2_fill_2 FILLER_0_71_726 ();
 sg13g2_fill_2 FILLER_0_71_750 ();
 sg13g2_fill_8 FILLER_0_71_766 ();
 sg13g2_fill_8 FILLER_0_71_774 ();
 sg13g2_fill_4 FILLER_0_71_782 ();
 sg13g2_fill_1 FILLER_0_71_786 ();
 sg13g2_fill_8 FILLER_0_71_791 ();
 sg13g2_fill_8 FILLER_0_71_799 ();
 sg13g2_fill_4 FILLER_0_71_842 ();
 sg13g2_fill_8 FILLER_0_71_850 ();
 sg13g2_fill_2 FILLER_0_71_858 ();
 sg13g2_fill_2 FILLER_0_71_907 ();
 sg13g2_fill_1 FILLER_0_71_909 ();
 sg13g2_fill_2 FILLER_0_71_920 ();
 sg13g2_fill_1 FILLER_0_71_941 ();
 sg13g2_decap_8 FILLER_0_71_950 ();
 sg13g2_fill_8 FILLER_0_71_966 ();
 sg13g2_fill_8 FILLER_0_71_974 ();
 sg13g2_fill_2 FILLER_0_71_982 ();
 sg13g2_fill_4 FILLER_0_71_989 ();
 sg13g2_fill_1 FILLER_0_71_993 ();
 sg13g2_fill_8 FILLER_0_71_1030 ();
 sg13g2_fill_8 FILLER_0_71_1038 ();
 sg13g2_fill_8 FILLER_0_71_1046 ();
 sg13g2_fill_8 FILLER_0_71_1054 ();
 sg13g2_fill_8 FILLER_0_71_1062 ();
 sg13g2_fill_8 FILLER_0_71_1070 ();
 sg13g2_fill_8 FILLER_0_71_1078 ();
 sg13g2_fill_8 FILLER_0_71_1086 ();
 sg13g2_fill_8 FILLER_0_71_1094 ();
 sg13g2_fill_8 FILLER_0_71_1102 ();
 sg13g2_fill_8 FILLER_0_71_1110 ();
 sg13g2_fill_8 FILLER_0_71_1118 ();
 sg13g2_fill_8 FILLER_0_71_1126 ();
 sg13g2_fill_8 FILLER_0_71_1134 ();
 sg13g2_fill_8 FILLER_0_71_1142 ();
 sg13g2_fill_8 FILLER_0_71_1150 ();
 sg13g2_fill_8 FILLER_0_71_1158 ();
 sg13g2_fill_8 FILLER_0_71_1166 ();
 sg13g2_fill_8 FILLER_0_71_1174 ();
 sg13g2_fill_8 FILLER_0_71_1182 ();
 sg13g2_fill_8 FILLER_0_71_1190 ();
 sg13g2_fill_8 FILLER_0_71_1198 ();
 sg13g2_fill_8 FILLER_0_71_1206 ();
 sg13g2_fill_8 FILLER_0_71_1214 ();
 sg13g2_fill_4 FILLER_0_71_1222 ();
 sg13g2_fill_2 FILLER_0_71_1226 ();
 sg13g2_fill_2 FILLER_0_72_0 ();
 sg13g2_fill_1 FILLER_0_72_2 ();
 sg13g2_fill_2 FILLER_0_72_44 ();
 sg13g2_fill_1 FILLER_0_72_46 ();
 sg13g2_fill_8 FILLER_0_72_86 ();
 sg13g2_fill_4 FILLER_0_72_94 ();
 sg13g2_fill_8 FILLER_0_72_102 ();
 sg13g2_fill_8 FILLER_0_72_110 ();
 sg13g2_fill_1 FILLER_0_72_118 ();
 sg13g2_fill_4 FILLER_0_72_123 ();
 sg13g2_fill_2 FILLER_0_72_127 ();
 sg13g2_fill_2 FILLER_0_72_134 ();
 sg13g2_fill_1 FILLER_0_72_136 ();
 sg13g2_fill_2 FILLER_0_72_141 ();
 sg13g2_fill_1 FILLER_0_72_143 ();
 sg13g2_fill_2 FILLER_0_72_148 ();
 sg13g2_fill_1 FILLER_0_72_188 ();
 sg13g2_decap_8 FILLER_0_72_202 ();
 sg13g2_fill_4 FILLER_0_72_250 ();
 sg13g2_fill_1 FILLER_0_72_254 ();
 sg13g2_fill_8 FILLER_0_72_286 ();
 sg13g2_fill_2 FILLER_0_72_294 ();
 sg13g2_fill_1 FILLER_0_72_296 ();
 sg13g2_fill_8 FILLER_0_72_306 ();
 sg13g2_fill_8 FILLER_0_72_314 ();
 sg13g2_fill_2 FILLER_0_72_322 ();
 sg13g2_fill_4 FILLER_0_72_329 ();
 sg13g2_fill_2 FILLER_0_72_333 ();
 sg13g2_fill_2 FILLER_0_72_340 ();
 sg13g2_fill_8 FILLER_0_72_356 ();
 sg13g2_fill_2 FILLER_0_72_364 ();
 sg13g2_fill_1 FILLER_0_72_366 ();
 sg13g2_fill_4 FILLER_0_72_371 ();
 sg13g2_fill_8 FILLER_0_72_406 ();
 sg13g2_fill_8 FILLER_0_72_414 ();
 sg13g2_fill_8 FILLER_0_72_422 ();
 sg13g2_fill_8 FILLER_0_72_430 ();
 sg13g2_fill_8 FILLER_0_72_438 ();
 sg13g2_fill_1 FILLER_0_72_446 ();
 sg13g2_fill_2 FILLER_0_72_485 ();
 sg13g2_fill_1 FILLER_0_72_487 ();
 sg13g2_fill_1 FILLER_0_72_498 ();
 sg13g2_fill_8 FILLER_0_72_504 ();
 sg13g2_fill_1 FILLER_0_72_520 ();
 sg13g2_fill_1 FILLER_0_72_547 ();
 sg13g2_fill_8 FILLER_0_72_584 ();
 sg13g2_fill_4 FILLER_0_72_592 ();
 sg13g2_fill_1 FILLER_0_72_601 ();
 sg13g2_fill_1 FILLER_0_72_612 ();
 sg13g2_fill_1 FILLER_0_72_628 ();
 sg13g2_fill_2 FILLER_0_72_637 ();
 sg13g2_fill_1 FILLER_0_72_639 ();
 sg13g2_fill_4 FILLER_0_72_645 ();
 sg13g2_fill_1 FILLER_0_72_649 ();
 sg13g2_fill_8 FILLER_0_72_654 ();
 sg13g2_fill_8 FILLER_0_72_662 ();
 sg13g2_fill_8 FILLER_0_72_670 ();
 sg13g2_fill_4 FILLER_0_72_678 ();
 sg13g2_fill_1 FILLER_0_72_682 ();
 sg13g2_fill_2 FILLER_0_72_688 ();
 sg13g2_fill_1 FILLER_0_72_690 ();
 sg13g2_fill_8 FILLER_0_72_757 ();
 sg13g2_fill_8 FILLER_0_72_765 ();
 sg13g2_fill_1 FILLER_0_72_773 ();
 sg13g2_fill_1 FILLER_0_72_804 ();
 sg13g2_fill_1 FILLER_0_72_815 ();
 sg13g2_fill_1 FILLER_0_72_831 ();
 sg13g2_fill_8 FILLER_0_72_836 ();
 sg13g2_fill_8 FILLER_0_72_844 ();
 sg13g2_fill_8 FILLER_0_72_852 ();
 sg13g2_fill_8 FILLER_0_72_860 ();
 sg13g2_fill_2 FILLER_0_72_868 ();
 sg13g2_fill_1 FILLER_0_72_870 ();
 sg13g2_fill_4 FILLER_0_72_875 ();
 sg13g2_fill_1 FILLER_0_72_879 ();
 sg13g2_fill_4 FILLER_0_72_916 ();
 sg13g2_fill_2 FILLER_0_72_951 ();
 sg13g2_fill_4 FILLER_0_72_983 ();
 sg13g2_fill_8 FILLER_0_72_1021 ();
 sg13g2_fill_8 FILLER_0_72_1029 ();
 sg13g2_fill_8 FILLER_0_72_1037 ();
 sg13g2_fill_8 FILLER_0_72_1045 ();
 sg13g2_fill_8 FILLER_0_72_1053 ();
 sg13g2_fill_8 FILLER_0_72_1061 ();
 sg13g2_fill_8 FILLER_0_72_1069 ();
 sg13g2_fill_8 FILLER_0_72_1077 ();
 sg13g2_fill_8 FILLER_0_72_1085 ();
 sg13g2_fill_8 FILLER_0_72_1093 ();
 sg13g2_fill_8 FILLER_0_72_1101 ();
 sg13g2_fill_8 FILLER_0_72_1109 ();
 sg13g2_fill_8 FILLER_0_72_1117 ();
 sg13g2_fill_8 FILLER_0_72_1125 ();
 sg13g2_fill_8 FILLER_0_72_1133 ();
 sg13g2_fill_8 FILLER_0_72_1141 ();
 sg13g2_fill_8 FILLER_0_72_1149 ();
 sg13g2_fill_8 FILLER_0_72_1157 ();
 sg13g2_fill_8 FILLER_0_72_1165 ();
 sg13g2_fill_8 FILLER_0_72_1173 ();
 sg13g2_fill_8 FILLER_0_72_1181 ();
 sg13g2_fill_8 FILLER_0_72_1189 ();
 sg13g2_fill_8 FILLER_0_72_1197 ();
 sg13g2_fill_8 FILLER_0_72_1205 ();
 sg13g2_fill_8 FILLER_0_72_1213 ();
 sg13g2_decap_8 FILLER_0_72_1221 ();
 sg13g2_fill_8 FILLER_0_73_0 ();
 sg13g2_fill_2 FILLER_0_73_8 ();
 sg13g2_fill_1 FILLER_0_73_10 ();
 sg13g2_fill_1 FILLER_0_73_15 ();
 sg13g2_fill_1 FILLER_0_73_88 ();
 sg13g2_fill_2 FILLER_0_73_112 ();
 sg13g2_fill_1 FILLER_0_73_114 ();
 sg13g2_fill_4 FILLER_0_73_145 ();
 sg13g2_fill_1 FILLER_0_73_149 ();
 sg13g2_fill_2 FILLER_0_73_158 ();
 sg13g2_fill_1 FILLER_0_73_160 ();
 sg13g2_fill_4 FILLER_0_73_171 ();
 sg13g2_fill_2 FILLER_0_73_175 ();
 sg13g2_fill_4 FILLER_0_73_187 ();
 sg13g2_fill_2 FILLER_0_73_191 ();
 sg13g2_fill_4 FILLER_0_73_197 ();
 sg13g2_fill_1 FILLER_0_73_201 ();
 sg13g2_fill_8 FILLER_0_73_232 ();
 sg13g2_fill_8 FILLER_0_73_240 ();
 sg13g2_fill_2 FILLER_0_73_248 ();
 sg13g2_fill_2 FILLER_0_73_260 ();
 sg13g2_fill_1 FILLER_0_73_262 ();
 sg13g2_fill_8 FILLER_0_73_333 ();
 sg13g2_fill_8 FILLER_0_73_341 ();
 sg13g2_fill_2 FILLER_0_73_349 ();
 sg13g2_fill_8 FILLER_0_73_359 ();
 sg13g2_fill_1 FILLER_0_73_367 ();
 sg13g2_fill_4 FILLER_0_73_378 ();
 sg13g2_fill_2 FILLER_0_73_382 ();
 sg13g2_fill_2 FILLER_0_73_394 ();
 sg13g2_fill_1 FILLER_0_73_396 ();
 sg13g2_fill_2 FILLER_0_73_402 ();
 sg13g2_fill_1 FILLER_0_73_404 ();
 sg13g2_fill_8 FILLER_0_73_409 ();
 sg13g2_fill_8 FILLER_0_73_417 ();
 sg13g2_fill_8 FILLER_0_73_425 ();
 sg13g2_fill_8 FILLER_0_73_433 ();
 sg13g2_fill_4 FILLER_0_73_441 ();
 sg13g2_fill_1 FILLER_0_73_445 ();
 sg13g2_fill_2 FILLER_0_73_451 ();
 sg13g2_fill_2 FILLER_0_73_479 ();
 sg13g2_fill_2 FILLER_0_73_486 ();
 sg13g2_fill_1 FILLER_0_73_488 ();
 sg13g2_fill_1 FILLER_0_73_515 ();
 sg13g2_fill_4 FILLER_0_73_541 ();
 sg13g2_fill_2 FILLER_0_73_545 ();
 sg13g2_fill_2 FILLER_0_73_552 ();
 sg13g2_fill_2 FILLER_0_73_558 ();
 sg13g2_fill_2 FILLER_0_73_612 ();
 sg13g2_fill_1 FILLER_0_73_614 ();
 sg13g2_decap_8 FILLER_0_73_625 ();
 sg13g2_fill_4 FILLER_0_73_642 ();
 sg13g2_fill_1 FILLER_0_73_646 ();
 sg13g2_fill_8 FILLER_0_73_652 ();
 sg13g2_fill_8 FILLER_0_73_660 ();
 sg13g2_fill_8 FILLER_0_73_713 ();
 sg13g2_fill_2 FILLER_0_73_721 ();
 sg13g2_fill_1 FILLER_0_73_723 ();
 sg13g2_fill_8 FILLER_0_73_753 ();
 sg13g2_fill_8 FILLER_0_73_761 ();
 sg13g2_fill_4 FILLER_0_73_769 ();
 sg13g2_fill_2 FILLER_0_73_773 ();
 sg13g2_fill_4 FILLER_0_73_779 ();
 sg13g2_fill_1 FILLER_0_73_783 ();
 sg13g2_fill_1 FILLER_0_73_789 ();
 sg13g2_fill_2 FILLER_0_73_865 ();
 sg13g2_fill_8 FILLER_0_73_877 ();
 sg13g2_fill_8 FILLER_0_73_885 ();
 sg13g2_fill_2 FILLER_0_73_893 ();
 sg13g2_fill_2 FILLER_0_73_952 ();
 sg13g2_fill_4 FILLER_0_73_980 ();
 sg13g2_fill_8 FILLER_0_73_1015 ();
 sg13g2_fill_8 FILLER_0_73_1023 ();
 sg13g2_fill_8 FILLER_0_73_1031 ();
 sg13g2_fill_8 FILLER_0_73_1039 ();
 sg13g2_fill_8 FILLER_0_73_1047 ();
 sg13g2_fill_8 FILLER_0_73_1055 ();
 sg13g2_fill_8 FILLER_0_73_1063 ();
 sg13g2_fill_8 FILLER_0_73_1071 ();
 sg13g2_fill_8 FILLER_0_73_1079 ();
 sg13g2_fill_8 FILLER_0_73_1087 ();
 sg13g2_fill_8 FILLER_0_73_1095 ();
 sg13g2_fill_8 FILLER_0_73_1103 ();
 sg13g2_fill_8 FILLER_0_73_1111 ();
 sg13g2_fill_8 FILLER_0_73_1119 ();
 sg13g2_fill_8 FILLER_0_73_1127 ();
 sg13g2_fill_8 FILLER_0_73_1135 ();
 sg13g2_fill_8 FILLER_0_73_1143 ();
 sg13g2_fill_8 FILLER_0_73_1151 ();
 sg13g2_fill_8 FILLER_0_73_1159 ();
 sg13g2_fill_8 FILLER_0_73_1167 ();
 sg13g2_fill_8 FILLER_0_73_1175 ();
 sg13g2_fill_8 FILLER_0_73_1183 ();
 sg13g2_fill_8 FILLER_0_73_1191 ();
 sg13g2_fill_8 FILLER_0_73_1199 ();
 sg13g2_fill_8 FILLER_0_73_1207 ();
 sg13g2_fill_8 FILLER_0_73_1215 ();
 sg13g2_fill_4 FILLER_0_73_1223 ();
 sg13g2_fill_1 FILLER_0_73_1227 ();
 sg13g2_fill_2 FILLER_0_74_0 ();
 sg13g2_fill_1 FILLER_0_74_2 ();
 sg13g2_fill_1 FILLER_0_74_7 ();
 sg13g2_fill_4 FILLER_0_74_13 ();
 sg13g2_decap_8 FILLER_0_74_52 ();
 sg13g2_fill_2 FILLER_0_74_69 ();
 sg13g2_fill_1 FILLER_0_74_71 ();
 sg13g2_fill_1 FILLER_0_74_82 ();
 sg13g2_fill_2 FILLER_0_74_109 ();
 sg13g2_fill_1 FILLER_0_74_137 ();
 sg13g2_fill_4 FILLER_0_74_174 ();
 sg13g2_fill_1 FILLER_0_74_217 ();
 sg13g2_fill_8 FILLER_0_74_285 ();
 sg13g2_fill_1 FILLER_0_74_293 ();
 sg13g2_fill_4 FILLER_0_74_324 ();
 sg13g2_fill_4 FILLER_0_74_354 ();
 sg13g2_fill_2 FILLER_0_74_358 ();
 sg13g2_fill_4 FILLER_0_74_383 ();
 sg13g2_fill_1 FILLER_0_74_387 ();
 sg13g2_fill_8 FILLER_0_74_424 ();
 sg13g2_fill_8 FILLER_0_74_432 ();
 sg13g2_fill_8 FILLER_0_74_440 ();
 sg13g2_fill_4 FILLER_0_74_448 ();
 sg13g2_fill_4 FILLER_0_74_456 ();
 sg13g2_fill_8 FILLER_0_74_484 ();
 sg13g2_fill_2 FILLER_0_74_492 ();
 sg13g2_fill_1 FILLER_0_74_494 ();
 sg13g2_fill_8 FILLER_0_74_499 ();
 sg13g2_fill_8 FILLER_0_74_507 ();
 sg13g2_decap_8 FILLER_0_74_515 ();
 sg13g2_fill_8 FILLER_0_74_530 ();
 sg13g2_fill_8 FILLER_0_74_538 ();
 sg13g2_fill_8 FILLER_0_74_546 ();
 sg13g2_fill_8 FILLER_0_74_554 ();
 sg13g2_decap_8 FILLER_0_74_562 ();
 sg13g2_fill_4 FILLER_0_74_577 ();
 sg13g2_fill_4 FILLER_0_74_585 ();
 sg13g2_fill_2 FILLER_0_74_675 ();
 sg13g2_fill_4 FILLER_0_74_681 ();
 sg13g2_fill_4 FILLER_0_74_690 ();
 sg13g2_fill_8 FILLER_0_74_704 ();
 sg13g2_decap_8 FILLER_0_74_764 ();
 sg13g2_fill_2 FILLER_0_74_775 ();
 sg13g2_fill_1 FILLER_0_74_797 ();
 sg13g2_fill_2 FILLER_0_74_808 ();
 sg13g2_fill_1 FILLER_0_74_810 ();
 sg13g2_fill_2 FILLER_0_74_820 ();
 sg13g2_fill_1 FILLER_0_74_827 ();
 sg13g2_fill_1 FILLER_0_74_854 ();
 sg13g2_fill_2 FILLER_0_74_881 ();
 sg13g2_fill_1 FILLER_0_74_883 ();
 sg13g2_fill_8 FILLER_0_74_889 ();
 sg13g2_fill_8 FILLER_0_74_897 ();
 sg13g2_fill_4 FILLER_0_74_905 ();
 sg13g2_fill_1 FILLER_0_74_909 ();
 sg13g2_fill_8 FILLER_0_74_914 ();
 sg13g2_fill_1 FILLER_0_74_932 ();
 sg13g2_fill_8 FILLER_0_74_937 ();
 sg13g2_fill_1 FILLER_0_74_966 ();
 sg13g2_fill_1 FILLER_0_74_977 ();
 sg13g2_fill_1 FILLER_0_74_988 ();
 sg13g2_fill_2 FILLER_0_74_1003 ();
 sg13g2_fill_8 FILLER_0_74_1009 ();
 sg13g2_fill_8 FILLER_0_74_1017 ();
 sg13g2_fill_8 FILLER_0_74_1025 ();
 sg13g2_fill_8 FILLER_0_74_1033 ();
 sg13g2_fill_8 FILLER_0_74_1041 ();
 sg13g2_fill_8 FILLER_0_74_1049 ();
 sg13g2_fill_8 FILLER_0_74_1057 ();
 sg13g2_fill_8 FILLER_0_74_1065 ();
 sg13g2_fill_8 FILLER_0_74_1073 ();
 sg13g2_fill_8 FILLER_0_74_1081 ();
 sg13g2_fill_8 FILLER_0_74_1089 ();
 sg13g2_fill_8 FILLER_0_74_1097 ();
 sg13g2_fill_8 FILLER_0_74_1105 ();
 sg13g2_fill_8 FILLER_0_74_1113 ();
 sg13g2_fill_8 FILLER_0_74_1121 ();
 sg13g2_fill_8 FILLER_0_74_1129 ();
 sg13g2_fill_8 FILLER_0_74_1137 ();
 sg13g2_fill_8 FILLER_0_74_1145 ();
 sg13g2_fill_8 FILLER_0_74_1153 ();
 sg13g2_fill_8 FILLER_0_74_1161 ();
 sg13g2_fill_8 FILLER_0_74_1169 ();
 sg13g2_fill_8 FILLER_0_74_1177 ();
 sg13g2_fill_8 FILLER_0_74_1185 ();
 sg13g2_fill_8 FILLER_0_74_1193 ();
 sg13g2_fill_8 FILLER_0_74_1201 ();
 sg13g2_fill_8 FILLER_0_74_1209 ();
 sg13g2_fill_8 FILLER_0_74_1217 ();
 sg13g2_fill_2 FILLER_0_74_1225 ();
 sg13g2_fill_1 FILLER_0_74_1227 ();
 sg13g2_fill_1 FILLER_0_75_0 ();
 sg13g2_fill_8 FILLER_0_75_49 ();
 sg13g2_fill_1 FILLER_0_75_111 ();
 sg13g2_fill_8 FILLER_0_75_125 ();
 sg13g2_fill_4 FILLER_0_75_133 ();
 sg13g2_fill_2 FILLER_0_75_137 ();
 sg13g2_fill_1 FILLER_0_75_143 ();
 sg13g2_fill_4 FILLER_0_75_211 ();
 sg13g2_fill_1 FILLER_0_75_215 ();
 sg13g2_fill_2 FILLER_0_75_221 ();
 sg13g2_fill_1 FILLER_0_75_256 ();
 sg13g2_fill_4 FILLER_0_75_261 ();
 sg13g2_fill_4 FILLER_0_75_291 ();
 sg13g2_fill_2 FILLER_0_75_295 ();
 sg13g2_fill_1 FILLER_0_75_323 ();
 sg13g2_fill_2 FILLER_0_75_401 ();
 sg13g2_fill_8 FILLER_0_75_429 ();
 sg13g2_fill_8 FILLER_0_75_437 ();
 sg13g2_fill_8 FILLER_0_75_445 ();
 sg13g2_fill_8 FILLER_0_75_453 ();
 sg13g2_fill_8 FILLER_0_75_461 ();
 sg13g2_fill_8 FILLER_0_75_469 ();
 sg13g2_fill_8 FILLER_0_75_477 ();
 sg13g2_fill_1 FILLER_0_75_494 ();
 sg13g2_fill_8 FILLER_0_75_538 ();
 sg13g2_fill_1 FILLER_0_75_546 ();
 sg13g2_fill_2 FILLER_0_75_573 ();
 sg13g2_fill_1 FILLER_0_75_575 ();
 sg13g2_fill_8 FILLER_0_75_584 ();
 sg13g2_fill_4 FILLER_0_75_592 ();
 sg13g2_fill_1 FILLER_0_75_601 ();
 sg13g2_fill_2 FILLER_0_75_606 ();
 sg13g2_fill_1 FILLER_0_75_608 ();
 sg13g2_fill_2 FILLER_0_75_613 ();
 sg13g2_fill_1 FILLER_0_75_615 ();
 sg13g2_fill_1 FILLER_0_75_620 ();
 sg13g2_fill_2 FILLER_0_75_625 ();
 sg13g2_fill_1 FILLER_0_75_637 ();
 sg13g2_fill_4 FILLER_0_75_664 ();
 sg13g2_fill_2 FILLER_0_75_668 ();
 sg13g2_fill_1 FILLER_0_75_696 ();
 sg13g2_fill_1 FILLER_0_75_707 ();
 sg13g2_fill_8 FILLER_0_75_722 ();
 sg13g2_fill_1 FILLER_0_75_761 ();
 sg13g2_fill_8 FILLER_0_75_793 ();
 sg13g2_fill_8 FILLER_0_75_801 ();
 sg13g2_fill_8 FILLER_0_75_814 ();
 sg13g2_fill_4 FILLER_0_75_822 ();
 sg13g2_fill_1 FILLER_0_75_826 ();
 sg13g2_fill_4 FILLER_0_75_831 ();
 sg13g2_fill_1 FILLER_0_75_835 ();
 sg13g2_fill_8 FILLER_0_75_840 ();
 sg13g2_fill_2 FILLER_0_75_848 ();
 sg13g2_fill_1 FILLER_0_75_850 ();
 sg13g2_fill_1 FILLER_0_75_877 ();
 sg13g2_fill_1 FILLER_0_75_888 ();
 sg13g2_fill_1 FILLER_0_75_915 ();
 sg13g2_fill_1 FILLER_0_75_921 ();
 sg13g2_fill_1 FILLER_0_75_932 ();
 sg13g2_fill_8 FILLER_0_75_937 ();
 sg13g2_fill_8 FILLER_0_75_949 ();
 sg13g2_fill_2 FILLER_0_75_957 ();
 sg13g2_fill_1 FILLER_0_75_959 ();
 sg13g2_fill_4 FILLER_0_75_964 ();
 sg13g2_fill_8 FILLER_0_75_978 ();
 sg13g2_fill_8 FILLER_0_75_986 ();
 sg13g2_fill_8 FILLER_0_75_994 ();
 sg13g2_fill_8 FILLER_0_75_1002 ();
 sg13g2_fill_8 FILLER_0_75_1010 ();
 sg13g2_fill_8 FILLER_0_75_1018 ();
 sg13g2_fill_8 FILLER_0_75_1026 ();
 sg13g2_fill_8 FILLER_0_75_1034 ();
 sg13g2_fill_8 FILLER_0_75_1042 ();
 sg13g2_fill_8 FILLER_0_75_1050 ();
 sg13g2_fill_8 FILLER_0_75_1058 ();
 sg13g2_fill_8 FILLER_0_75_1066 ();
 sg13g2_fill_8 FILLER_0_75_1074 ();
 sg13g2_fill_8 FILLER_0_75_1082 ();
 sg13g2_fill_8 FILLER_0_75_1090 ();
 sg13g2_fill_8 FILLER_0_75_1098 ();
 sg13g2_fill_8 FILLER_0_75_1106 ();
 sg13g2_fill_8 FILLER_0_75_1114 ();
 sg13g2_fill_8 FILLER_0_75_1122 ();
 sg13g2_fill_8 FILLER_0_75_1130 ();
 sg13g2_fill_8 FILLER_0_75_1138 ();
 sg13g2_fill_8 FILLER_0_75_1146 ();
 sg13g2_fill_8 FILLER_0_75_1154 ();
 sg13g2_fill_8 FILLER_0_75_1162 ();
 sg13g2_fill_8 FILLER_0_75_1170 ();
 sg13g2_fill_8 FILLER_0_75_1178 ();
 sg13g2_fill_8 FILLER_0_75_1186 ();
 sg13g2_fill_8 FILLER_0_75_1194 ();
 sg13g2_fill_8 FILLER_0_75_1202 ();
 sg13g2_fill_8 FILLER_0_75_1210 ();
 sg13g2_fill_8 FILLER_0_75_1218 ();
 sg13g2_fill_2 FILLER_0_75_1226 ();
 sg13g2_fill_1 FILLER_0_76_0 ();
 sg13g2_fill_8 FILLER_0_76_42 ();
 sg13g2_fill_8 FILLER_0_76_50 ();
 sg13g2_decap_8 FILLER_0_76_58 ();
 sg13g2_fill_8 FILLER_0_76_73 ();
 sg13g2_fill_4 FILLER_0_76_81 ();
 sg13g2_fill_1 FILLER_0_76_85 ();
 sg13g2_fill_8 FILLER_0_76_94 ();
 sg13g2_fill_8 FILLER_0_76_102 ();
 sg13g2_fill_4 FILLER_0_76_110 ();
 sg13g2_decap_8 FILLER_0_76_129 ();
 sg13g2_fill_2 FILLER_0_76_173 ();
 sg13g2_fill_8 FILLER_0_76_209 ();
 sg13g2_fill_8 FILLER_0_76_217 ();
 sg13g2_fill_8 FILLER_0_76_225 ();
 sg13g2_fill_1 FILLER_0_76_233 ();
 sg13g2_fill_8 FILLER_0_76_238 ();
 sg13g2_fill_8 FILLER_0_76_246 ();
 sg13g2_fill_1 FILLER_0_76_254 ();
 sg13g2_fill_4 FILLER_0_76_259 ();
 sg13g2_fill_2 FILLER_0_76_268 ();
 sg13g2_fill_8 FILLER_0_76_278 ();
 sg13g2_fill_8 FILLER_0_76_286 ();
 sg13g2_fill_1 FILLER_0_76_294 ();
 sg13g2_fill_4 FILLER_0_76_300 ();
 sg13g2_fill_1 FILLER_0_76_304 ();
 sg13g2_fill_2 FILLER_0_76_314 ();
 sg13g2_fill_1 FILLER_0_76_331 ();
 sg13g2_fill_8 FILLER_0_76_351 ();
 sg13g2_decap_8 FILLER_0_76_359 ();
 sg13g2_fill_8 FILLER_0_76_370 ();
 sg13g2_fill_1 FILLER_0_76_378 ();
 sg13g2_fill_8 FILLER_0_76_414 ();
 sg13g2_fill_8 FILLER_0_76_422 ();
 sg13g2_fill_8 FILLER_0_76_430 ();
 sg13g2_fill_8 FILLER_0_76_438 ();
 sg13g2_fill_8 FILLER_0_76_446 ();
 sg13g2_fill_8 FILLER_0_76_454 ();
 sg13g2_fill_8 FILLER_0_76_462 ();
 sg13g2_fill_8 FILLER_0_76_470 ();
 sg13g2_fill_2 FILLER_0_76_478 ();
 sg13g2_fill_1 FILLER_0_76_506 ();
 sg13g2_fill_2 FILLER_0_76_511 ();
 sg13g2_fill_1 FILLER_0_76_539 ();
 sg13g2_fill_1 FILLER_0_76_544 ();
 sg13g2_fill_1 FILLER_0_76_591 ();
 sg13g2_fill_8 FILLER_0_76_596 ();
 sg13g2_fill_8 FILLER_0_76_604 ();
 sg13g2_fill_8 FILLER_0_76_612 ();
 sg13g2_decap_8 FILLER_0_76_620 ();
 sg13g2_fill_2 FILLER_0_76_631 ();
 sg13g2_fill_1 FILLER_0_76_633 ();
 sg13g2_fill_8 FILLER_0_76_658 ();
 sg13g2_fill_1 FILLER_0_76_666 ();
 sg13g2_fill_2 FILLER_0_76_675 ();
 sg13g2_fill_1 FILLER_0_76_677 ();
 sg13g2_fill_1 FILLER_0_76_704 ();
 sg13g2_fill_8 FILLER_0_76_715 ();
 sg13g2_fill_2 FILLER_0_76_723 ();
 sg13g2_fill_1 FILLER_0_76_725 ();
 sg13g2_decap_8 FILLER_0_76_736 ();
 sg13g2_fill_2 FILLER_0_76_747 ();
 sg13g2_fill_2 FILLER_0_76_753 ();
 sg13g2_fill_1 FILLER_0_76_755 ();
 sg13g2_fill_2 FILLER_0_76_782 ();
 sg13g2_fill_4 FILLER_0_76_789 ();
 sg13g2_fill_4 FILLER_0_76_819 ();
 sg13g2_fill_2 FILLER_0_76_842 ();
 sg13g2_fill_2 FILLER_0_76_853 ();
 sg13g2_fill_1 FILLER_0_76_855 ();
 sg13g2_fill_2 FILLER_0_76_865 ();
 sg13g2_fill_2 FILLER_0_76_877 ();
 sg13g2_fill_1 FILLER_0_76_879 ();
 sg13g2_fill_1 FILLER_0_76_890 ();
 sg13g2_fill_2 FILLER_0_76_917 ();
 sg13g2_fill_2 FILLER_0_76_945 ();
 sg13g2_fill_2 FILLER_0_76_959 ();
 sg13g2_fill_1 FILLER_0_76_961 ();
 sg13g2_fill_8 FILLER_0_76_1003 ();
 sg13g2_fill_8 FILLER_0_76_1011 ();
 sg13g2_fill_8 FILLER_0_76_1019 ();
 sg13g2_fill_8 FILLER_0_76_1027 ();
 sg13g2_fill_8 FILLER_0_76_1035 ();
 sg13g2_fill_8 FILLER_0_76_1043 ();
 sg13g2_fill_8 FILLER_0_76_1051 ();
 sg13g2_fill_8 FILLER_0_76_1059 ();
 sg13g2_fill_8 FILLER_0_76_1067 ();
 sg13g2_fill_8 FILLER_0_76_1075 ();
 sg13g2_fill_8 FILLER_0_76_1083 ();
 sg13g2_fill_8 FILLER_0_76_1091 ();
 sg13g2_fill_8 FILLER_0_76_1099 ();
 sg13g2_fill_8 FILLER_0_76_1107 ();
 sg13g2_fill_8 FILLER_0_76_1115 ();
 sg13g2_fill_8 FILLER_0_76_1123 ();
 sg13g2_fill_8 FILLER_0_76_1131 ();
 sg13g2_fill_8 FILLER_0_76_1139 ();
 sg13g2_fill_8 FILLER_0_76_1147 ();
 sg13g2_fill_8 FILLER_0_76_1155 ();
 sg13g2_fill_8 FILLER_0_76_1163 ();
 sg13g2_fill_8 FILLER_0_76_1171 ();
 sg13g2_fill_8 FILLER_0_76_1179 ();
 sg13g2_fill_8 FILLER_0_76_1187 ();
 sg13g2_fill_8 FILLER_0_76_1195 ();
 sg13g2_fill_8 FILLER_0_76_1203 ();
 sg13g2_fill_8 FILLER_0_76_1211 ();
 sg13g2_fill_8 FILLER_0_76_1219 ();
 sg13g2_fill_1 FILLER_0_76_1227 ();
 sg13g2_fill_8 FILLER_0_77_0 ();
 sg13g2_fill_2 FILLER_0_77_8 ();
 sg13g2_fill_2 FILLER_0_77_14 ();
 sg13g2_fill_8 FILLER_0_77_46 ();
 sg13g2_fill_8 FILLER_0_77_54 ();
 sg13g2_decap_8 FILLER_0_77_67 ();
 sg13g2_fill_8 FILLER_0_77_84 ();
 sg13g2_fill_8 FILLER_0_77_92 ();
 sg13g2_fill_8 FILLER_0_77_100 ();
 sg13g2_fill_2 FILLER_0_77_108 ();
 sg13g2_fill_2 FILLER_0_77_134 ();
 sg13g2_fill_8 FILLER_0_77_166 ();
 sg13g2_fill_8 FILLER_0_77_174 ();
 sg13g2_fill_1 FILLER_0_77_182 ();
 sg13g2_fill_8 FILLER_0_77_202 ();
 sg13g2_fill_8 FILLER_0_77_210 ();
 sg13g2_fill_8 FILLER_0_77_218 ();
 sg13g2_fill_8 FILLER_0_77_240 ();
 sg13g2_fill_1 FILLER_0_77_248 ();
 sg13g2_fill_2 FILLER_0_77_257 ();
 sg13g2_fill_1 FILLER_0_77_274 ();
 sg13g2_fill_8 FILLER_0_77_285 ();
 sg13g2_fill_8 FILLER_0_77_293 ();
 sg13g2_fill_4 FILLER_0_77_301 ();
 sg13g2_fill_1 FILLER_0_77_323 ();
 sg13g2_fill_8 FILLER_0_77_329 ();
 sg13g2_fill_4 FILLER_0_77_337 ();
 sg13g2_fill_8 FILLER_0_77_345 ();
 sg13g2_fill_8 FILLER_0_77_353 ();
 sg13g2_fill_1 FILLER_0_77_361 ();
 sg13g2_fill_4 FILLER_0_77_385 ();
 sg13g2_fill_1 FILLER_0_77_389 ();
 sg13g2_decap_8 FILLER_0_77_394 ();
 sg13g2_fill_8 FILLER_0_77_409 ();
 sg13g2_fill_4 FILLER_0_77_417 ();
 sg13g2_fill_1 FILLER_0_77_421 ();
 sg13g2_fill_4 FILLER_0_77_437 ();
 sg13g2_fill_8 FILLER_0_77_445 ();
 sg13g2_fill_4 FILLER_0_77_468 ();
 sg13g2_fill_2 FILLER_0_77_472 ();
 sg13g2_fill_1 FILLER_0_77_525 ();
 sg13g2_fill_1 FILLER_0_77_557 ();
 sg13g2_fill_2 FILLER_0_77_562 ();
 sg13g2_fill_2 FILLER_0_77_569 ();
 sg13g2_fill_2 FILLER_0_77_575 ();
 sg13g2_fill_1 FILLER_0_77_577 ();
 sg13g2_fill_2 FILLER_0_77_582 ();
 sg13g2_fill_2 FILLER_0_77_610 ();
 sg13g2_fill_1 FILLER_0_77_612 ();
 sg13g2_fill_2 FILLER_0_77_617 ();
 sg13g2_fill_1 FILLER_0_77_619 ();
 sg13g2_fill_1 FILLER_0_77_625 ();
 sg13g2_fill_2 FILLER_0_77_644 ();
 sg13g2_fill_1 FILLER_0_77_646 ();
 sg13g2_fill_2 FILLER_0_77_657 ();
 sg13g2_fill_8 FILLER_0_77_664 ();
 sg13g2_fill_2 FILLER_0_77_672 ();
 sg13g2_fill_8 FILLER_0_77_682 ();
 sg13g2_fill_8 FILLER_0_77_690 ();
 sg13g2_fill_2 FILLER_0_77_698 ();
 sg13g2_fill_8 FILLER_0_77_736 ();
 sg13g2_decap_8 FILLER_0_77_744 ();
 sg13g2_fill_2 FILLER_0_77_765 ();
 sg13g2_fill_1 FILLER_0_77_775 ();
 sg13g2_fill_1 FILLER_0_77_802 ();
 sg13g2_fill_2 FILLER_0_77_842 ();
 sg13g2_fill_1 FILLER_0_77_844 ();
 sg13g2_fill_2 FILLER_0_77_849 ();
 sg13g2_fill_2 FILLER_0_77_856 ();
 sg13g2_fill_1 FILLER_0_77_858 ();
 sg13g2_fill_4 FILLER_0_77_871 ();
 sg13g2_fill_2 FILLER_0_77_899 ();
 sg13g2_fill_8 FILLER_0_77_913 ();
 sg13g2_fill_8 FILLER_0_77_921 ();
 sg13g2_fill_4 FILLER_0_77_929 ();
 sg13g2_fill_8 FILLER_0_77_1020 ();
 sg13g2_fill_8 FILLER_0_77_1028 ();
 sg13g2_fill_8 FILLER_0_77_1036 ();
 sg13g2_fill_8 FILLER_0_77_1044 ();
 sg13g2_fill_8 FILLER_0_77_1052 ();
 sg13g2_fill_8 FILLER_0_77_1060 ();
 sg13g2_fill_8 FILLER_0_77_1068 ();
 sg13g2_fill_8 FILLER_0_77_1076 ();
 sg13g2_fill_8 FILLER_0_77_1084 ();
 sg13g2_fill_8 FILLER_0_77_1092 ();
 sg13g2_fill_8 FILLER_0_77_1100 ();
 sg13g2_fill_8 FILLER_0_77_1108 ();
 sg13g2_fill_8 FILLER_0_77_1116 ();
 sg13g2_fill_8 FILLER_0_77_1124 ();
 sg13g2_fill_8 FILLER_0_77_1132 ();
 sg13g2_fill_8 FILLER_0_77_1140 ();
 sg13g2_fill_8 FILLER_0_77_1148 ();
 sg13g2_fill_8 FILLER_0_77_1156 ();
 sg13g2_fill_8 FILLER_0_77_1164 ();
 sg13g2_fill_8 FILLER_0_77_1172 ();
 sg13g2_fill_8 FILLER_0_77_1180 ();
 sg13g2_fill_8 FILLER_0_77_1188 ();
 sg13g2_fill_8 FILLER_0_77_1196 ();
 sg13g2_fill_8 FILLER_0_77_1204 ();
 sg13g2_fill_8 FILLER_0_77_1212 ();
 sg13g2_fill_8 FILLER_0_77_1220 ();
 sg13g2_fill_8 FILLER_0_78_0 ();
 sg13g2_fill_8 FILLER_0_78_8 ();
 sg13g2_fill_4 FILLER_0_78_16 ();
 sg13g2_fill_2 FILLER_0_78_20 ();
 sg13g2_fill_8 FILLER_0_78_47 ();
 sg13g2_fill_4 FILLER_0_78_55 ();
 sg13g2_fill_1 FILLER_0_78_90 ();
 sg13g2_fill_4 FILLER_0_78_142 ();
 sg13g2_fill_1 FILLER_0_78_146 ();
 sg13g2_fill_4 FILLER_0_78_178 ();
 sg13g2_fill_2 FILLER_0_78_213 ();
 sg13g2_fill_8 FILLER_0_78_287 ();
 sg13g2_fill_2 FILLER_0_78_295 ();
 sg13g2_fill_1 FILLER_0_78_297 ();
 sg13g2_fill_4 FILLER_0_78_302 ();
 sg13g2_fill_2 FILLER_0_78_310 ();
 sg13g2_fill_1 FILLER_0_78_312 ();
 sg13g2_fill_2 FILLER_0_78_327 ();
 sg13g2_fill_2 FILLER_0_78_360 ();
 sg13g2_fill_1 FILLER_0_78_362 ();
 sg13g2_decap_8 FILLER_0_78_393 ();
 sg13g2_fill_1 FILLER_0_78_431 ();
 sg13g2_fill_2 FILLER_0_78_458 ();
 sg13g2_fill_1 FILLER_0_78_486 ();
 sg13g2_fill_1 FILLER_0_78_506 ();
 sg13g2_fill_1 FILLER_0_78_511 ();
 sg13g2_fill_2 FILLER_0_78_521 ();
 sg13g2_fill_2 FILLER_0_78_528 ();
 sg13g2_fill_2 FILLER_0_78_540 ();
 sg13g2_fill_2 FILLER_0_78_550 ();
 sg13g2_fill_1 FILLER_0_78_552 ();
 sg13g2_fill_8 FILLER_0_78_583 ();
 sg13g2_fill_1 FILLER_0_78_595 ();
 sg13g2_fill_2 FILLER_0_78_622 ();
 sg13g2_fill_2 FILLER_0_78_650 ();
 sg13g2_fill_1 FILLER_0_78_652 ();
 sg13g2_fill_8 FILLER_0_78_684 ();
 sg13g2_fill_8 FILLER_0_78_692 ();
 sg13g2_decap_8 FILLER_0_78_700 ();
 sg13g2_fill_4 FILLER_0_78_712 ();
 sg13g2_fill_1 FILLER_0_78_716 ();
 sg13g2_fill_8 FILLER_0_78_721 ();
 sg13g2_fill_8 FILLER_0_78_729 ();
 sg13g2_fill_4 FILLER_0_78_737 ();
 sg13g2_fill_2 FILLER_0_78_741 ();
 sg13g2_fill_1 FILLER_0_78_769 ();
 sg13g2_fill_1 FILLER_0_78_775 ();
 sg13g2_fill_1 FILLER_0_78_786 ();
 sg13g2_fill_1 FILLER_0_78_791 ();
 sg13g2_fill_1 FILLER_0_78_797 ();
 sg13g2_fill_2 FILLER_0_78_843 ();
 sg13g2_fill_1 FILLER_0_78_936 ();
 sg13g2_fill_2 FILLER_0_78_941 ();
 sg13g2_fill_1 FILLER_0_78_947 ();
 sg13g2_fill_2 FILLER_0_78_977 ();
 sg13g2_fill_1 FILLER_0_78_979 ();
 sg13g2_fill_2 FILLER_0_78_990 ();
 sg13g2_fill_2 FILLER_0_78_1002 ();
 sg13g2_fill_8 FILLER_0_78_1008 ();
 sg13g2_fill_8 FILLER_0_78_1016 ();
 sg13g2_fill_8 FILLER_0_78_1024 ();
 sg13g2_fill_8 FILLER_0_78_1032 ();
 sg13g2_fill_8 FILLER_0_78_1040 ();
 sg13g2_fill_8 FILLER_0_78_1048 ();
 sg13g2_fill_8 FILLER_0_78_1056 ();
 sg13g2_fill_8 FILLER_0_78_1064 ();
 sg13g2_fill_8 FILLER_0_78_1072 ();
 sg13g2_fill_8 FILLER_0_78_1080 ();
 sg13g2_fill_8 FILLER_0_78_1088 ();
 sg13g2_fill_8 FILLER_0_78_1096 ();
 sg13g2_fill_8 FILLER_0_78_1104 ();
 sg13g2_fill_8 FILLER_0_78_1112 ();
 sg13g2_fill_8 FILLER_0_78_1120 ();
 sg13g2_fill_8 FILLER_0_78_1128 ();
 sg13g2_fill_8 FILLER_0_78_1136 ();
 sg13g2_fill_8 FILLER_0_78_1144 ();
 sg13g2_fill_8 FILLER_0_78_1152 ();
 sg13g2_fill_8 FILLER_0_78_1160 ();
 sg13g2_fill_8 FILLER_0_78_1168 ();
 sg13g2_fill_8 FILLER_0_78_1176 ();
 sg13g2_fill_8 FILLER_0_78_1184 ();
 sg13g2_fill_8 FILLER_0_78_1192 ();
 sg13g2_fill_8 FILLER_0_78_1200 ();
 sg13g2_fill_8 FILLER_0_78_1208 ();
 sg13g2_fill_8 FILLER_0_78_1216 ();
 sg13g2_fill_4 FILLER_0_78_1224 ();
 sg13g2_fill_8 FILLER_0_79_0 ();
 sg13g2_fill_8 FILLER_0_79_8 ();
 sg13g2_fill_4 FILLER_0_79_16 ();
 sg13g2_fill_8 FILLER_0_79_87 ();
 sg13g2_fill_2 FILLER_0_79_95 ();
 sg13g2_fill_1 FILLER_0_79_97 ();
 sg13g2_fill_8 FILLER_0_79_141 ();
 sg13g2_fill_2 FILLER_0_79_149 ();
 sg13g2_fill_8 FILLER_0_79_165 ();
 sg13g2_fill_4 FILLER_0_79_173 ();
 sg13g2_fill_8 FILLER_0_79_192 ();
 sg13g2_fill_8 FILLER_0_79_200 ();
 sg13g2_fill_2 FILLER_0_79_208 ();
 sg13g2_fill_1 FILLER_0_79_210 ();
 sg13g2_fill_1 FILLER_0_79_252 ();
 sg13g2_fill_2 FILLER_0_79_315 ();
 sg13g2_fill_1 FILLER_0_79_317 ();
 sg13g2_fill_1 FILLER_0_79_328 ();
 sg13g2_fill_1 FILLER_0_79_355 ();
 sg13g2_fill_1 FILLER_0_79_370 ();
 sg13g2_fill_1 FILLER_0_79_376 ();
 sg13g2_fill_1 FILLER_0_79_403 ();
 sg13g2_fill_1 FILLER_0_79_430 ();
 sg13g2_fill_1 FILLER_0_79_467 ();
 sg13g2_fill_8 FILLER_0_79_472 ();
 sg13g2_fill_8 FILLER_0_79_480 ();
 sg13g2_fill_1 FILLER_0_79_488 ();
 sg13g2_fill_8 FILLER_0_79_509 ();
 sg13g2_fill_8 FILLER_0_79_517 ();
 sg13g2_fill_8 FILLER_0_79_525 ();
 sg13g2_fill_8 FILLER_0_79_533 ();
 sg13g2_fill_4 FILLER_0_79_541 ();
 sg13g2_fill_1 FILLER_0_79_553 ();
 sg13g2_fill_2 FILLER_0_79_580 ();
 sg13g2_fill_2 FILLER_0_79_590 ();
 sg13g2_fill_1 FILLER_0_79_592 ();
 sg13g2_fill_2 FILLER_0_79_611 ();
 sg13g2_fill_4 FILLER_0_79_618 ();
 sg13g2_fill_2 FILLER_0_79_658 ();
 sg13g2_fill_8 FILLER_0_79_690 ();
 sg13g2_fill_8 FILLER_0_79_698 ();
 sg13g2_fill_8 FILLER_0_79_706 ();
 sg13g2_fill_1 FILLER_0_79_714 ();
 sg13g2_fill_8 FILLER_0_79_723 ();
 sg13g2_fill_8 FILLER_0_79_731 ();
 sg13g2_fill_8 FILLER_0_79_739 ();
 sg13g2_fill_2 FILLER_0_79_747 ();
 sg13g2_fill_1 FILLER_0_79_749 ();
 sg13g2_fill_8 FILLER_0_79_754 ();
 sg13g2_fill_8 FILLER_0_79_762 ();
 sg13g2_fill_1 FILLER_0_79_770 ();
 sg13g2_fill_8 FILLER_0_79_776 ();
 sg13g2_fill_8 FILLER_0_79_784 ();
 sg13g2_fill_8 FILLER_0_79_792 ();
 sg13g2_fill_8 FILLER_0_79_804 ();
 sg13g2_decap_8 FILLER_0_79_812 ();
 sg13g2_fill_1 FILLER_0_79_859 ();
 sg13g2_fill_1 FILLER_0_79_886 ();
 sg13g2_fill_1 FILLER_0_79_891 ();
 sg13g2_fill_1 FILLER_0_79_896 ();
 sg13g2_fill_2 FILLER_0_79_954 ();
 sg13g2_fill_1 FILLER_0_79_956 ();
 sg13g2_fill_1 FILLER_0_79_1005 ();
 sg13g2_fill_8 FILLER_0_79_1010 ();
 sg13g2_fill_8 FILLER_0_79_1018 ();
 sg13g2_fill_8 FILLER_0_79_1026 ();
 sg13g2_fill_8 FILLER_0_79_1034 ();
 sg13g2_fill_8 FILLER_0_79_1042 ();
 sg13g2_fill_8 FILLER_0_79_1050 ();
 sg13g2_fill_8 FILLER_0_79_1058 ();
 sg13g2_fill_8 FILLER_0_79_1066 ();
 sg13g2_fill_8 FILLER_0_79_1074 ();
 sg13g2_fill_8 FILLER_0_79_1082 ();
 sg13g2_fill_8 FILLER_0_79_1090 ();
 sg13g2_fill_8 FILLER_0_79_1098 ();
 sg13g2_fill_8 FILLER_0_79_1106 ();
 sg13g2_fill_8 FILLER_0_79_1114 ();
 sg13g2_fill_8 FILLER_0_79_1122 ();
 sg13g2_fill_8 FILLER_0_79_1130 ();
 sg13g2_fill_8 FILLER_0_79_1138 ();
 sg13g2_fill_8 FILLER_0_79_1146 ();
 sg13g2_fill_8 FILLER_0_79_1154 ();
 sg13g2_fill_8 FILLER_0_79_1162 ();
 sg13g2_fill_8 FILLER_0_79_1170 ();
 sg13g2_fill_8 FILLER_0_79_1178 ();
 sg13g2_fill_8 FILLER_0_79_1186 ();
 sg13g2_fill_8 FILLER_0_79_1194 ();
 sg13g2_fill_8 FILLER_0_79_1202 ();
 sg13g2_fill_8 FILLER_0_79_1210 ();
 sg13g2_fill_8 FILLER_0_79_1218 ();
 sg13g2_fill_2 FILLER_0_79_1226 ();
 sg13g2_fill_8 FILLER_0_80_0 ();
 sg13g2_fill_8 FILLER_0_80_8 ();
 sg13g2_fill_8 FILLER_0_80_16 ();
 sg13g2_fill_4 FILLER_0_80_24 ();
 sg13g2_fill_2 FILLER_0_80_28 ();
 sg13g2_fill_1 FILLER_0_80_60 ();
 sg13g2_fill_2 FILLER_0_80_66 ();
 sg13g2_fill_2 FILLER_0_80_72 ();
 sg13g2_fill_8 FILLER_0_80_78 ();
 sg13g2_fill_4 FILLER_0_80_86 ();
 sg13g2_fill_8 FILLER_0_80_121 ();
 sg13g2_fill_8 FILLER_0_80_129 ();
 sg13g2_fill_8 FILLER_0_80_137 ();
 sg13g2_fill_8 FILLER_0_80_145 ();
 sg13g2_fill_8 FILLER_0_80_153 ();
 sg13g2_fill_1 FILLER_0_80_213 ();
 sg13g2_fill_1 FILLER_0_80_240 ();
 sg13g2_fill_4 FILLER_0_80_281 ();
 sg13g2_fill_1 FILLER_0_80_285 ();
 sg13g2_fill_4 FILLER_0_80_331 ();
 sg13g2_fill_1 FILLER_0_80_335 ();
 sg13g2_fill_1 FILLER_0_80_344 ();
 sg13g2_fill_1 FILLER_0_80_376 ();
 sg13g2_fill_1 FILLER_0_80_391 ();
 sg13g2_fill_2 FILLER_0_80_402 ();
 sg13g2_fill_2 FILLER_0_80_408 ();
 sg13g2_fill_1 FILLER_0_80_414 ();
 sg13g2_fill_1 FILLER_0_80_425 ();
 sg13g2_fill_1 FILLER_0_80_436 ();
 sg13g2_fill_4 FILLER_0_80_442 ();
 sg13g2_fill_8 FILLER_0_80_458 ();
 sg13g2_fill_8 FILLER_0_80_466 ();
 sg13g2_fill_2 FILLER_0_80_505 ();
 sg13g2_fill_4 FILLER_0_80_512 ();
 sg13g2_fill_2 FILLER_0_80_516 ();
 sg13g2_fill_4 FILLER_0_80_522 ();
 sg13g2_fill_2 FILLER_0_80_526 ();
 sg13g2_fill_1 FILLER_0_80_536 ();
 sg13g2_fill_1 FILLER_0_80_563 ();
 sg13g2_fill_1 FILLER_0_80_569 ();
 sg13g2_fill_1 FILLER_0_80_615 ();
 sg13g2_fill_2 FILLER_0_80_629 ();
 sg13g2_fill_1 FILLER_0_80_635 ();
 sg13g2_fill_2 FILLER_0_80_646 ();
 sg13g2_fill_1 FILLER_0_80_658 ();
 sg13g2_fill_8 FILLER_0_80_685 ();
 sg13g2_fill_8 FILLER_0_80_693 ();
 sg13g2_fill_8 FILLER_0_80_701 ();
 sg13g2_fill_8 FILLER_0_80_709 ();
 sg13g2_fill_8 FILLER_0_80_717 ();
 sg13g2_fill_8 FILLER_0_80_725 ();
 sg13g2_fill_8 FILLER_0_80_733 ();
 sg13g2_fill_8 FILLER_0_80_741 ();
 sg13g2_fill_8 FILLER_0_80_749 ();
 sg13g2_fill_8 FILLER_0_80_757 ();
 sg13g2_fill_8 FILLER_0_80_765 ();
 sg13g2_fill_4 FILLER_0_80_773 ();
 sg13g2_fill_2 FILLER_0_80_777 ();
 sg13g2_fill_1 FILLER_0_80_789 ();
 sg13g2_fill_8 FILLER_0_80_800 ();
 sg13g2_fill_8 FILLER_0_80_808 ();
 sg13g2_fill_8 FILLER_0_80_816 ();
 sg13g2_fill_2 FILLER_0_80_824 ();
 sg13g2_fill_1 FILLER_0_80_834 ();
 sg13g2_fill_1 FILLER_0_80_845 ();
 sg13g2_fill_1 FILLER_0_80_856 ();
 sg13g2_fill_2 FILLER_0_80_862 ();
 sg13g2_fill_1 FILLER_0_80_868 ();
 sg13g2_fill_1 FILLER_0_80_879 ();
 sg13g2_fill_1 FILLER_0_80_888 ();
 sg13g2_fill_1 FILLER_0_80_893 ();
 sg13g2_fill_1 FILLER_0_80_920 ();
 sg13g2_fill_2 FILLER_0_80_926 ();
 sg13g2_fill_2 FILLER_0_80_936 ();
 sg13g2_fill_2 FILLER_0_80_948 ();
 sg13g2_fill_1 FILLER_0_80_955 ();
 sg13g2_fill_2 FILLER_0_80_982 ();
 sg13g2_fill_1 FILLER_0_80_984 ();
 sg13g2_fill_4 FILLER_0_80_989 ();
 sg13g2_fill_1 FILLER_0_80_993 ();
 sg13g2_fill_8 FILLER_0_80_1020 ();
 sg13g2_fill_8 FILLER_0_80_1028 ();
 sg13g2_fill_8 FILLER_0_80_1036 ();
 sg13g2_fill_8 FILLER_0_80_1044 ();
 sg13g2_fill_8 FILLER_0_80_1052 ();
 sg13g2_fill_8 FILLER_0_80_1060 ();
 sg13g2_fill_8 FILLER_0_80_1068 ();
 sg13g2_fill_8 FILLER_0_80_1076 ();
 sg13g2_fill_8 FILLER_0_80_1084 ();
 sg13g2_fill_8 FILLER_0_80_1092 ();
 sg13g2_fill_8 FILLER_0_80_1100 ();
 sg13g2_fill_8 FILLER_0_80_1108 ();
 sg13g2_fill_8 FILLER_0_80_1116 ();
 sg13g2_fill_8 FILLER_0_80_1124 ();
 sg13g2_fill_8 FILLER_0_80_1132 ();
 sg13g2_fill_8 FILLER_0_80_1140 ();
 sg13g2_fill_8 FILLER_0_80_1148 ();
 sg13g2_fill_8 FILLER_0_80_1156 ();
 sg13g2_fill_8 FILLER_0_80_1164 ();
 sg13g2_fill_8 FILLER_0_80_1172 ();
 sg13g2_fill_8 FILLER_0_80_1180 ();
 sg13g2_fill_8 FILLER_0_80_1188 ();
 sg13g2_fill_8 FILLER_0_80_1196 ();
 sg13g2_fill_8 FILLER_0_80_1204 ();
 sg13g2_fill_8 FILLER_0_80_1212 ();
 sg13g2_fill_8 FILLER_0_80_1220 ();
 sg13g2_fill_8 FILLER_0_81_0 ();
 sg13g2_fill_8 FILLER_0_81_8 ();
 sg13g2_fill_8 FILLER_0_81_16 ();
 sg13g2_fill_8 FILLER_0_81_24 ();
 sg13g2_fill_2 FILLER_0_81_32 ();
 sg13g2_fill_2 FILLER_0_81_39 ();
 sg13g2_fill_8 FILLER_0_81_55 ();
 sg13g2_fill_8 FILLER_0_81_89 ();
 sg13g2_decap_8 FILLER_0_81_97 ();
 sg13g2_fill_8 FILLER_0_81_108 ();
 sg13g2_decap_8 FILLER_0_81_116 ();
 sg13g2_fill_8 FILLER_0_81_127 ();
 sg13g2_fill_1 FILLER_0_81_139 ();
 sg13g2_fill_2 FILLER_0_81_166 ();
 sg13g2_fill_1 FILLER_0_81_172 ();
 sg13g2_fill_1 FILLER_0_81_178 ();
 sg13g2_fill_1 FILLER_0_81_189 ();
 sg13g2_fill_8 FILLER_0_81_204 ();
 sg13g2_fill_4 FILLER_0_81_212 ();
 sg13g2_fill_2 FILLER_0_81_216 ();
 sg13g2_fill_1 FILLER_0_81_222 ();
 sg13g2_decap_8 FILLER_0_81_227 ();
 sg13g2_fill_1 FILLER_0_81_244 ();
 sg13g2_fill_2 FILLER_0_81_258 ();
 sg13g2_fill_1 FILLER_0_81_260 ();
 sg13g2_fill_2 FILLER_0_81_265 ();
 sg13g2_fill_1 FILLER_0_81_271 ();
 sg13g2_fill_1 FILLER_0_81_276 ();
 sg13g2_fill_1 FILLER_0_81_285 ();
 sg13g2_fill_1 FILLER_0_81_291 ();
 sg13g2_fill_4 FILLER_0_81_313 ();
 sg13g2_fill_8 FILLER_0_81_335 ();
 sg13g2_fill_8 FILLER_0_81_343 ();
 sg13g2_fill_1 FILLER_0_81_351 ();
 sg13g2_fill_4 FILLER_0_81_356 ();
 sg13g2_fill_2 FILLER_0_81_364 ();
 sg13g2_fill_2 FILLER_0_81_374 ();
 sg13g2_fill_1 FILLER_0_81_376 ();
 sg13g2_fill_4 FILLER_0_81_387 ();
 sg13g2_fill_2 FILLER_0_81_427 ();
 sg13g2_fill_1 FILLER_0_81_429 ();
 sg13g2_fill_8 FILLER_0_81_466 ();
 sg13g2_fill_8 FILLER_0_81_474 ();
 sg13g2_fill_1 FILLER_0_81_482 ();
 sg13g2_fill_2 FILLER_0_81_487 ();
 sg13g2_fill_2 FILLER_0_81_494 ();
 sg13g2_fill_1 FILLER_0_81_496 ();
 sg13g2_fill_1 FILLER_0_81_538 ();
 sg13g2_fill_2 FILLER_0_81_543 ();
 sg13g2_fill_2 FILLER_0_81_549 ();
 sg13g2_fill_2 FILLER_0_81_556 ();
 sg13g2_decap_8 FILLER_0_81_568 ();
 sg13g2_fill_2 FILLER_0_81_585 ();
 sg13g2_fill_8 FILLER_0_81_591 ();
 sg13g2_fill_8 FILLER_0_81_630 ();
 sg13g2_fill_8 FILLER_0_81_638 ();
 sg13g2_decap_8 FILLER_0_81_646 ();
 sg13g2_fill_4 FILLER_0_81_658 ();
 sg13g2_fill_2 FILLER_0_81_662 ();
 sg13g2_fill_4 FILLER_0_81_672 ();
 sg13g2_fill_1 FILLER_0_81_676 ();
 sg13g2_fill_8 FILLER_0_81_685 ();
 sg13g2_fill_8 FILLER_0_81_693 ();
 sg13g2_fill_8 FILLER_0_81_701 ();
 sg13g2_fill_8 FILLER_0_81_709 ();
 sg13g2_fill_8 FILLER_0_81_717 ();
 sg13g2_fill_8 FILLER_0_81_725 ();
 sg13g2_fill_4 FILLER_0_81_733 ();
 sg13g2_fill_4 FILLER_0_81_741 ();
 sg13g2_fill_1 FILLER_0_81_750 ();
 sg13g2_fill_1 FILLER_0_81_761 ();
 sg13g2_fill_2 FILLER_0_81_767 ();
 sg13g2_fill_2 FILLER_0_81_773 ();
 sg13g2_fill_1 FILLER_0_81_775 ();
 sg13g2_fill_1 FILLER_0_81_786 ();
 sg13g2_fill_2 FILLER_0_81_813 ();
 sg13g2_fill_1 FILLER_0_81_815 ();
 sg13g2_fill_4 FILLER_0_81_820 ();
 sg13g2_fill_1 FILLER_0_81_824 ();
 sg13g2_fill_8 FILLER_0_81_829 ();
 sg13g2_decap_8 FILLER_0_81_837 ();
 sg13g2_decap_8 FILLER_0_81_848 ();
 sg13g2_fill_8 FILLER_0_81_859 ();
 sg13g2_fill_8 FILLER_0_81_867 ();
 sg13g2_fill_8 FILLER_0_81_875 ();
 sg13g2_decap_8 FILLER_0_81_883 ();
 sg13g2_fill_2 FILLER_0_81_900 ();
 sg13g2_fill_2 FILLER_0_81_912 ();
 sg13g2_fill_4 FILLER_0_81_924 ();
 sg13g2_fill_1 FILLER_0_81_966 ();
 sg13g2_fill_8 FILLER_0_81_971 ();
 sg13g2_fill_8 FILLER_0_81_979 ();
 sg13g2_fill_2 FILLER_0_81_987 ();
 sg13g2_fill_1 FILLER_0_81_989 ();
 sg13g2_fill_8 FILLER_0_81_1015 ();
 sg13g2_fill_8 FILLER_0_81_1023 ();
 sg13g2_fill_8 FILLER_0_81_1031 ();
 sg13g2_fill_8 FILLER_0_81_1039 ();
 sg13g2_fill_8 FILLER_0_81_1047 ();
 sg13g2_fill_8 FILLER_0_81_1055 ();
 sg13g2_fill_8 FILLER_0_81_1063 ();
 sg13g2_fill_8 FILLER_0_81_1071 ();
 sg13g2_fill_8 FILLER_0_81_1079 ();
 sg13g2_fill_8 FILLER_0_81_1087 ();
 sg13g2_fill_8 FILLER_0_81_1095 ();
 sg13g2_fill_8 FILLER_0_81_1103 ();
 sg13g2_fill_8 FILLER_0_81_1111 ();
 sg13g2_fill_8 FILLER_0_81_1119 ();
 sg13g2_fill_8 FILLER_0_81_1127 ();
 sg13g2_fill_8 FILLER_0_81_1135 ();
 sg13g2_fill_8 FILLER_0_81_1143 ();
 sg13g2_fill_8 FILLER_0_81_1151 ();
 sg13g2_fill_8 FILLER_0_81_1159 ();
 sg13g2_fill_8 FILLER_0_81_1167 ();
 sg13g2_fill_8 FILLER_0_81_1175 ();
 sg13g2_fill_8 FILLER_0_81_1183 ();
 sg13g2_fill_8 FILLER_0_81_1191 ();
 sg13g2_fill_8 FILLER_0_81_1199 ();
 sg13g2_fill_8 FILLER_0_81_1207 ();
 sg13g2_fill_8 FILLER_0_81_1215 ();
 sg13g2_fill_4 FILLER_0_81_1223 ();
 sg13g2_fill_1 FILLER_0_81_1227 ();
 sg13g2_fill_8 FILLER_0_82_0 ();
 sg13g2_fill_8 FILLER_0_82_8 ();
 sg13g2_fill_8 FILLER_0_82_16 ();
 sg13g2_fill_8 FILLER_0_82_24 ();
 sg13g2_fill_4 FILLER_0_82_32 ();
 sg13g2_fill_1 FILLER_0_82_36 ();
 sg13g2_fill_8 FILLER_0_82_45 ();
 sg13g2_fill_8 FILLER_0_82_53 ();
 sg13g2_fill_8 FILLER_0_82_61 ();
 sg13g2_fill_1 FILLER_0_82_73 ();
 sg13g2_fill_8 FILLER_0_82_100 ();
 sg13g2_fill_2 FILLER_0_82_108 ();
 sg13g2_fill_8 FILLER_0_82_156 ();
 sg13g2_fill_4 FILLER_0_82_164 ();
 sg13g2_fill_2 FILLER_0_82_168 ();
 sg13g2_fill_2 FILLER_0_82_183 ();
 sg13g2_fill_1 FILLER_0_82_185 ();
 sg13g2_fill_8 FILLER_0_82_200 ();
 sg13g2_decap_8 FILLER_0_82_208 ();
 sg13g2_fill_2 FILLER_0_82_241 ();
 sg13g2_fill_1 FILLER_0_82_243 ();
 sg13g2_fill_8 FILLER_0_82_284 ();
 sg13g2_fill_1 FILLER_0_82_292 ();
 sg13g2_fill_8 FILLER_0_82_333 ();
 sg13g2_fill_8 FILLER_0_82_341 ();
 sg13g2_fill_8 FILLER_0_82_349 ();
 sg13g2_fill_2 FILLER_0_82_357 ();
 sg13g2_fill_2 FILLER_0_82_400 ();
 sg13g2_fill_1 FILLER_0_82_402 ();
 sg13g2_fill_8 FILLER_0_82_407 ();
 sg13g2_fill_4 FILLER_0_82_415 ();
 sg13g2_fill_2 FILLER_0_82_419 ();
 sg13g2_fill_2 FILLER_0_82_426 ();
 sg13g2_fill_4 FILLER_0_82_469 ();
 sg13g2_fill_1 FILLER_0_82_473 ();
 sg13g2_fill_2 FILLER_0_82_526 ();
 sg13g2_fill_1 FILLER_0_82_528 ();
 sg13g2_fill_2 FILLER_0_82_555 ();
 sg13g2_fill_2 FILLER_0_82_577 ();
 sg13g2_fill_1 FILLER_0_82_579 ();
 sg13g2_fill_8 FILLER_0_82_590 ();
 sg13g2_fill_8 FILLER_0_82_598 ();
 sg13g2_fill_8 FILLER_0_82_652 ();
 sg13g2_fill_2 FILLER_0_82_660 ();
 sg13g2_fill_8 FILLER_0_82_666 ();
 sg13g2_fill_8 FILLER_0_82_674 ();
 sg13g2_fill_8 FILLER_0_82_682 ();
 sg13g2_fill_8 FILLER_0_82_690 ();
 sg13g2_fill_8 FILLER_0_82_698 ();
 sg13g2_fill_8 FILLER_0_82_706 ();
 sg13g2_fill_8 FILLER_0_82_714 ();
 sg13g2_fill_8 FILLER_0_82_722 ();
 sg13g2_fill_1 FILLER_0_82_730 ();
 sg13g2_fill_8 FILLER_0_82_845 ();
 sg13g2_fill_8 FILLER_0_82_853 ();
 sg13g2_fill_8 FILLER_0_82_861 ();
 sg13g2_decap_8 FILLER_0_82_869 ();
 sg13g2_fill_8 FILLER_0_82_912 ();
 sg13g2_fill_2 FILLER_0_82_920 ();
 sg13g2_fill_1 FILLER_0_82_922 ();
 sg13g2_fill_4 FILLER_0_82_943 ();
 sg13g2_decap_8 FILLER_0_82_957 ();
 sg13g2_fill_8 FILLER_0_82_969 ();
 sg13g2_fill_8 FILLER_0_82_977 ();
 sg13g2_fill_1 FILLER_0_82_985 ();
 sg13g2_fill_8 FILLER_0_82_1029 ();
 sg13g2_fill_8 FILLER_0_82_1037 ();
 sg13g2_fill_8 FILLER_0_82_1045 ();
 sg13g2_fill_8 FILLER_0_82_1053 ();
 sg13g2_fill_8 FILLER_0_82_1061 ();
 sg13g2_fill_8 FILLER_0_82_1069 ();
 sg13g2_fill_8 FILLER_0_82_1077 ();
 sg13g2_fill_8 FILLER_0_82_1085 ();
 sg13g2_fill_8 FILLER_0_82_1093 ();
 sg13g2_fill_8 FILLER_0_82_1101 ();
 sg13g2_fill_8 FILLER_0_82_1109 ();
 sg13g2_fill_8 FILLER_0_82_1117 ();
 sg13g2_fill_8 FILLER_0_82_1125 ();
 sg13g2_fill_8 FILLER_0_82_1133 ();
 sg13g2_fill_8 FILLER_0_82_1141 ();
 sg13g2_fill_8 FILLER_0_82_1149 ();
 sg13g2_fill_8 FILLER_0_82_1157 ();
 sg13g2_fill_8 FILLER_0_82_1165 ();
 sg13g2_fill_8 FILLER_0_82_1173 ();
 sg13g2_fill_8 FILLER_0_82_1181 ();
 sg13g2_fill_8 FILLER_0_82_1189 ();
 sg13g2_fill_8 FILLER_0_82_1197 ();
 sg13g2_fill_8 FILLER_0_82_1205 ();
 sg13g2_fill_8 FILLER_0_82_1213 ();
 sg13g2_decap_8 FILLER_0_82_1221 ();
 sg13g2_fill_8 FILLER_0_83_0 ();
 sg13g2_decap_8 FILLER_0_83_8 ();
 sg13g2_fill_8 FILLER_0_83_19 ();
 sg13g2_fill_8 FILLER_0_83_58 ();
 sg13g2_fill_8 FILLER_0_83_66 ();
 sg13g2_fill_2 FILLER_0_83_74 ();
 sg13g2_fill_8 FILLER_0_83_147 ();
 sg13g2_fill_1 FILLER_0_83_155 ();
 sg13g2_fill_1 FILLER_0_83_170 ();
 sg13g2_fill_1 FILLER_0_83_181 ();
 sg13g2_fill_1 FILLER_0_83_192 ();
 sg13g2_fill_1 FILLER_0_83_219 ();
 sg13g2_fill_2 FILLER_0_83_246 ();
 sg13g2_fill_2 FILLER_0_83_266 ();
 sg13g2_fill_1 FILLER_0_83_268 ();
 sg13g2_fill_4 FILLER_0_83_295 ();
 sg13g2_fill_1 FILLER_0_83_299 ();
 sg13g2_fill_1 FILLER_0_83_339 ();
 sg13g2_fill_8 FILLER_0_83_344 ();
 sg13g2_fill_8 FILLER_0_83_352 ();
 sg13g2_fill_2 FILLER_0_83_360 ();
 sg13g2_fill_2 FILLER_0_83_410 ();
 sg13g2_fill_1 FILLER_0_83_427 ();
 sg13g2_fill_1 FILLER_0_83_436 ();
 sg13g2_fill_4 FILLER_0_83_477 ();
 sg13g2_fill_2 FILLER_0_83_481 ();
 sg13g2_fill_4 FILLER_0_83_487 ();
 sg13g2_fill_2 FILLER_0_83_491 ();
 sg13g2_fill_2 FILLER_0_83_526 ();
 sg13g2_fill_1 FILLER_0_83_528 ();
 sg13g2_decap_8 FILLER_0_83_539 ();
 sg13g2_fill_4 FILLER_0_83_572 ();
 sg13g2_fill_2 FILLER_0_83_599 ();
 sg13g2_fill_2 FILLER_0_83_611 ();
 sg13g2_fill_1 FILLER_0_83_613 ();
 sg13g2_fill_4 FILLER_0_83_644 ();
 sg13g2_fill_1 FILLER_0_83_648 ();
 sg13g2_fill_8 FILLER_0_83_680 ();
 sg13g2_fill_8 FILLER_0_83_688 ();
 sg13g2_fill_8 FILLER_0_83_696 ();
 sg13g2_fill_8 FILLER_0_83_704 ();
 sg13g2_fill_8 FILLER_0_83_712 ();
 sg13g2_fill_8 FILLER_0_83_720 ();
 sg13g2_fill_2 FILLER_0_83_808 ();
 sg13g2_fill_8 FILLER_0_83_872 ();
 sg13g2_fill_1 FILLER_0_83_880 ();
 sg13g2_fill_4 FILLER_0_83_915 ();
 sg13g2_fill_2 FILLER_0_83_919 ();
 sg13g2_fill_8 FILLER_0_83_1017 ();
 sg13g2_fill_8 FILLER_0_83_1025 ();
 sg13g2_fill_8 FILLER_0_83_1033 ();
 sg13g2_fill_8 FILLER_0_83_1041 ();
 sg13g2_fill_8 FILLER_0_83_1049 ();
 sg13g2_fill_8 FILLER_0_83_1057 ();
 sg13g2_fill_8 FILLER_0_83_1065 ();
 sg13g2_fill_8 FILLER_0_83_1073 ();
 sg13g2_fill_8 FILLER_0_83_1081 ();
 sg13g2_fill_8 FILLER_0_83_1089 ();
 sg13g2_fill_8 FILLER_0_83_1097 ();
 sg13g2_fill_8 FILLER_0_83_1105 ();
 sg13g2_fill_8 FILLER_0_83_1113 ();
 sg13g2_fill_8 FILLER_0_83_1121 ();
 sg13g2_fill_8 FILLER_0_83_1129 ();
 sg13g2_fill_8 FILLER_0_83_1137 ();
 sg13g2_fill_8 FILLER_0_83_1145 ();
 sg13g2_fill_8 FILLER_0_83_1153 ();
 sg13g2_fill_8 FILLER_0_83_1161 ();
 sg13g2_fill_8 FILLER_0_83_1169 ();
 sg13g2_fill_8 FILLER_0_83_1177 ();
 sg13g2_fill_8 FILLER_0_83_1185 ();
 sg13g2_fill_8 FILLER_0_83_1193 ();
 sg13g2_fill_8 FILLER_0_83_1201 ();
 sg13g2_fill_8 FILLER_0_83_1209 ();
 sg13g2_fill_8 FILLER_0_83_1217 ();
 sg13g2_fill_2 FILLER_0_83_1225 ();
 sg13g2_fill_1 FILLER_0_83_1227 ();
 sg13g2_fill_8 FILLER_0_84_0 ();
 sg13g2_fill_2 FILLER_0_84_34 ();
 sg13g2_fill_1 FILLER_0_84_36 ();
 sg13g2_fill_4 FILLER_0_84_68 ();
 sg13g2_fill_1 FILLER_0_84_72 ();
 sg13g2_fill_1 FILLER_0_84_102 ();
 sg13g2_fill_2 FILLER_0_84_117 ();
 sg13g2_fill_1 FILLER_0_84_119 ();
 sg13g2_fill_2 FILLER_0_84_130 ();
 sg13g2_fill_2 FILLER_0_84_142 ();
 sg13g2_fill_4 FILLER_0_84_180 ();
 sg13g2_fill_2 FILLER_0_84_223 ();
 sg13g2_fill_1 FILLER_0_84_225 ();
 sg13g2_fill_2 FILLER_0_84_230 ();
 sg13g2_fill_1 FILLER_0_84_232 ();
 sg13g2_fill_1 FILLER_0_84_259 ();
 sg13g2_fill_1 FILLER_0_84_296 ();
 sg13g2_fill_4 FILLER_0_84_359 ();
 sg13g2_fill_1 FILLER_0_84_363 ();
 sg13g2_fill_4 FILLER_0_84_402 ();
 sg13g2_fill_4 FILLER_0_84_432 ();
 sg13g2_fill_8 FILLER_0_84_513 ();
 sg13g2_fill_8 FILLER_0_84_521 ();
 sg13g2_fill_8 FILLER_0_84_529 ();
 sg13g2_fill_8 FILLER_0_84_537 ();
 sg13g2_fill_2 FILLER_0_84_545 ();
 sg13g2_fill_1 FILLER_0_84_547 ();
 sg13g2_fill_4 FILLER_0_84_613 ();
 sg13g2_fill_1 FILLER_0_84_617 ();
 sg13g2_fill_1 FILLER_0_84_628 ();
 sg13g2_fill_8 FILLER_0_84_639 ();
 sg13g2_fill_8 FILLER_0_84_647 ();
 sg13g2_fill_8 FILLER_0_84_655 ();
 sg13g2_fill_8 FILLER_0_84_663 ();
 sg13g2_fill_8 FILLER_0_84_671 ();
 sg13g2_fill_8 FILLER_0_84_679 ();
 sg13g2_fill_8 FILLER_0_84_687 ();
 sg13g2_fill_8 FILLER_0_84_695 ();
 sg13g2_fill_8 FILLER_0_84_703 ();
 sg13g2_fill_8 FILLER_0_84_711 ();
 sg13g2_fill_8 FILLER_0_84_719 ();
 sg13g2_decap_8 FILLER_0_84_727 ();
 sg13g2_fill_8 FILLER_0_84_738 ();
 sg13g2_fill_4 FILLER_0_84_746 ();
 sg13g2_fill_1 FILLER_0_84_765 ();
 sg13g2_fill_8 FILLER_0_84_771 ();
 sg13g2_fill_8 FILLER_0_84_793 ();
 sg13g2_fill_8 FILLER_0_84_801 ();
 sg13g2_fill_2 FILLER_0_84_809 ();
 sg13g2_fill_2 FILLER_0_84_816 ();
 sg13g2_fill_1 FILLER_0_84_818 ();
 sg13g2_fill_2 FILLER_0_84_824 ();
 sg13g2_fill_1 FILLER_0_84_826 ();
 sg13g2_fill_1 FILLER_0_84_837 ();
 sg13g2_fill_4 FILLER_0_84_868 ();
 sg13g2_fill_1 FILLER_0_84_890 ();
 sg13g2_fill_1 FILLER_0_84_896 ();
 sg13g2_fill_2 FILLER_0_84_901 ();
 sg13g2_fill_2 FILLER_0_84_913 ();
 sg13g2_fill_2 FILLER_0_84_919 ();
 sg13g2_fill_1 FILLER_0_84_921 ();
 sg13g2_fill_8 FILLER_0_84_948 ();
 sg13g2_fill_2 FILLER_0_84_956 ();
 sg13g2_fill_1 FILLER_0_84_993 ();
 sg13g2_fill_8 FILLER_0_84_1020 ();
 sg13g2_fill_8 FILLER_0_84_1028 ();
 sg13g2_fill_8 FILLER_0_84_1036 ();
 sg13g2_fill_8 FILLER_0_84_1044 ();
 sg13g2_fill_8 FILLER_0_84_1052 ();
 sg13g2_fill_8 FILLER_0_84_1060 ();
 sg13g2_fill_8 FILLER_0_84_1068 ();
 sg13g2_fill_8 FILLER_0_84_1076 ();
 sg13g2_fill_8 FILLER_0_84_1084 ();
 sg13g2_fill_8 FILLER_0_84_1092 ();
 sg13g2_fill_8 FILLER_0_84_1100 ();
 sg13g2_fill_8 FILLER_0_84_1108 ();
 sg13g2_fill_8 FILLER_0_84_1116 ();
 sg13g2_fill_8 FILLER_0_84_1124 ();
 sg13g2_fill_8 FILLER_0_84_1132 ();
 sg13g2_fill_8 FILLER_0_84_1140 ();
 sg13g2_fill_8 FILLER_0_84_1148 ();
 sg13g2_fill_8 FILLER_0_84_1156 ();
 sg13g2_fill_8 FILLER_0_84_1164 ();
 sg13g2_fill_8 FILLER_0_84_1172 ();
 sg13g2_fill_8 FILLER_0_84_1180 ();
 sg13g2_fill_8 FILLER_0_84_1188 ();
 sg13g2_fill_8 FILLER_0_84_1196 ();
 sg13g2_fill_8 FILLER_0_84_1204 ();
 sg13g2_fill_8 FILLER_0_84_1212 ();
 sg13g2_fill_8 FILLER_0_84_1220 ();
 sg13g2_fill_4 FILLER_0_85_0 ();
 sg13g2_fill_2 FILLER_0_85_13 ();
 sg13g2_fill_1 FILLER_0_85_30 ();
 sg13g2_fill_1 FILLER_0_85_49 ();
 sg13g2_fill_2 FILLER_0_85_76 ();
 sg13g2_fill_4 FILLER_0_85_198 ();
 sg13g2_fill_1 FILLER_0_85_202 ();
 sg13g2_fill_8 FILLER_0_85_211 ();
 sg13g2_fill_2 FILLER_0_85_219 ();
 sg13g2_fill_1 FILLER_0_85_240 ();
 sg13g2_fill_2 FILLER_0_85_245 ();
 sg13g2_fill_1 FILLER_0_85_247 ();
 sg13g2_fill_2 FILLER_0_85_258 ();
 sg13g2_fill_1 FILLER_0_85_260 ();
 sg13g2_fill_8 FILLER_0_85_289 ();
 sg13g2_decap_8 FILLER_0_85_297 ();
 sg13g2_fill_8 FILLER_0_85_338 ();
 sg13g2_fill_4 FILLER_0_85_346 ();
 sg13g2_fill_8 FILLER_0_85_354 ();
 sg13g2_fill_8 FILLER_0_85_362 ();
 sg13g2_fill_1 FILLER_0_85_370 ();
 sg13g2_fill_8 FILLER_0_85_389 ();
 sg13g2_fill_8 FILLER_0_85_397 ();
 sg13g2_fill_4 FILLER_0_85_405 ();
 sg13g2_fill_2 FILLER_0_85_409 ();
 sg13g2_fill_8 FILLER_0_85_415 ();
 sg13g2_fill_8 FILLER_0_85_423 ();
 sg13g2_fill_8 FILLER_0_85_431 ();
 sg13g2_fill_4 FILLER_0_85_439 ();
 sg13g2_fill_2 FILLER_0_85_443 ();
 sg13g2_fill_2 FILLER_0_85_450 ();
 sg13g2_fill_4 FILLER_0_85_479 ();
 sg13g2_fill_1 FILLER_0_85_487 ();
 sg13g2_fill_2 FILLER_0_85_493 ();
 sg13g2_fill_2 FILLER_0_85_505 ();
 sg13g2_fill_2 FILLER_0_85_533 ();
 sg13g2_fill_8 FILLER_0_85_539 ();
 sg13g2_fill_8 FILLER_0_85_547 ();
 sg13g2_fill_8 FILLER_0_85_555 ();
 sg13g2_fill_1 FILLER_0_85_563 ();
 sg13g2_fill_8 FILLER_0_85_568 ();
 sg13g2_fill_8 FILLER_0_85_606 ();
 sg13g2_fill_8 FILLER_0_85_614 ();
 sg13g2_fill_1 FILLER_0_85_622 ();
 sg13g2_fill_8 FILLER_0_85_627 ();
 sg13g2_fill_2 FILLER_0_85_635 ();
 sg13g2_fill_8 FILLER_0_85_647 ();
 sg13g2_fill_8 FILLER_0_85_655 ();
 sg13g2_fill_4 FILLER_0_85_663 ();
 sg13g2_fill_1 FILLER_0_85_667 ();
 sg13g2_fill_8 FILLER_0_85_682 ();
 sg13g2_fill_8 FILLER_0_85_690 ();
 sg13g2_fill_4 FILLER_0_85_698 ();
 sg13g2_fill_1 FILLER_0_85_702 ();
 sg13g2_fill_8 FILLER_0_85_707 ();
 sg13g2_fill_8 FILLER_0_85_715 ();
 sg13g2_fill_1 FILLER_0_85_723 ();
 sg13g2_fill_8 FILLER_0_85_767 ();
 sg13g2_fill_8 FILLER_0_85_775 ();
 sg13g2_fill_8 FILLER_0_85_783 ();
 sg13g2_fill_8 FILLER_0_85_791 ();
 sg13g2_fill_1 FILLER_0_85_799 ();
 sg13g2_fill_4 FILLER_0_85_813 ();
 sg13g2_fill_2 FILLER_0_85_851 ();
 sg13g2_fill_1 FILLER_0_85_905 ();
 sg13g2_fill_8 FILLER_0_85_911 ();
 sg13g2_fill_4 FILLER_0_85_919 ();
 sg13g2_fill_4 FILLER_0_85_928 ();
 sg13g2_fill_1 FILLER_0_85_932 ();
 sg13g2_fill_1 FILLER_0_85_951 ();
 sg13g2_fill_2 FILLER_0_85_983 ();
 sg13g2_fill_1 FILLER_0_85_989 ();
 sg13g2_fill_2 FILLER_0_85_994 ();
 sg13g2_fill_1 FILLER_0_85_996 ();
 sg13g2_fill_2 FILLER_0_85_1002 ();
 sg13g2_fill_1 FILLER_0_85_1004 ();
 sg13g2_fill_8 FILLER_0_85_1009 ();
 sg13g2_fill_8 FILLER_0_85_1017 ();
 sg13g2_fill_8 FILLER_0_85_1025 ();
 sg13g2_fill_8 FILLER_0_85_1033 ();
 sg13g2_fill_8 FILLER_0_85_1041 ();
 sg13g2_fill_8 FILLER_0_85_1049 ();
 sg13g2_fill_8 FILLER_0_85_1057 ();
 sg13g2_fill_8 FILLER_0_85_1065 ();
 sg13g2_fill_8 FILLER_0_85_1073 ();
 sg13g2_fill_8 FILLER_0_85_1081 ();
 sg13g2_fill_8 FILLER_0_85_1089 ();
 sg13g2_fill_8 FILLER_0_85_1097 ();
 sg13g2_fill_8 FILLER_0_85_1105 ();
 sg13g2_fill_8 FILLER_0_85_1113 ();
 sg13g2_fill_8 FILLER_0_85_1121 ();
 sg13g2_fill_8 FILLER_0_85_1129 ();
 sg13g2_fill_8 FILLER_0_85_1137 ();
 sg13g2_fill_8 FILLER_0_85_1145 ();
 sg13g2_fill_8 FILLER_0_85_1153 ();
 sg13g2_fill_8 FILLER_0_85_1161 ();
 sg13g2_fill_8 FILLER_0_85_1169 ();
 sg13g2_fill_8 FILLER_0_85_1177 ();
 sg13g2_fill_8 FILLER_0_85_1185 ();
 sg13g2_fill_8 FILLER_0_85_1193 ();
 sg13g2_fill_8 FILLER_0_85_1201 ();
 sg13g2_fill_8 FILLER_0_85_1209 ();
 sg13g2_fill_8 FILLER_0_85_1217 ();
 sg13g2_fill_2 FILLER_0_85_1225 ();
 sg13g2_fill_1 FILLER_0_85_1227 ();
 sg13g2_fill_1 FILLER_0_86_36 ();
 sg13g2_fill_1 FILLER_0_86_41 ();
 sg13g2_fill_2 FILLER_0_86_86 ();
 sg13g2_fill_2 FILLER_0_86_92 ();
 sg13g2_fill_4 FILLER_0_86_99 ();
 sg13g2_fill_8 FILLER_0_86_107 ();
 sg13g2_fill_2 FILLER_0_86_115 ();
 sg13g2_fill_1 FILLER_0_86_117 ();
 sg13g2_fill_1 FILLER_0_86_126 ();
 sg13g2_fill_2 FILLER_0_86_163 ();
 sg13g2_fill_4 FILLER_0_86_169 ();
 sg13g2_fill_1 FILLER_0_86_173 ();
 sg13g2_decap_8 FILLER_0_86_183 ();
 sg13g2_fill_8 FILLER_0_86_195 ();
 sg13g2_fill_8 FILLER_0_86_203 ();
 sg13g2_fill_8 FILLER_0_86_211 ();
 sg13g2_fill_8 FILLER_0_86_219 ();
 sg13g2_fill_8 FILLER_0_86_227 ();
 sg13g2_fill_8 FILLER_0_86_235 ();
 sg13g2_fill_8 FILLER_0_86_243 ();
 sg13g2_fill_8 FILLER_0_86_251 ();
 sg13g2_fill_4 FILLER_0_86_259 ();
 sg13g2_fill_1 FILLER_0_86_263 ();
 sg13g2_fill_8 FILLER_0_86_289 ();
 sg13g2_fill_8 FILLER_0_86_297 ();
 sg13g2_fill_8 FILLER_0_86_305 ();
 sg13g2_fill_4 FILLER_0_86_313 ();
 sg13g2_fill_2 FILLER_0_86_317 ();
 sg13g2_fill_4 FILLER_0_86_323 ();
 sg13g2_fill_1 FILLER_0_86_327 ();
 sg13g2_fill_8 FILLER_0_86_333 ();
 sg13g2_fill_2 FILLER_0_86_341 ();
 sg13g2_fill_4 FILLER_0_86_374 ();
 sg13g2_fill_8 FILLER_0_86_382 ();
 sg13g2_fill_4 FILLER_0_86_390 ();
 sg13g2_fill_2 FILLER_0_86_394 ();
 sg13g2_fill_8 FILLER_0_86_406 ();
 sg13g2_fill_4 FILLER_0_86_414 ();
 sg13g2_fill_8 FILLER_0_86_444 ();
 sg13g2_fill_2 FILLER_0_86_452 ();
 sg13g2_fill_1 FILLER_0_86_459 ();
 sg13g2_fill_8 FILLER_0_86_464 ();
 sg13g2_fill_8 FILLER_0_86_472 ();
 sg13g2_fill_2 FILLER_0_86_480 ();
 sg13g2_fill_1 FILLER_0_86_482 ();
 sg13g2_fill_1 FILLER_0_86_502 ();
 sg13g2_fill_1 FILLER_0_86_544 ();
 sg13g2_fill_8 FILLER_0_86_571 ();
 sg13g2_fill_2 FILLER_0_86_579 ();
 sg13g2_fill_1 FILLER_0_86_581 ();
 sg13g2_fill_8 FILLER_0_86_586 ();
 sg13g2_fill_8 FILLER_0_86_594 ();
 sg13g2_fill_4 FILLER_0_86_602 ();
 sg13g2_fill_2 FILLER_0_86_637 ();
 sg13g2_fill_1 FILLER_0_86_639 ();
 sg13g2_fill_4 FILLER_0_86_679 ();
 sg13g2_fill_1 FILLER_0_86_683 ();
 sg13g2_fill_8 FILLER_0_86_719 ();
 sg13g2_fill_4 FILLER_0_86_727 ();
 sg13g2_fill_1 FILLER_0_86_731 ();
 sg13g2_fill_1 FILLER_0_86_762 ();
 sg13g2_fill_8 FILLER_0_86_839 ();
 sg13g2_fill_2 FILLER_0_86_847 ();
 sg13g2_fill_1 FILLER_0_86_849 ();
 sg13g2_decap_8 FILLER_0_86_855 ();
 sg13g2_fill_8 FILLER_0_86_866 ();
 sg13g2_fill_8 FILLER_0_86_874 ();
 sg13g2_fill_4 FILLER_0_86_882 ();
 sg13g2_fill_1 FILLER_0_86_886 ();
 sg13g2_fill_8 FILLER_0_86_917 ();
 sg13g2_fill_4 FILLER_0_86_930 ();
 sg13g2_fill_1 FILLER_0_86_934 ();
 sg13g2_fill_8 FILLER_0_86_945 ();
 sg13g2_fill_8 FILLER_0_86_973 ();
 sg13g2_fill_8 FILLER_0_86_981 ();
 sg13g2_fill_8 FILLER_0_86_989 ();
 sg13g2_fill_8 FILLER_0_86_997 ();
 sg13g2_fill_8 FILLER_0_86_1005 ();
 sg13g2_fill_8 FILLER_0_86_1013 ();
 sg13g2_fill_8 FILLER_0_86_1021 ();
 sg13g2_fill_8 FILLER_0_86_1029 ();
 sg13g2_fill_8 FILLER_0_86_1037 ();
 sg13g2_fill_8 FILLER_0_86_1045 ();
 sg13g2_fill_8 FILLER_0_86_1053 ();
 sg13g2_fill_8 FILLER_0_86_1061 ();
 sg13g2_fill_8 FILLER_0_86_1069 ();
 sg13g2_fill_8 FILLER_0_86_1077 ();
 sg13g2_fill_8 FILLER_0_86_1085 ();
 sg13g2_fill_8 FILLER_0_86_1093 ();
 sg13g2_fill_8 FILLER_0_86_1101 ();
 sg13g2_fill_8 FILLER_0_86_1109 ();
 sg13g2_fill_8 FILLER_0_86_1117 ();
 sg13g2_fill_8 FILLER_0_86_1125 ();
 sg13g2_fill_8 FILLER_0_86_1133 ();
 sg13g2_fill_8 FILLER_0_86_1141 ();
 sg13g2_fill_8 FILLER_0_86_1149 ();
 sg13g2_fill_8 FILLER_0_86_1157 ();
 sg13g2_fill_8 FILLER_0_86_1165 ();
 sg13g2_fill_8 FILLER_0_86_1173 ();
 sg13g2_fill_8 FILLER_0_86_1181 ();
 sg13g2_fill_8 FILLER_0_86_1189 ();
 sg13g2_fill_8 FILLER_0_86_1197 ();
 sg13g2_fill_8 FILLER_0_86_1205 ();
 sg13g2_fill_8 FILLER_0_86_1213 ();
 sg13g2_decap_8 FILLER_0_86_1221 ();
 sg13g2_fill_4 FILLER_0_87_0 ();
 sg13g2_fill_1 FILLER_0_87_4 ();
 sg13g2_fill_4 FILLER_0_87_36 ();
 sg13g2_fill_8 FILLER_0_87_52 ();
 sg13g2_fill_8 FILLER_0_87_60 ();
 sg13g2_fill_2 FILLER_0_87_68 ();
 sg13g2_fill_2 FILLER_0_87_82 ();
 sg13g2_fill_2 FILLER_0_87_124 ();
 sg13g2_fill_4 FILLER_0_87_145 ();
 sg13g2_fill_8 FILLER_0_87_157 ();
 sg13g2_fill_8 FILLER_0_87_165 ();
 sg13g2_fill_8 FILLER_0_87_173 ();
 sg13g2_fill_8 FILLER_0_87_181 ();
 sg13g2_fill_8 FILLER_0_87_189 ();
 sg13g2_fill_2 FILLER_0_87_197 ();
 sg13g2_fill_8 FILLER_0_87_204 ();
 sg13g2_fill_8 FILLER_0_87_212 ();
 sg13g2_fill_1 FILLER_0_87_220 ();
 sg13g2_fill_8 FILLER_0_87_226 ();
 sg13g2_fill_8 FILLER_0_87_234 ();
 sg13g2_fill_4 FILLER_0_87_242 ();
 sg13g2_fill_2 FILLER_0_87_246 ();
 sg13g2_fill_1 FILLER_0_87_288 ();
 sg13g2_fill_8 FILLER_0_87_299 ();
 sg13g2_fill_8 FILLER_0_87_321 ();
 sg13g2_fill_2 FILLER_0_87_329 ();
 sg13g2_fill_1 FILLER_0_87_331 ();
 sg13g2_fill_2 FILLER_0_87_367 ();
 sg13g2_fill_1 FILLER_0_87_462 ();
 sg13g2_fill_8 FILLER_0_87_467 ();
 sg13g2_fill_1 FILLER_0_87_475 ();
 sg13g2_fill_1 FILLER_0_87_502 ();
 sg13g2_fill_2 FILLER_0_87_536 ();
 sg13g2_fill_1 FILLER_0_87_538 ();
 sg13g2_fill_8 FILLER_0_87_574 ();
 sg13g2_fill_8 FILLER_0_87_582 ();
 sg13g2_fill_2 FILLER_0_87_590 ();
 sg13g2_fill_1 FILLER_0_87_592 ();
 sg13g2_fill_1 FILLER_0_87_619 ();
 sg13g2_fill_8 FILLER_0_87_646 ();
 sg13g2_fill_1 FILLER_0_87_685 ();
 sg13g2_fill_8 FILLER_0_87_722 ();
 sg13g2_decap_8 FILLER_0_87_730 ();
 sg13g2_fill_1 FILLER_0_87_766 ();
 sg13g2_fill_2 FILLER_0_87_798 ();
 sg13g2_fill_2 FILLER_0_87_830 ();
 sg13g2_fill_4 FILLER_0_87_842 ();
 sg13g2_fill_8 FILLER_0_87_861 ();
 sg13g2_fill_8 FILLER_0_87_869 ();
 sg13g2_fill_2 FILLER_0_87_877 ();
 sg13g2_fill_1 FILLER_0_87_879 ();
 sg13g2_fill_8 FILLER_0_87_885 ();
 sg13g2_fill_1 FILLER_0_87_893 ();
 sg13g2_fill_4 FILLER_0_87_899 ();
 sg13g2_fill_2 FILLER_0_87_903 ();
 sg13g2_fill_2 FILLER_0_87_915 ();
 sg13g2_fill_1 FILLER_0_87_917 ();
 sg13g2_fill_8 FILLER_0_87_983 ();
 sg13g2_fill_8 FILLER_0_87_991 ();
 sg13g2_fill_8 FILLER_0_87_999 ();
 sg13g2_fill_8 FILLER_0_87_1007 ();
 sg13g2_fill_8 FILLER_0_87_1015 ();
 sg13g2_fill_8 FILLER_0_87_1023 ();
 sg13g2_fill_8 FILLER_0_87_1031 ();
 sg13g2_fill_8 FILLER_0_87_1039 ();
 sg13g2_fill_8 FILLER_0_87_1047 ();
 sg13g2_fill_8 FILLER_0_87_1055 ();
 sg13g2_fill_8 FILLER_0_87_1063 ();
 sg13g2_fill_8 FILLER_0_87_1071 ();
 sg13g2_fill_8 FILLER_0_87_1079 ();
 sg13g2_fill_8 FILLER_0_87_1087 ();
 sg13g2_fill_8 FILLER_0_87_1095 ();
 sg13g2_fill_8 FILLER_0_87_1103 ();
 sg13g2_fill_8 FILLER_0_87_1111 ();
 sg13g2_fill_8 FILLER_0_87_1119 ();
 sg13g2_fill_8 FILLER_0_87_1127 ();
 sg13g2_fill_8 FILLER_0_87_1135 ();
 sg13g2_fill_8 FILLER_0_87_1143 ();
 sg13g2_fill_8 FILLER_0_87_1151 ();
 sg13g2_fill_8 FILLER_0_87_1159 ();
 sg13g2_fill_8 FILLER_0_87_1167 ();
 sg13g2_fill_8 FILLER_0_87_1175 ();
 sg13g2_fill_8 FILLER_0_87_1183 ();
 sg13g2_fill_8 FILLER_0_87_1191 ();
 sg13g2_fill_8 FILLER_0_87_1199 ();
 sg13g2_fill_8 FILLER_0_87_1207 ();
 sg13g2_fill_8 FILLER_0_87_1215 ();
 sg13g2_fill_4 FILLER_0_87_1223 ();
 sg13g2_fill_1 FILLER_0_87_1227 ();
 sg13g2_fill_8 FILLER_0_88_0 ();
 sg13g2_fill_4 FILLER_0_88_8 ();
 sg13g2_fill_8 FILLER_0_88_16 ();
 sg13g2_fill_1 FILLER_0_88_24 ();
 sg13g2_fill_4 FILLER_0_88_66 ();
 sg13g2_fill_1 FILLER_0_88_70 ();
 sg13g2_fill_8 FILLER_0_88_75 ();
 sg13g2_decap_8 FILLER_0_88_83 ();
 sg13g2_fill_8 FILLER_0_88_94 ();
 sg13g2_fill_8 FILLER_0_88_102 ();
 sg13g2_fill_8 FILLER_0_88_110 ();
 sg13g2_fill_8 FILLER_0_88_118 ();
 sg13g2_fill_8 FILLER_0_88_126 ();
 sg13g2_fill_8 FILLER_0_88_134 ();
 sg13g2_fill_2 FILLER_0_88_142 ();
 sg13g2_fill_1 FILLER_0_88_144 ();
 sg13g2_fill_1 FILLER_0_88_153 ();
 sg13g2_fill_1 FILLER_0_88_162 ();
 sg13g2_fill_1 FILLER_0_88_168 ();
 sg13g2_fill_1 FILLER_0_88_195 ();
 sg13g2_fill_1 FILLER_0_88_226 ();
 sg13g2_fill_2 FILLER_0_88_253 ();
 sg13g2_fill_1 FILLER_0_88_286 ();
 sg13g2_fill_8 FILLER_0_88_333 ();
 sg13g2_fill_2 FILLER_0_88_407 ();
 sg13g2_fill_1 FILLER_0_88_419 ();
 sg13g2_fill_1 FILLER_0_88_430 ();
 sg13g2_fill_2 FILLER_0_88_436 ();
 sg13g2_fill_2 FILLER_0_88_448 ();
 sg13g2_fill_1 FILLER_0_88_450 ();
 sg13g2_fill_2 FILLER_0_88_481 ();
 sg13g2_fill_1 FILLER_0_88_483 ();
 sg13g2_fill_4 FILLER_0_88_524 ();
 sg13g2_fill_2 FILLER_0_88_528 ();
 sg13g2_fill_8 FILLER_0_88_564 ();
 sg13g2_fill_8 FILLER_0_88_572 ();
 sg13g2_fill_8 FILLER_0_88_580 ();
 sg13g2_fill_8 FILLER_0_88_588 ();
 sg13g2_fill_2 FILLER_0_88_596 ();
 sg13g2_fill_1 FILLER_0_88_642 ();
 sg13g2_fill_2 FILLER_0_88_703 ();
 sg13g2_fill_2 FILLER_0_88_720 ();
 sg13g2_fill_8 FILLER_0_88_726 ();
 sg13g2_fill_8 FILLER_0_88_734 ();
 sg13g2_fill_2 FILLER_0_88_742 ();
 sg13g2_fill_1 FILLER_0_88_744 ();
 sg13g2_fill_2 FILLER_0_88_749 ();
 sg13g2_fill_2 FILLER_0_88_755 ();
 sg13g2_fill_2 FILLER_0_88_767 ();
 sg13g2_fill_2 FILLER_0_88_774 ();
 sg13g2_fill_1 FILLER_0_88_776 ();
 sg13g2_fill_2 FILLER_0_88_781 ();
 sg13g2_fill_1 FILLER_0_88_783 ();
 sg13g2_fill_2 FILLER_0_88_788 ();
 sg13g2_fill_1 FILLER_0_88_790 ();
 sg13g2_fill_1 FILLER_0_88_809 ();
 sg13g2_fill_1 FILLER_0_88_888 ();
 sg13g2_fill_1 FILLER_0_88_894 ();
 sg13g2_fill_1 FILLER_0_88_905 ();
 sg13g2_fill_1 FILLER_0_88_916 ();
 sg13g2_fill_1 FILLER_0_88_921 ();
 sg13g2_decap_8 FILLER_0_88_949 ();
 sg13g2_fill_8 FILLER_0_88_987 ();
 sg13g2_fill_8 FILLER_0_88_995 ();
 sg13g2_fill_8 FILLER_0_88_1003 ();
 sg13g2_fill_8 FILLER_0_88_1011 ();
 sg13g2_fill_8 FILLER_0_88_1019 ();
 sg13g2_fill_8 FILLER_0_88_1027 ();
 sg13g2_fill_8 FILLER_0_88_1035 ();
 sg13g2_fill_8 FILLER_0_88_1043 ();
 sg13g2_fill_8 FILLER_0_88_1051 ();
 sg13g2_fill_8 FILLER_0_88_1059 ();
 sg13g2_fill_8 FILLER_0_88_1067 ();
 sg13g2_fill_8 FILLER_0_88_1075 ();
 sg13g2_fill_8 FILLER_0_88_1083 ();
 sg13g2_fill_8 FILLER_0_88_1091 ();
 sg13g2_fill_8 FILLER_0_88_1099 ();
 sg13g2_fill_8 FILLER_0_88_1107 ();
 sg13g2_fill_8 FILLER_0_88_1115 ();
 sg13g2_fill_8 FILLER_0_88_1123 ();
 sg13g2_fill_8 FILLER_0_88_1131 ();
 sg13g2_fill_8 FILLER_0_88_1139 ();
 sg13g2_fill_8 FILLER_0_88_1147 ();
 sg13g2_fill_8 FILLER_0_88_1155 ();
 sg13g2_fill_8 FILLER_0_88_1163 ();
 sg13g2_fill_8 FILLER_0_88_1171 ();
 sg13g2_fill_8 FILLER_0_88_1179 ();
 sg13g2_fill_8 FILLER_0_88_1187 ();
 sg13g2_fill_8 FILLER_0_88_1195 ();
 sg13g2_fill_8 FILLER_0_88_1203 ();
 sg13g2_fill_8 FILLER_0_88_1211 ();
 sg13g2_fill_8 FILLER_0_88_1219 ();
 sg13g2_fill_1 FILLER_0_88_1227 ();
 sg13g2_fill_8 FILLER_0_89_0 ();
 sg13g2_fill_8 FILLER_0_89_8 ();
 sg13g2_fill_1 FILLER_0_89_20 ();
 sg13g2_fill_1 FILLER_0_89_31 ();
 sg13g2_fill_1 FILLER_0_89_47 ();
 sg13g2_fill_4 FILLER_0_89_52 ();
 sg13g2_fill_2 FILLER_0_89_61 ();
 sg13g2_fill_1 FILLER_0_89_63 ();
 sg13g2_fill_2 FILLER_0_89_100 ();
 sg13g2_fill_2 FILLER_0_89_107 ();
 sg13g2_fill_2 FILLER_0_89_119 ();
 sg13g2_fill_4 FILLER_0_89_131 ();
 sg13g2_fill_2 FILLER_0_89_135 ();
 sg13g2_decap_8 FILLER_0_89_251 ();
 sg13g2_fill_1 FILLER_0_89_267 ();
 sg13g2_decap_8 FILLER_0_89_325 ();
 sg13g2_fill_4 FILLER_0_89_368 ();
 sg13g2_fill_2 FILLER_0_89_372 ();
 sg13g2_fill_4 FILLER_0_89_378 ();
 sg13g2_fill_2 FILLER_0_89_382 ();
 sg13g2_fill_8 FILLER_0_89_388 ();
 sg13g2_fill_2 FILLER_0_89_396 ();
 sg13g2_fill_1 FILLER_0_89_398 ();
 sg13g2_fill_4 FILLER_0_89_413 ();
 sg13g2_fill_4 FILLER_0_89_422 ();
 sg13g2_fill_2 FILLER_0_89_430 ();
 sg13g2_fill_1 FILLER_0_89_432 ();
 sg13g2_fill_8 FILLER_0_89_437 ();
 sg13g2_fill_2 FILLER_0_89_445 ();
 sg13g2_fill_1 FILLER_0_89_447 ();
 sg13g2_fill_4 FILLER_0_89_474 ();
 sg13g2_fill_8 FILLER_0_89_514 ();
 sg13g2_fill_4 FILLER_0_89_522 ();
 sg13g2_fill_1 FILLER_0_89_526 ();
 sg13g2_fill_8 FILLER_0_89_557 ();
 sg13g2_fill_2 FILLER_0_89_565 ();
 sg13g2_fill_1 FILLER_0_89_567 ();
 sg13g2_fill_2 FILLER_0_89_599 ();
 sg13g2_fill_1 FILLER_0_89_601 ();
 sg13g2_fill_2 FILLER_0_89_610 ();
 sg13g2_fill_1 FILLER_0_89_626 ();
 sg13g2_fill_8 FILLER_0_89_631 ();
 sg13g2_fill_8 FILLER_0_89_639 ();
 sg13g2_fill_1 FILLER_0_89_647 ();
 sg13g2_fill_2 FILLER_0_89_657 ();
 sg13g2_fill_8 FILLER_0_89_669 ();
 sg13g2_fill_8 FILLER_0_89_677 ();
 sg13g2_fill_8 FILLER_0_89_685 ();
 sg13g2_fill_4 FILLER_0_89_693 ();
 sg13g2_fill_1 FILLER_0_89_697 ();
 sg13g2_fill_2 FILLER_0_89_708 ();
 sg13g2_fill_1 FILLER_0_89_710 ();
 sg13g2_fill_8 FILLER_0_89_768 ();
 sg13g2_fill_8 FILLER_0_89_776 ();
 sg13g2_fill_8 FILLER_0_89_784 ();
 sg13g2_fill_2 FILLER_0_89_792 ();
 sg13g2_fill_1 FILLER_0_89_794 ();
 sg13g2_fill_4 FILLER_0_89_803 ();
 sg13g2_fill_2 FILLER_0_89_823 ();
 sg13g2_fill_1 FILLER_0_89_825 ();
 sg13g2_fill_2 FILLER_0_89_830 ();
 sg13g2_fill_1 FILLER_0_89_832 ();
 sg13g2_fill_2 FILLER_0_89_845 ();
 sg13g2_fill_2 FILLER_0_89_873 ();
 sg13g2_fill_1 FILLER_0_89_875 ();
 sg13g2_fill_2 FILLER_0_89_902 ();
 sg13g2_fill_1 FILLER_0_89_904 ();
 sg13g2_decap_8 FILLER_0_89_931 ();
 sg13g2_fill_8 FILLER_0_89_972 ();
 sg13g2_fill_8 FILLER_0_89_980 ();
 sg13g2_fill_8 FILLER_0_89_988 ();
 sg13g2_fill_8 FILLER_0_89_996 ();
 sg13g2_fill_8 FILLER_0_89_1004 ();
 sg13g2_fill_8 FILLER_0_89_1012 ();
 sg13g2_fill_8 FILLER_0_89_1020 ();
 sg13g2_fill_8 FILLER_0_89_1028 ();
 sg13g2_fill_8 FILLER_0_89_1036 ();
 sg13g2_fill_8 FILLER_0_89_1044 ();
 sg13g2_fill_8 FILLER_0_89_1052 ();
 sg13g2_fill_8 FILLER_0_89_1060 ();
 sg13g2_fill_8 FILLER_0_89_1068 ();
 sg13g2_fill_8 FILLER_0_89_1076 ();
 sg13g2_fill_8 FILLER_0_89_1084 ();
 sg13g2_fill_8 FILLER_0_89_1092 ();
 sg13g2_fill_8 FILLER_0_89_1100 ();
 sg13g2_fill_8 FILLER_0_89_1108 ();
 sg13g2_fill_8 FILLER_0_89_1116 ();
 sg13g2_fill_8 FILLER_0_89_1124 ();
 sg13g2_fill_8 FILLER_0_89_1132 ();
 sg13g2_fill_8 FILLER_0_89_1140 ();
 sg13g2_fill_8 FILLER_0_89_1148 ();
 sg13g2_fill_8 FILLER_0_89_1156 ();
 sg13g2_fill_8 FILLER_0_89_1164 ();
 sg13g2_fill_8 FILLER_0_89_1172 ();
 sg13g2_fill_8 FILLER_0_89_1180 ();
 sg13g2_fill_8 FILLER_0_89_1188 ();
 sg13g2_fill_8 FILLER_0_89_1196 ();
 sg13g2_fill_8 FILLER_0_89_1204 ();
 sg13g2_fill_8 FILLER_0_89_1212 ();
 sg13g2_fill_8 FILLER_0_89_1220 ();
 sg13g2_fill_4 FILLER_0_90_0 ();
 sg13g2_fill_2 FILLER_0_90_4 ();
 sg13g2_fill_2 FILLER_0_90_37 ();
 sg13g2_fill_8 FILLER_0_90_69 ();
 sg13g2_fill_1 FILLER_0_90_81 ();
 sg13g2_fill_2 FILLER_0_90_134 ();
 sg13g2_fill_2 FILLER_0_90_198 ();
 sg13g2_fill_1 FILLER_0_90_200 ();
 sg13g2_fill_1 FILLER_0_90_211 ();
 sg13g2_fill_2 FILLER_0_90_241 ();
 sg13g2_fill_8 FILLER_0_90_251 ();
 sg13g2_fill_8 FILLER_0_90_259 ();
 sg13g2_fill_8 FILLER_0_90_267 ();
 sg13g2_fill_8 FILLER_0_90_279 ();
 sg13g2_fill_2 FILLER_0_90_287 ();
 sg13g2_fill_1 FILLER_0_90_289 ();
 sg13g2_fill_8 FILLER_0_90_316 ();
 sg13g2_fill_8 FILLER_0_90_324 ();
 sg13g2_fill_2 FILLER_0_90_332 ();
 sg13g2_fill_1 FILLER_0_90_334 ();
 sg13g2_fill_4 FILLER_0_90_343 ();
 sg13g2_fill_1 FILLER_0_90_347 ();
 sg13g2_fill_1 FILLER_0_90_368 ();
 sg13g2_fill_4 FILLER_0_90_395 ();
 sg13g2_fill_2 FILLER_0_90_399 ();
 sg13g2_fill_8 FILLER_0_90_410 ();
 sg13g2_fill_8 FILLER_0_90_418 ();
 sg13g2_fill_8 FILLER_0_90_436 ();
 sg13g2_fill_2 FILLER_0_90_444 ();
 sg13g2_fill_8 FILLER_0_90_475 ();
 sg13g2_fill_2 FILLER_0_90_483 ();
 sg13g2_fill_8 FILLER_0_90_489 ();
 sg13g2_fill_2 FILLER_0_90_497 ();
 sg13g2_fill_1 FILLER_0_90_499 ();
 sg13g2_fill_8 FILLER_0_90_504 ();
 sg13g2_fill_4 FILLER_0_90_512 ();
 sg13g2_fill_1 FILLER_0_90_516 ();
 sg13g2_fill_4 FILLER_0_90_522 ();
 sg13g2_fill_2 FILLER_0_90_526 ();
 sg13g2_fill_2 FILLER_0_90_533 ();
 sg13g2_decap_8 FILLER_0_90_555 ();
 sg13g2_fill_8 FILLER_0_90_634 ();
 sg13g2_decap_8 FILLER_0_90_642 ();
 sg13g2_fill_2 FILLER_0_90_661 ();
 sg13g2_fill_8 FILLER_0_90_667 ();
 sg13g2_fill_4 FILLER_0_90_675 ();
 sg13g2_decap_8 FILLER_0_90_683 ();
 sg13g2_fill_4 FILLER_0_90_726 ();
 sg13g2_fill_1 FILLER_0_90_730 ();
 sg13g2_fill_2 FILLER_0_90_772 ();
 sg13g2_fill_1 FILLER_0_90_797 ();
 sg13g2_fill_8 FILLER_0_90_808 ();
 sg13g2_fill_4 FILLER_0_90_816 ();
 sg13g2_fill_2 FILLER_0_90_820 ();
 sg13g2_fill_8 FILLER_0_90_832 ();
 sg13g2_fill_4 FILLER_0_90_840 ();
 sg13g2_fill_2 FILLER_0_90_844 ();
 sg13g2_fill_2 FILLER_0_90_855 ();
 sg13g2_fill_1 FILLER_0_90_857 ();
 sg13g2_fill_1 FILLER_0_90_868 ();
 sg13g2_fill_1 FILLER_0_90_873 ();
 sg13g2_fill_1 FILLER_0_90_884 ();
 sg13g2_fill_2 FILLER_0_90_895 ();
 sg13g2_fill_8 FILLER_0_90_928 ();
 sg13g2_fill_8 FILLER_0_90_936 ();
 sg13g2_fill_2 FILLER_0_90_944 ();
 sg13g2_fill_8 FILLER_0_90_950 ();
 sg13g2_fill_8 FILLER_0_90_958 ();
 sg13g2_fill_8 FILLER_0_90_966 ();
 sg13g2_fill_8 FILLER_0_90_974 ();
 sg13g2_fill_8 FILLER_0_90_982 ();
 sg13g2_fill_8 FILLER_0_90_990 ();
 sg13g2_fill_8 FILLER_0_90_998 ();
 sg13g2_fill_8 FILLER_0_90_1006 ();
 sg13g2_fill_8 FILLER_0_90_1014 ();
 sg13g2_fill_8 FILLER_0_90_1022 ();
 sg13g2_fill_8 FILLER_0_90_1030 ();
 sg13g2_fill_8 FILLER_0_90_1038 ();
 sg13g2_fill_8 FILLER_0_90_1046 ();
 sg13g2_fill_8 FILLER_0_90_1054 ();
 sg13g2_fill_8 FILLER_0_90_1062 ();
 sg13g2_fill_8 FILLER_0_90_1070 ();
 sg13g2_fill_8 FILLER_0_90_1078 ();
 sg13g2_fill_8 FILLER_0_90_1086 ();
 sg13g2_fill_8 FILLER_0_90_1094 ();
 sg13g2_fill_8 FILLER_0_90_1102 ();
 sg13g2_fill_8 FILLER_0_90_1110 ();
 sg13g2_fill_8 FILLER_0_90_1118 ();
 sg13g2_fill_8 FILLER_0_90_1126 ();
 sg13g2_fill_8 FILLER_0_90_1134 ();
 sg13g2_fill_8 FILLER_0_90_1142 ();
 sg13g2_fill_8 FILLER_0_90_1150 ();
 sg13g2_fill_8 FILLER_0_90_1158 ();
 sg13g2_fill_8 FILLER_0_90_1166 ();
 sg13g2_fill_8 FILLER_0_90_1174 ();
 sg13g2_fill_8 FILLER_0_90_1182 ();
 sg13g2_fill_8 FILLER_0_90_1190 ();
 sg13g2_fill_8 FILLER_0_90_1198 ();
 sg13g2_fill_8 FILLER_0_90_1206 ();
 sg13g2_fill_8 FILLER_0_90_1214 ();
 sg13g2_fill_4 FILLER_0_90_1222 ();
 sg13g2_fill_2 FILLER_0_90_1226 ();
 sg13g2_fill_1 FILLER_0_91_0 ();
 sg13g2_fill_1 FILLER_0_91_27 ();
 sg13g2_fill_1 FILLER_0_91_38 ();
 sg13g2_fill_2 FILLER_0_91_47 ();
 sg13g2_fill_2 FILLER_0_91_57 ();
 sg13g2_fill_1 FILLER_0_91_59 ();
 sg13g2_fill_8 FILLER_0_91_69 ();
 sg13g2_fill_8 FILLER_0_91_77 ();
 sg13g2_fill_2 FILLER_0_91_85 ();
 sg13g2_fill_2 FILLER_0_91_135 ();
 sg13g2_fill_1 FILLER_0_91_156 ();
 sg13g2_fill_8 FILLER_0_91_172 ();
 sg13g2_fill_1 FILLER_0_91_190 ();
 sg13g2_fill_8 FILLER_0_91_196 ();
 sg13g2_fill_4 FILLER_0_91_204 ();
 sg13g2_fill_1 FILLER_0_91_208 ();
 sg13g2_fill_8 FILLER_0_91_213 ();
 sg13g2_fill_1 FILLER_0_91_221 ();
 sg13g2_fill_4 FILLER_0_91_227 ();
 sg13g2_fill_8 FILLER_0_91_239 ();
 sg13g2_fill_8 FILLER_0_91_247 ();
 sg13g2_decap_8 FILLER_0_91_255 ();
 sg13g2_fill_4 FILLER_0_91_266 ();
 sg13g2_fill_1 FILLER_0_91_270 ();
 sg13g2_fill_8 FILLER_0_91_276 ();
 sg13g2_fill_8 FILLER_0_91_284 ();
 sg13g2_fill_4 FILLER_0_91_292 ();
 sg13g2_fill_2 FILLER_0_91_296 ();
 sg13g2_fill_4 FILLER_0_91_302 ();
 sg13g2_fill_2 FILLER_0_91_306 ();
 sg13g2_fill_8 FILLER_0_91_312 ();
 sg13g2_fill_8 FILLER_0_91_320 ();
 sg13g2_fill_1 FILLER_0_91_328 ();
 sg13g2_fill_4 FILLER_0_91_365 ();
 sg13g2_fill_1 FILLER_0_91_369 ();
 sg13g2_fill_8 FILLER_0_91_378 ();
 sg13g2_fill_8 FILLER_0_91_386 ();
 sg13g2_fill_8 FILLER_0_91_394 ();
 sg13g2_fill_1 FILLER_0_91_402 ();
 sg13g2_fill_2 FILLER_0_91_438 ();
 sg13g2_fill_1 FILLER_0_91_440 ();
 sg13g2_fill_1 FILLER_0_91_446 ();
 sg13g2_fill_1 FILLER_0_91_457 ();
 sg13g2_fill_1 FILLER_0_91_484 ();
 sg13g2_fill_2 FILLER_0_91_489 ();
 sg13g2_fill_1 FILLER_0_91_491 ();
 sg13g2_fill_8 FILLER_0_91_497 ();
 sg13g2_fill_8 FILLER_0_91_505 ();
 sg13g2_fill_1 FILLER_0_91_575 ();
 sg13g2_fill_1 FILLER_0_91_581 ();
 sg13g2_fill_4 FILLER_0_91_586 ();
 sg13g2_fill_8 FILLER_0_91_594 ();
 sg13g2_fill_8 FILLER_0_91_641 ();
 sg13g2_fill_2 FILLER_0_91_712 ();
 sg13g2_fill_8 FILLER_0_91_718 ();
 sg13g2_decap_8 FILLER_0_91_726 ();
 sg13g2_fill_8 FILLER_0_91_853 ();
 sg13g2_fill_8 FILLER_0_91_861 ();
 sg13g2_fill_8 FILLER_0_91_869 ();
 sg13g2_decap_8 FILLER_0_91_877 ();
 sg13g2_fill_8 FILLER_0_91_888 ();
 sg13g2_fill_4 FILLER_0_91_896 ();
 sg13g2_fill_2 FILLER_0_91_900 ();
 sg13g2_fill_2 FILLER_0_91_907 ();
 sg13g2_fill_1 FILLER_0_91_909 ();
 sg13g2_fill_4 FILLER_0_91_914 ();
 sg13g2_fill_2 FILLER_0_91_918 ();
 sg13g2_fill_8 FILLER_0_91_929 ();
 sg13g2_fill_8 FILLER_0_91_937 ();
 sg13g2_fill_2 FILLER_0_91_945 ();
 sg13g2_fill_1 FILLER_0_91_947 ();
 sg13g2_fill_8 FILLER_0_91_958 ();
 sg13g2_fill_2 FILLER_0_91_966 ();
 sg13g2_fill_1 FILLER_0_91_968 ();
 sg13g2_fill_8 FILLER_0_91_986 ();
 sg13g2_fill_8 FILLER_0_91_994 ();
 sg13g2_fill_8 FILLER_0_91_1002 ();
 sg13g2_fill_8 FILLER_0_91_1010 ();
 sg13g2_fill_8 FILLER_0_91_1018 ();
 sg13g2_fill_8 FILLER_0_91_1026 ();
 sg13g2_fill_8 FILLER_0_91_1034 ();
 sg13g2_fill_8 FILLER_0_91_1042 ();
 sg13g2_fill_8 FILLER_0_91_1050 ();
 sg13g2_fill_2 FILLER_0_91_1058 ();
 sg13g2_fill_1 FILLER_0_91_1060 ();
 sg13g2_fill_8 FILLER_0_91_1065 ();
 sg13g2_fill_8 FILLER_0_91_1073 ();
 sg13g2_fill_8 FILLER_0_91_1081 ();
 sg13g2_fill_8 FILLER_0_91_1089 ();
 sg13g2_fill_8 FILLER_0_91_1097 ();
 sg13g2_fill_8 FILLER_0_91_1105 ();
 sg13g2_fill_8 FILLER_0_91_1113 ();
 sg13g2_fill_8 FILLER_0_91_1121 ();
 sg13g2_fill_8 FILLER_0_91_1129 ();
 sg13g2_fill_8 FILLER_0_91_1137 ();
 sg13g2_fill_8 FILLER_0_91_1145 ();
 sg13g2_fill_8 FILLER_0_91_1153 ();
 sg13g2_fill_8 FILLER_0_91_1161 ();
 sg13g2_fill_8 FILLER_0_91_1169 ();
 sg13g2_fill_8 FILLER_0_91_1177 ();
 sg13g2_fill_8 FILLER_0_91_1185 ();
 sg13g2_fill_8 FILLER_0_91_1193 ();
 sg13g2_fill_8 FILLER_0_91_1201 ();
 sg13g2_fill_8 FILLER_0_91_1209 ();
 sg13g2_fill_8 FILLER_0_91_1217 ();
 sg13g2_fill_2 FILLER_0_91_1225 ();
 sg13g2_fill_1 FILLER_0_91_1227 ();
 sg13g2_fill_2 FILLER_0_92_0 ();
 sg13g2_fill_2 FILLER_0_92_52 ();
 sg13g2_fill_1 FILLER_0_92_54 ();
 sg13g2_fill_4 FILLER_0_92_93 ();
 sg13g2_fill_1 FILLER_0_92_97 ();
 sg13g2_fill_1 FILLER_0_92_130 ();
 sg13g2_fill_2 FILLER_0_92_161 ();
 sg13g2_fill_1 FILLER_0_92_163 ();
 sg13g2_fill_8 FILLER_0_92_168 ();
 sg13g2_fill_4 FILLER_0_92_176 ();
 sg13g2_fill_2 FILLER_0_92_180 ();
 sg13g2_fill_1 FILLER_0_92_213 ();
 sg13g2_fill_4 FILLER_0_92_250 ();
 sg13g2_fill_1 FILLER_0_92_254 ();
 sg13g2_fill_8 FILLER_0_92_291 ();
 sg13g2_fill_8 FILLER_0_92_299 ();
 sg13g2_fill_8 FILLER_0_92_307 ();
 sg13g2_fill_8 FILLER_0_92_315 ();
 sg13g2_fill_1 FILLER_0_92_331 ();
 sg13g2_fill_2 FILLER_0_92_358 ();
 sg13g2_fill_1 FILLER_0_92_360 ();
 sg13g2_fill_2 FILLER_0_92_366 ();
 sg13g2_fill_1 FILLER_0_92_368 ();
 sg13g2_fill_4 FILLER_0_92_395 ();
 sg13g2_fill_1 FILLER_0_92_473 ();
 sg13g2_fill_2 FILLER_0_92_484 ();
 sg13g2_fill_1 FILLER_0_92_486 ();
 sg13g2_fill_2 FILLER_0_92_495 ();
 sg13g2_fill_8 FILLER_0_92_588 ();
 sg13g2_fill_8 FILLER_0_92_596 ();
 sg13g2_fill_8 FILLER_0_92_604 ();
 sg13g2_fill_1 FILLER_0_92_612 ();
 sg13g2_fill_2 FILLER_0_92_617 ();
 sg13g2_fill_1 FILLER_0_92_676 ();
 sg13g2_fill_8 FILLER_0_92_708 ();
 sg13g2_fill_8 FILLER_0_92_716 ();
 sg13g2_fill_8 FILLER_0_92_724 ();
 sg13g2_decap_8 FILLER_0_92_732 ();
 sg13g2_fill_2 FILLER_0_92_770 ();
 sg13g2_fill_2 FILLER_0_92_860 ();
 sg13g2_fill_1 FILLER_0_92_862 ();
 sg13g2_fill_1 FILLER_0_92_867 ();
 sg13g2_fill_2 FILLER_0_92_871 ();
 sg13g2_fill_8 FILLER_0_92_878 ();
 sg13g2_fill_1 FILLER_0_92_886 ();
 sg13g2_fill_4 FILLER_0_92_905 ();
 sg13g2_fill_1 FILLER_0_92_909 ();
 sg13g2_fill_1 FILLER_0_92_928 ();
 sg13g2_fill_2 FILLER_0_92_952 ();
 sg13g2_fill_2 FILLER_0_92_959 ();
 sg13g2_fill_1 FILLER_0_92_973 ();
 sg13g2_fill_1 FILLER_0_92_979 ();
 sg13g2_fill_8 FILLER_0_92_988 ();
 sg13g2_fill_8 FILLER_0_92_996 ();
 sg13g2_fill_8 FILLER_0_92_1004 ();
 sg13g2_fill_8 FILLER_0_92_1012 ();
 sg13g2_fill_1 FILLER_0_92_1020 ();
 sg13g2_fill_8 FILLER_0_92_1025 ();
 sg13g2_fill_2 FILLER_0_92_1038 ();
 sg13g2_fill_8 FILLER_0_92_1077 ();
 sg13g2_fill_8 FILLER_0_92_1085 ();
 sg13g2_fill_8 FILLER_0_92_1093 ();
 sg13g2_fill_8 FILLER_0_92_1101 ();
 sg13g2_fill_8 FILLER_0_92_1109 ();
 sg13g2_fill_8 FILLER_0_92_1117 ();
 sg13g2_fill_8 FILLER_0_92_1125 ();
 sg13g2_fill_8 FILLER_0_92_1133 ();
 sg13g2_fill_8 FILLER_0_92_1141 ();
 sg13g2_fill_8 FILLER_0_92_1149 ();
 sg13g2_fill_8 FILLER_0_92_1157 ();
 sg13g2_fill_8 FILLER_0_92_1165 ();
 sg13g2_fill_8 FILLER_0_92_1173 ();
 sg13g2_fill_8 FILLER_0_92_1181 ();
 sg13g2_fill_8 FILLER_0_92_1189 ();
 sg13g2_fill_8 FILLER_0_92_1197 ();
 sg13g2_fill_8 FILLER_0_92_1205 ();
 sg13g2_fill_8 FILLER_0_92_1213 ();
 sg13g2_decap_8 FILLER_0_92_1221 ();
 sg13g2_fill_8 FILLER_0_93_0 ();
 sg13g2_fill_2 FILLER_0_93_8 ();
 sg13g2_fill_4 FILLER_0_93_28 ();
 sg13g2_fill_8 FILLER_0_93_36 ();
 sg13g2_fill_1 FILLER_0_93_44 ();
 sg13g2_fill_1 FILLER_0_93_85 ();
 sg13g2_fill_2 FILLER_0_93_109 ();
 sg13g2_fill_2 FILLER_0_93_136 ();
 sg13g2_fill_1 FILLER_0_93_138 ();
 sg13g2_fill_2 FILLER_0_93_162 ();
 sg13g2_fill_2 FILLER_0_93_199 ();
 sg13g2_fill_2 FILLER_0_93_253 ();
 sg13g2_fill_2 FILLER_0_93_260 ();
 sg13g2_fill_1 FILLER_0_93_262 ();
 sg13g2_fill_1 FILLER_0_93_273 ();
 sg13g2_fill_2 FILLER_0_93_300 ();
 sg13g2_fill_2 FILLER_0_93_341 ();
 sg13g2_fill_1 FILLER_0_93_369 ();
 sg13g2_fill_2 FILLER_0_93_400 ();
 sg13g2_fill_1 FILLER_0_93_402 ();
 sg13g2_fill_1 FILLER_0_93_413 ();
 sg13g2_fill_1 FILLER_0_93_418 ();
 sg13g2_fill_8 FILLER_0_93_427 ();
 sg13g2_fill_1 FILLER_0_93_435 ();
 sg13g2_fill_2 FILLER_0_93_466 ();
 sg13g2_fill_2 FILLER_0_93_503 ();
 sg13g2_fill_1 FILLER_0_93_509 ();
 sg13g2_fill_2 FILLER_0_93_514 ();
 sg13g2_decap_8 FILLER_0_93_530 ();
 sg13g2_fill_8 FILLER_0_93_595 ();
 sg13g2_fill_4 FILLER_0_93_608 ();
 sg13g2_fill_1 FILLER_0_93_612 ();
 sg13g2_fill_1 FILLER_0_93_623 ();
 sg13g2_fill_1 FILLER_0_93_634 ();
 sg13g2_fill_2 FILLER_0_93_645 ();
 sg13g2_fill_1 FILLER_0_93_647 ();
 sg13g2_fill_2 FILLER_0_93_653 ();
 sg13g2_fill_1 FILLER_0_93_655 ();
 sg13g2_fill_8 FILLER_0_93_666 ();
 sg13g2_fill_4 FILLER_0_93_674 ();
 sg13g2_fill_1 FILLER_0_93_678 ();
 sg13g2_fill_4 FILLER_0_93_691 ();
 sg13g2_fill_2 FILLER_0_93_695 ();
 sg13g2_fill_2 FILLER_0_93_742 ();
 sg13g2_fill_1 FILLER_0_93_748 ();
 sg13g2_fill_1 FILLER_0_93_759 ();
 sg13g2_fill_1 FILLER_0_93_810 ();
 sg13g2_fill_1 FILLER_0_93_849 ();
 sg13g2_fill_1 FILLER_0_93_927 ();
 sg13g2_fill_1 FILLER_0_93_933 ();
 sg13g2_fill_2 FILLER_0_93_939 ();
 sg13g2_fill_1 FILLER_0_93_941 ();
 sg13g2_fill_1 FILLER_0_93_948 ();
 sg13g2_fill_1 FILLER_0_93_958 ();
 sg13g2_fill_8 FILLER_0_93_1004 ();
 sg13g2_fill_2 FILLER_0_93_1012 ();
 sg13g2_fill_2 FILLER_0_93_1040 ();
 sg13g2_fill_2 FILLER_0_93_1057 ();
 sg13g2_fill_1 FILLER_0_93_1059 ();
 sg13g2_fill_8 FILLER_0_93_1078 ();
 sg13g2_fill_8 FILLER_0_93_1086 ();
 sg13g2_fill_8 FILLER_0_93_1094 ();
 sg13g2_fill_8 FILLER_0_93_1102 ();
 sg13g2_fill_8 FILLER_0_93_1110 ();
 sg13g2_fill_8 FILLER_0_93_1118 ();
 sg13g2_fill_8 FILLER_0_93_1126 ();
 sg13g2_fill_8 FILLER_0_93_1134 ();
 sg13g2_fill_8 FILLER_0_93_1142 ();
 sg13g2_fill_8 FILLER_0_93_1150 ();
 sg13g2_fill_8 FILLER_0_93_1158 ();
 sg13g2_fill_8 FILLER_0_93_1166 ();
 sg13g2_fill_8 FILLER_0_93_1174 ();
 sg13g2_fill_8 FILLER_0_93_1182 ();
 sg13g2_fill_8 FILLER_0_93_1190 ();
 sg13g2_fill_8 FILLER_0_93_1198 ();
 sg13g2_fill_8 FILLER_0_93_1206 ();
 sg13g2_fill_8 FILLER_0_93_1214 ();
 sg13g2_fill_4 FILLER_0_93_1222 ();
 sg13g2_fill_2 FILLER_0_93_1226 ();
 sg13g2_fill_1 FILLER_0_94_0 ();
 sg13g2_fill_4 FILLER_0_94_27 ();
 sg13g2_fill_1 FILLER_0_94_31 ();
 sg13g2_fill_8 FILLER_0_94_37 ();
 sg13g2_fill_8 FILLER_0_94_45 ();
 sg13g2_fill_1 FILLER_0_94_53 ();
 sg13g2_fill_2 FILLER_0_94_59 ();
 sg13g2_fill_1 FILLER_0_94_81 ();
 sg13g2_fill_1 FILLER_0_94_92 ();
 sg13g2_fill_2 FILLER_0_94_119 ();
 sg13g2_fill_4 FILLER_0_94_151 ();
 sg13g2_fill_1 FILLER_0_94_155 ();
 sg13g2_fill_4 FILLER_0_94_168 ();
 sg13g2_fill_1 FILLER_0_94_172 ();
 sg13g2_fill_1 FILLER_0_94_239 ();
 sg13g2_decap_8 FILLER_0_94_244 ();
 sg13g2_fill_1 FILLER_0_94_306 ();
 sg13g2_fill_2 FILLER_0_94_341 ();
 sg13g2_fill_1 FILLER_0_94_352 ();
 sg13g2_fill_1 FILLER_0_94_373 ();
 sg13g2_fill_8 FILLER_0_94_396 ();
 sg13g2_fill_1 FILLER_0_94_404 ();
 sg13g2_fill_2 FILLER_0_94_409 ();
 sg13g2_fill_8 FILLER_0_94_415 ();
 sg13g2_fill_8 FILLER_0_94_423 ();
 sg13g2_fill_2 FILLER_0_94_431 ();
 sg13g2_fill_1 FILLER_0_94_433 ();
 sg13g2_fill_2 FILLER_0_94_447 ();
 sg13g2_fill_2 FILLER_0_94_453 ();
 sg13g2_fill_1 FILLER_0_94_455 ();
 sg13g2_fill_1 FILLER_0_94_470 ();
 sg13g2_fill_8 FILLER_0_94_510 ();
 sg13g2_fill_8 FILLER_0_94_518 ();
 sg13g2_fill_8 FILLER_0_94_526 ();
 sg13g2_fill_4 FILLER_0_94_534 ();
 sg13g2_fill_2 FILLER_0_94_554 ();
 sg13g2_fill_1 FILLER_0_94_556 ();
 sg13g2_fill_2 FILLER_0_94_587 ();
 sg13g2_fill_1 FILLER_0_94_589 ();
 sg13g2_fill_8 FILLER_0_94_672 ();
 sg13g2_fill_4 FILLER_0_94_680 ();
 sg13g2_fill_1 FILLER_0_94_684 ();
 sg13g2_fill_1 FILLER_0_94_704 ();
 sg13g2_fill_2 FILLER_0_94_729 ();
 sg13g2_fill_1 FILLER_0_94_731 ();
 sg13g2_fill_8 FILLER_0_94_748 ();
 sg13g2_fill_4 FILLER_0_94_756 ();
 sg13g2_fill_2 FILLER_0_94_760 ();
 sg13g2_fill_2 FILLER_0_94_767 ();
 sg13g2_fill_8 FILLER_0_94_773 ();
 sg13g2_fill_1 FILLER_0_94_781 ();
 sg13g2_fill_8 FILLER_0_94_786 ();
 sg13g2_fill_4 FILLER_0_94_794 ();
 sg13g2_fill_1 FILLER_0_94_798 ();
 sg13g2_fill_8 FILLER_0_94_803 ();
 sg13g2_fill_8 FILLER_0_94_811 ();
 sg13g2_fill_8 FILLER_0_94_819 ();
 sg13g2_fill_8 FILLER_0_94_827 ();
 sg13g2_fill_1 FILLER_0_94_835 ();
 sg13g2_fill_4 FILLER_0_94_846 ();
 sg13g2_fill_4 FILLER_0_94_885 ();
 sg13g2_fill_2 FILLER_0_94_895 ();
 sg13g2_fill_4 FILLER_0_94_901 ();
 sg13g2_fill_1 FILLER_0_94_910 ();
 sg13g2_fill_1 FILLER_0_94_916 ();
 sg13g2_fill_8 FILLER_0_94_951 ();
 sg13g2_fill_1 FILLER_0_94_959 ();
 sg13g2_fill_1 FILLER_0_94_965 ();
 sg13g2_fill_8 FILLER_0_94_1000 ();
 sg13g2_fill_2 FILLER_0_94_1008 ();
 sg13g2_fill_1 FILLER_0_94_1010 ();
 sg13g2_fill_1 FILLER_0_94_1015 ();
 sg13g2_fill_1 FILLER_0_94_1046 ();
 sg13g2_fill_2 FILLER_0_94_1068 ();
 sg13g2_fill_2 FILLER_0_94_1081 ();
 sg13g2_fill_8 FILLER_0_94_1109 ();
 sg13g2_fill_8 FILLER_0_94_1117 ();
 sg13g2_fill_8 FILLER_0_94_1125 ();
 sg13g2_fill_8 FILLER_0_94_1133 ();
 sg13g2_fill_8 FILLER_0_94_1141 ();
 sg13g2_fill_8 FILLER_0_94_1149 ();
 sg13g2_fill_8 FILLER_0_94_1157 ();
 sg13g2_fill_8 FILLER_0_94_1165 ();
 sg13g2_fill_8 FILLER_0_94_1173 ();
 sg13g2_fill_8 FILLER_0_94_1181 ();
 sg13g2_fill_8 FILLER_0_94_1189 ();
 sg13g2_fill_8 FILLER_0_94_1197 ();
 sg13g2_fill_8 FILLER_0_94_1205 ();
 sg13g2_fill_8 FILLER_0_94_1213 ();
 sg13g2_decap_8 FILLER_0_94_1221 ();
 sg13g2_fill_8 FILLER_0_95_0 ();
 sg13g2_fill_2 FILLER_0_95_8 ();
 sg13g2_fill_2 FILLER_0_95_66 ();
 sg13g2_fill_1 FILLER_0_95_68 ();
 sg13g2_fill_2 FILLER_0_95_95 ();
 sg13g2_fill_2 FILLER_0_95_101 ();
 sg13g2_fill_1 FILLER_0_95_129 ();
 sg13g2_fill_2 FILLER_0_95_134 ();
 sg13g2_fill_1 FILLER_0_95_140 ();
 sg13g2_fill_2 FILLER_0_95_167 ();
 sg13g2_fill_8 FILLER_0_95_195 ();
 sg13g2_fill_8 FILLER_0_95_203 ();
 sg13g2_fill_8 FILLER_0_95_211 ();
 sg13g2_fill_8 FILLER_0_95_219 ();
 sg13g2_fill_8 FILLER_0_95_227 ();
 sg13g2_fill_8 FILLER_0_95_235 ();
 sg13g2_fill_8 FILLER_0_95_243 ();
 sg13g2_fill_2 FILLER_0_95_274 ();
 sg13g2_fill_8 FILLER_0_95_285 ();
 sg13g2_fill_8 FILLER_0_95_293 ();
 sg13g2_fill_4 FILLER_0_95_301 ();
 sg13g2_fill_1 FILLER_0_95_320 ();
 sg13g2_fill_8 FILLER_0_95_325 ();
 sg13g2_fill_8 FILLER_0_95_333 ();
 sg13g2_fill_8 FILLER_0_95_341 ();
 sg13g2_fill_2 FILLER_0_95_349 ();
 sg13g2_fill_1 FILLER_0_95_351 ();
 sg13g2_fill_4 FILLER_0_95_372 ();
 sg13g2_fill_1 FILLER_0_95_376 ();
 sg13g2_fill_1 FILLER_0_95_392 ();
 sg13g2_fill_8 FILLER_0_95_397 ();
 sg13g2_fill_1 FILLER_0_95_405 ();
 sg13g2_fill_4 FILLER_0_95_415 ();
 sg13g2_fill_8 FILLER_0_95_433 ();
 sg13g2_fill_2 FILLER_0_95_441 ();
 sg13g2_fill_8 FILLER_0_95_447 ();
 sg13g2_fill_4 FILLER_0_95_455 ();
 sg13g2_fill_2 FILLER_0_95_459 ();
 sg13g2_fill_4 FILLER_0_95_471 ();
 sg13g2_fill_8 FILLER_0_95_499 ();
 sg13g2_fill_1 FILLER_0_95_507 ();
 sg13g2_fill_4 FILLER_0_95_512 ();
 sg13g2_fill_4 FILLER_0_95_530 ();
 sg13g2_fill_8 FILLER_0_95_575 ();
 sg13g2_fill_4 FILLER_0_95_583 ();
 sg13g2_fill_2 FILLER_0_95_587 ();
 sg13g2_fill_2 FILLER_0_95_593 ();
 sg13g2_fill_1 FILLER_0_95_595 ();
 sg13g2_fill_4 FILLER_0_95_600 ();
 sg13g2_fill_2 FILLER_0_95_604 ();
 sg13g2_decap_8 FILLER_0_95_616 ();
 sg13g2_fill_1 FILLER_0_95_627 ();
 sg13g2_fill_2 FILLER_0_95_633 ();
 sg13g2_fill_2 FILLER_0_95_652 ();
 sg13g2_fill_8 FILLER_0_95_658 ();
 sg13g2_fill_8 FILLER_0_95_666 ();
 sg13g2_fill_8 FILLER_0_95_674 ();
 sg13g2_fill_4 FILLER_0_95_682 ();
 sg13g2_fill_1 FILLER_0_95_712 ();
 sg13g2_fill_2 FILLER_0_95_718 ();
 sg13g2_fill_2 FILLER_0_95_746 ();
 sg13g2_fill_2 FILLER_0_95_774 ();
 sg13g2_fill_1 FILLER_0_95_776 ();
 sg13g2_fill_2 FILLER_0_95_792 ();
 sg13g2_fill_8 FILLER_0_95_798 ();
 sg13g2_fill_2 FILLER_0_95_818 ();
 sg13g2_fill_1 FILLER_0_95_820 ();
 sg13g2_fill_2 FILLER_0_95_852 ();
 sg13g2_fill_1 FILLER_0_95_854 ();
 sg13g2_fill_1 FILLER_0_95_876 ();
 sg13g2_fill_2 FILLER_0_95_891 ();
 sg13g2_fill_2 FILLER_0_95_916 ();
 sg13g2_fill_2 FILLER_0_95_922 ();
 sg13g2_fill_1 FILLER_0_95_924 ();
 sg13g2_fill_4 FILLER_0_95_932 ();
 sg13g2_fill_2 FILLER_0_95_936 ();
 sg13g2_fill_8 FILLER_0_95_948 ();
 sg13g2_fill_4 FILLER_0_95_956 ();
 sg13g2_fill_2 FILLER_0_95_960 ();
 sg13g2_fill_2 FILLER_0_95_972 ();
 sg13g2_fill_2 FILLER_0_95_979 ();
 sg13g2_fill_4 FILLER_0_95_996 ();
 sg13g2_fill_2 FILLER_0_95_1000 ();
 sg13g2_fill_1 FILLER_0_95_1037 ();
 sg13g2_fill_2 FILLER_0_95_1043 ();
 sg13g2_fill_2 FILLER_0_95_1067 ();
 sg13g2_fill_1 FILLER_0_95_1082 ();
 sg13g2_fill_2 FILLER_0_95_1087 ();
 sg13g2_fill_1 FILLER_0_95_1089 ();
 sg13g2_fill_8 FILLER_0_95_1116 ();
 sg13g2_fill_8 FILLER_0_95_1124 ();
 sg13g2_fill_8 FILLER_0_95_1132 ();
 sg13g2_fill_8 FILLER_0_95_1140 ();
 sg13g2_fill_8 FILLER_0_95_1148 ();
 sg13g2_fill_8 FILLER_0_95_1156 ();
 sg13g2_fill_8 FILLER_0_95_1164 ();
 sg13g2_fill_8 FILLER_0_95_1172 ();
 sg13g2_fill_8 FILLER_0_95_1180 ();
 sg13g2_fill_8 FILLER_0_95_1188 ();
 sg13g2_fill_8 FILLER_0_95_1196 ();
 sg13g2_fill_8 FILLER_0_95_1204 ();
 sg13g2_fill_8 FILLER_0_95_1212 ();
 sg13g2_fill_8 FILLER_0_95_1220 ();
 sg13g2_fill_1 FILLER_0_96_0 ();
 sg13g2_fill_2 FILLER_0_96_27 ();
 sg13g2_fill_8 FILLER_0_96_85 ();
 sg13g2_fill_8 FILLER_0_96_93 ();
 sg13g2_fill_8 FILLER_0_96_101 ();
 sg13g2_fill_2 FILLER_0_96_109 ();
 sg13g2_fill_1 FILLER_0_96_111 ();
 sg13g2_fill_8 FILLER_0_96_116 ();
 sg13g2_fill_8 FILLER_0_96_124 ();
 sg13g2_fill_2 FILLER_0_96_132 ();
 sg13g2_fill_1 FILLER_0_96_134 ();
 sg13g2_fill_1 FILLER_0_96_144 ();
 sg13g2_fill_8 FILLER_0_96_155 ();
 sg13g2_fill_8 FILLER_0_96_163 ();
 sg13g2_fill_4 FILLER_0_96_171 ();
 sg13g2_fill_2 FILLER_0_96_184 ();
 sg13g2_fill_4 FILLER_0_96_206 ();
 sg13g2_fill_8 FILLER_0_96_236 ();
 sg13g2_fill_1 FILLER_0_96_248 ();
 sg13g2_fill_8 FILLER_0_96_275 ();
 sg13g2_fill_8 FILLER_0_96_283 ();
 sg13g2_fill_8 FILLER_0_96_291 ();
 sg13g2_fill_1 FILLER_0_96_299 ();
 sg13g2_fill_8 FILLER_0_96_319 ();
 sg13g2_decap_8 FILLER_0_96_327 ();
 sg13g2_fill_1 FILLER_0_96_370 ();
 sg13g2_fill_8 FILLER_0_96_376 ();
 sg13g2_fill_2 FILLER_0_96_384 ();
 sg13g2_fill_1 FILLER_0_96_412 ();
 sg13g2_decap_8 FILLER_0_96_472 ();
 sg13g2_fill_2 FILLER_0_96_536 ();
 sg13g2_fill_1 FILLER_0_96_538 ();
 sg13g2_fill_4 FILLER_0_96_575 ();
 sg13g2_fill_1 FILLER_0_96_579 ();
 sg13g2_fill_4 FILLER_0_96_606 ();
 sg13g2_fill_2 FILLER_0_96_610 ();
 sg13g2_fill_8 FILLER_0_96_617 ();
 sg13g2_fill_8 FILLER_0_96_625 ();
 sg13g2_fill_4 FILLER_0_96_633 ();
 sg13g2_fill_2 FILLER_0_96_637 ();
 sg13g2_fill_4 FILLER_0_96_669 ();
 sg13g2_fill_2 FILLER_0_96_673 ();
 sg13g2_fill_4 FILLER_0_96_706 ();
 sg13g2_fill_1 FILLER_0_96_710 ();
 sg13g2_fill_2 FILLER_0_96_749 ();
 sg13g2_fill_1 FILLER_0_96_751 ();
 sg13g2_fill_2 FILLER_0_96_786 ();
 sg13g2_fill_1 FILLER_0_96_788 ();
 sg13g2_fill_2 FILLER_0_96_798 ();
 sg13g2_fill_2 FILLER_0_96_810 ();
 sg13g2_fill_1 FILLER_0_96_812 ();
 sg13g2_fill_1 FILLER_0_96_823 ();
 sg13g2_fill_1 FILLER_0_96_859 ();
 sg13g2_fill_1 FILLER_0_96_865 ();
 sg13g2_fill_8 FILLER_0_96_882 ();
 sg13g2_fill_8 FILLER_0_96_890 ();
 sg13g2_fill_1 FILLER_0_96_898 ();
 sg13g2_fill_2 FILLER_0_96_908 ();
 sg13g2_fill_1 FILLER_0_96_910 ();
 sg13g2_fill_8 FILLER_0_96_916 ();
 sg13g2_fill_8 FILLER_0_96_924 ();
 sg13g2_fill_8 FILLER_0_96_932 ();
 sg13g2_fill_2 FILLER_0_96_940 ();
 sg13g2_fill_1 FILLER_0_96_968 ();
 sg13g2_fill_2 FILLER_0_96_976 ();
 sg13g2_fill_2 FILLER_0_96_988 ();
 sg13g2_fill_1 FILLER_0_96_994 ();
 sg13g2_fill_8 FILLER_0_96_1052 ();
 sg13g2_fill_2 FILLER_0_96_1060 ();
 sg13g2_fill_1 FILLER_0_96_1066 ();
 sg13g2_fill_8 FILLER_0_96_1071 ();
 sg13g2_fill_8 FILLER_0_96_1079 ();
 sg13g2_fill_1 FILLER_0_96_1087 ();
 sg13g2_fill_2 FILLER_0_96_1096 ();
 sg13g2_fill_8 FILLER_0_96_1102 ();
 sg13g2_fill_8 FILLER_0_96_1110 ();
 sg13g2_fill_8 FILLER_0_96_1118 ();
 sg13g2_fill_8 FILLER_0_96_1126 ();
 sg13g2_fill_8 FILLER_0_96_1134 ();
 sg13g2_fill_8 FILLER_0_96_1142 ();
 sg13g2_fill_8 FILLER_0_96_1150 ();
 sg13g2_fill_8 FILLER_0_96_1158 ();
 sg13g2_fill_8 FILLER_0_96_1166 ();
 sg13g2_fill_8 FILLER_0_96_1174 ();
 sg13g2_fill_8 FILLER_0_96_1182 ();
 sg13g2_fill_8 FILLER_0_96_1190 ();
 sg13g2_fill_8 FILLER_0_96_1198 ();
 sg13g2_fill_8 FILLER_0_96_1206 ();
 sg13g2_fill_8 FILLER_0_96_1214 ();
 sg13g2_fill_4 FILLER_0_96_1222 ();
 sg13g2_fill_2 FILLER_0_96_1226 ();
 sg13g2_fill_8 FILLER_0_97_0 ();
 sg13g2_fill_4 FILLER_0_97_55 ();
 sg13g2_fill_2 FILLER_0_97_59 ();
 sg13g2_fill_8 FILLER_0_97_65 ();
 sg13g2_fill_4 FILLER_0_97_73 ();
 sg13g2_fill_2 FILLER_0_97_77 ();
 sg13g2_fill_8 FILLER_0_97_83 ();
 sg13g2_fill_8 FILLER_0_97_95 ();
 sg13g2_fill_8 FILLER_0_97_103 ();
 sg13g2_fill_2 FILLER_0_97_111 ();
 sg13g2_fill_1 FILLER_0_97_113 ();
 sg13g2_fill_1 FILLER_0_97_119 ();
 sg13g2_fill_8 FILLER_0_97_124 ();
 sg13g2_fill_4 FILLER_0_97_145 ();
 sg13g2_fill_2 FILLER_0_97_149 ();
 sg13g2_fill_8 FILLER_0_97_155 ();
 sg13g2_fill_4 FILLER_0_97_163 ();
 sg13g2_fill_2 FILLER_0_97_167 ();
 sg13g2_fill_8 FILLER_0_97_173 ();
 sg13g2_fill_2 FILLER_0_97_181 ();
 sg13g2_fill_1 FILLER_0_97_193 ();
 sg13g2_fill_1 FILLER_0_97_204 ();
 sg13g2_fill_1 FILLER_0_97_262 ();
 sg13g2_fill_4 FILLER_0_97_268 ();
 sg13g2_fill_1 FILLER_0_97_272 ();
 sg13g2_fill_8 FILLER_0_97_283 ();
 sg13g2_decap_8 FILLER_0_97_291 ();
 sg13g2_fill_2 FILLER_0_97_329 ();
 sg13g2_fill_1 FILLER_0_97_331 ();
 sg13g2_fill_2 FILLER_0_97_358 ();
 sg13g2_fill_1 FILLER_0_97_360 ();
 sg13g2_fill_1 FILLER_0_97_397 ();
 sg13g2_fill_1 FILLER_0_97_406 ();
 sg13g2_fill_1 FILLER_0_97_433 ();
 sg13g2_fill_2 FILLER_0_97_485 ();
 sg13g2_fill_8 FILLER_0_97_497 ();
 sg13g2_fill_8 FILLER_0_97_505 ();
 sg13g2_fill_4 FILLER_0_97_522 ();
 sg13g2_fill_2 FILLER_0_97_526 ();
 sg13g2_fill_8 FILLER_0_97_536 ();
 sg13g2_fill_4 FILLER_0_97_553 ();
 sg13g2_fill_1 FILLER_0_97_562 ();
 sg13g2_fill_2 FILLER_0_97_573 ();
 sg13g2_fill_8 FILLER_0_97_579 ();
 sg13g2_fill_4 FILLER_0_97_595 ();
 sg13g2_fill_1 FILLER_0_97_608 ();
 sg13g2_fill_8 FILLER_0_97_624 ();
 sg13g2_fill_2 FILLER_0_97_632 ();
 sg13g2_fill_2 FILLER_0_97_644 ();
 sg13g2_fill_2 FILLER_0_97_651 ();
 sg13g2_fill_1 FILLER_0_97_653 ();
 sg13g2_fill_2 FILLER_0_97_688 ();
 sg13g2_fill_1 FILLER_0_97_694 ();
 sg13g2_fill_4 FILLER_0_97_705 ();
 sg13g2_decap_8 FILLER_0_97_734 ();
 sg13g2_fill_2 FILLER_0_97_753 ();
 sg13g2_fill_2 FILLER_0_97_774 ();
 sg13g2_fill_4 FILLER_0_97_780 ();
 sg13g2_fill_2 FILLER_0_97_788 ();
 sg13g2_fill_1 FILLER_0_97_820 ();
 sg13g2_fill_2 FILLER_0_97_826 ();
 sg13g2_fill_8 FILLER_0_97_854 ();
 sg13g2_fill_4 FILLER_0_97_862 ();
 sg13g2_fill_4 FILLER_0_97_871 ();
 sg13g2_fill_1 FILLER_0_97_939 ();
 sg13g2_fill_2 FILLER_0_97_1006 ();
 sg13g2_decap_8 FILLER_0_97_1012 ();
 sg13g2_fill_1 FILLER_0_97_1024 ();
 sg13g2_fill_2 FILLER_0_97_1030 ();
 sg13g2_fill_1 FILLER_0_97_1032 ();
 sg13g2_fill_4 FILLER_0_97_1037 ();
 sg13g2_fill_2 FILLER_0_97_1041 ();
 sg13g2_fill_2 FILLER_0_97_1048 ();
 sg13g2_fill_1 FILLER_0_97_1050 ();
 sg13g2_fill_2 FILLER_0_97_1056 ();
 sg13g2_fill_1 FILLER_0_97_1058 ();
 sg13g2_fill_2 FILLER_0_97_1085 ();
 sg13g2_fill_1 FILLER_0_97_1092 ();
 sg13g2_fill_8 FILLER_0_97_1102 ();
 sg13g2_fill_8 FILLER_0_97_1110 ();
 sg13g2_fill_8 FILLER_0_97_1118 ();
 sg13g2_fill_8 FILLER_0_97_1126 ();
 sg13g2_fill_8 FILLER_0_97_1134 ();
 sg13g2_fill_8 FILLER_0_97_1142 ();
 sg13g2_fill_8 FILLER_0_97_1150 ();
 sg13g2_fill_8 FILLER_0_97_1158 ();
 sg13g2_fill_8 FILLER_0_97_1166 ();
 sg13g2_fill_8 FILLER_0_97_1174 ();
 sg13g2_fill_8 FILLER_0_97_1182 ();
 sg13g2_fill_8 FILLER_0_97_1190 ();
 sg13g2_fill_8 FILLER_0_97_1198 ();
 sg13g2_fill_8 FILLER_0_97_1206 ();
 sg13g2_fill_8 FILLER_0_97_1214 ();
 sg13g2_fill_4 FILLER_0_97_1222 ();
 sg13g2_fill_2 FILLER_0_97_1226 ();
 sg13g2_fill_8 FILLER_0_98_0 ();
 sg13g2_fill_8 FILLER_0_98_8 ();
 sg13g2_fill_8 FILLER_0_98_16 ();
 sg13g2_fill_8 FILLER_0_98_24 ();
 sg13g2_fill_2 FILLER_0_98_32 ();
 sg13g2_fill_1 FILLER_0_98_34 ();
 sg13g2_fill_8 FILLER_0_98_39 ();
 sg13g2_fill_8 FILLER_0_98_47 ();
 sg13g2_fill_8 FILLER_0_98_55 ();
 sg13g2_decap_8 FILLER_0_98_63 ();
 sg13g2_fill_2 FILLER_0_98_110 ();
 sg13g2_fill_1 FILLER_0_98_112 ();
 sg13g2_fill_2 FILLER_0_98_139 ();
 sg13g2_fill_2 FILLER_0_98_167 ();
 sg13g2_fill_4 FILLER_0_98_195 ();
 sg13g2_fill_2 FILLER_0_98_204 ();
 sg13g2_fill_4 FILLER_0_98_215 ();
 sg13g2_fill_1 FILLER_0_98_219 ();
 sg13g2_fill_8 FILLER_0_98_224 ();
 sg13g2_fill_2 FILLER_0_98_232 ();
 sg13g2_fill_1 FILLER_0_98_234 ();
 sg13g2_fill_8 FILLER_0_98_239 ();
 sg13g2_decap_8 FILLER_0_98_247 ();
 sg13g2_fill_2 FILLER_0_98_258 ();
 sg13g2_fill_1 FILLER_0_98_260 ();
 sg13g2_fill_2 FILLER_0_98_287 ();
 sg13g2_fill_1 FILLER_0_98_338 ();
 sg13g2_fill_1 FILLER_0_98_369 ();
 sg13g2_fill_8 FILLER_0_98_389 ();
 sg13g2_fill_4 FILLER_0_98_397 ();
 sg13g2_fill_2 FILLER_0_98_401 ();
 sg13g2_fill_4 FILLER_0_98_411 ();
 sg13g2_fill_8 FILLER_0_98_419 ();
 sg13g2_fill_2 FILLER_0_98_427 ();
 sg13g2_fill_1 FILLER_0_98_429 ();
 sg13g2_fill_1 FILLER_0_98_469 ();
 sg13g2_fill_8 FILLER_0_98_531 ();
 sg13g2_fill_8 FILLER_0_98_539 ();
 sg13g2_fill_2 FILLER_0_98_547 ();
 sg13g2_fill_1 FILLER_0_98_564 ();
 sg13g2_fill_1 FILLER_0_98_591 ();
 sg13g2_fill_1 FILLER_0_98_618 ();
 sg13g2_fill_2 FILLER_0_98_645 ();
 sg13g2_fill_1 FILLER_0_98_657 ();
 sg13g2_fill_4 FILLER_0_98_675 ();
 sg13g2_fill_2 FILLER_0_98_709 ();
 sg13g2_fill_2 FILLER_0_98_715 ();
 sg13g2_fill_2 FILLER_0_98_722 ();
 sg13g2_fill_1 FILLER_0_98_724 ();
 sg13g2_fill_2 FILLER_0_98_730 ();
 sg13g2_fill_1 FILLER_0_98_732 ();
 sg13g2_fill_2 FILLER_0_98_737 ();
 sg13g2_fill_1 FILLER_0_98_739 ();
 sg13g2_fill_8 FILLER_0_98_750 ();
 sg13g2_fill_8 FILLER_0_98_758 ();
 sg13g2_fill_4 FILLER_0_98_766 ();
 sg13g2_fill_1 FILLER_0_98_770 ();
 sg13g2_fill_2 FILLER_0_98_775 ();
 sg13g2_fill_8 FILLER_0_98_789 ();
 sg13g2_fill_2 FILLER_0_98_797 ();
 sg13g2_fill_1 FILLER_0_98_799 ();
 sg13g2_fill_2 FILLER_0_98_804 ();
 sg13g2_fill_1 FILLER_0_98_806 ();
 sg13g2_fill_1 FILLER_0_98_812 ();
 sg13g2_fill_2 FILLER_0_98_842 ();
 sg13g2_fill_8 FILLER_0_98_848 ();
 sg13g2_fill_4 FILLER_0_98_856 ();
 sg13g2_fill_8 FILLER_0_98_895 ();
 sg13g2_decap_8 FILLER_0_98_903 ();
 sg13g2_fill_8 FILLER_0_98_926 ();
 sg13g2_fill_4 FILLER_0_98_934 ();
 sg13g2_fill_1 FILLER_0_98_938 ();
 sg13g2_fill_1 FILLER_0_98_970 ();
 sg13g2_fill_2 FILLER_0_98_975 ();
 sg13g2_fill_2 FILLER_0_98_982 ();
 sg13g2_fill_2 FILLER_0_98_988 ();
 sg13g2_fill_1 FILLER_0_98_990 ();
 sg13g2_decap_8 FILLER_0_98_1001 ();
 sg13g2_fill_2 FILLER_0_98_1013 ();
 sg13g2_fill_2 FILLER_0_98_1019 ();
 sg13g2_fill_1 FILLER_0_98_1035 ();
 sg13g2_fill_1 FILLER_0_98_1073 ();
 sg13g2_fill_1 FILLER_0_98_1083 ();
 sg13g2_fill_8 FILLER_0_98_1110 ();
 sg13g2_fill_8 FILLER_0_98_1118 ();
 sg13g2_fill_8 FILLER_0_98_1126 ();
 sg13g2_fill_8 FILLER_0_98_1134 ();
 sg13g2_fill_8 FILLER_0_98_1142 ();
 sg13g2_fill_8 FILLER_0_98_1150 ();
 sg13g2_fill_8 FILLER_0_98_1158 ();
 sg13g2_fill_8 FILLER_0_98_1166 ();
 sg13g2_fill_8 FILLER_0_98_1174 ();
 sg13g2_fill_8 FILLER_0_98_1182 ();
 sg13g2_fill_8 FILLER_0_98_1190 ();
 sg13g2_fill_8 FILLER_0_98_1198 ();
 sg13g2_fill_8 FILLER_0_98_1206 ();
 sg13g2_fill_8 FILLER_0_98_1214 ();
 sg13g2_fill_4 FILLER_0_98_1222 ();
 sg13g2_fill_2 FILLER_0_98_1226 ();
 sg13g2_fill_8 FILLER_0_99_0 ();
 sg13g2_fill_8 FILLER_0_99_8 ();
 sg13g2_fill_1 FILLER_0_99_16 ();
 sg13g2_fill_4 FILLER_0_99_47 ();
 sg13g2_fill_1 FILLER_0_99_51 ();
 sg13g2_fill_2 FILLER_0_99_98 ();
 sg13g2_fill_4 FILLER_0_99_136 ();
 sg13g2_fill_2 FILLER_0_99_170 ();
 sg13g2_fill_2 FILLER_0_99_177 ();
 sg13g2_fill_1 FILLER_0_99_179 ();
 sg13g2_fill_2 FILLER_0_99_206 ();
 sg13g2_fill_1 FILLER_0_99_208 ();
 sg13g2_fill_8 FILLER_0_99_235 ();
 sg13g2_fill_4 FILLER_0_99_243 ();
 sg13g2_fill_1 FILLER_0_99_247 ();
 sg13g2_fill_2 FILLER_0_99_263 ();
 sg13g2_fill_4 FILLER_0_99_269 ();
 sg13g2_fill_8 FILLER_0_99_283 ();
 sg13g2_fill_4 FILLER_0_99_291 ();
 sg13g2_fill_2 FILLER_0_99_299 ();
 sg13g2_fill_1 FILLER_0_99_301 ();
 sg13g2_fill_8 FILLER_0_99_328 ();
 sg13g2_fill_8 FILLER_0_99_336 ();
 sg13g2_fill_1 FILLER_0_99_344 ();
 sg13g2_fill_1 FILLER_0_99_360 ();
 sg13g2_fill_4 FILLER_0_99_418 ();
 sg13g2_fill_2 FILLER_0_99_422 ();
 sg13g2_fill_8 FILLER_0_99_437 ();
 sg13g2_fill_4 FILLER_0_99_445 ();
 sg13g2_fill_1 FILLER_0_99_449 ();
 sg13g2_fill_4 FILLER_0_99_454 ();
 sg13g2_fill_1 FILLER_0_99_458 ();
 sg13g2_fill_1 FILLER_0_99_467 ();
 sg13g2_fill_1 FILLER_0_99_499 ();
 sg13g2_fill_4 FILLER_0_99_519 ();
 sg13g2_fill_8 FILLER_0_99_540 ();
 sg13g2_fill_8 FILLER_0_99_548 ();
 sg13g2_fill_2 FILLER_0_99_556 ();
 sg13g2_fill_1 FILLER_0_99_598 ();
 sg13g2_fill_1 FILLER_0_99_625 ();
 sg13g2_fill_1 FILLER_0_99_630 ();
 sg13g2_fill_2 FILLER_0_99_641 ();
 sg13g2_fill_2 FILLER_0_99_661 ();
 sg13g2_fill_8 FILLER_0_99_667 ();
 sg13g2_fill_8 FILLER_0_99_675 ();
 sg13g2_fill_4 FILLER_0_99_683 ();
 sg13g2_fill_2 FILLER_0_99_687 ();
 sg13g2_fill_8 FILLER_0_99_697 ();
 sg13g2_fill_2 FILLER_0_99_709 ();
 sg13g2_fill_2 FILLER_0_99_721 ();
 sg13g2_fill_1 FILLER_0_99_723 ();
 sg13g2_fill_1 FILLER_0_99_776 ();
 sg13g2_fill_8 FILLER_0_99_803 ();
 sg13g2_fill_8 FILLER_0_99_816 ();
 sg13g2_fill_8 FILLER_0_99_824 ();
 sg13g2_fill_8 FILLER_0_99_832 ();
 sg13g2_fill_8 FILLER_0_99_840 ();
 sg13g2_fill_8 FILLER_0_99_848 ();
 sg13g2_fill_8 FILLER_0_99_856 ();
 sg13g2_fill_4 FILLER_0_99_864 ();
 sg13g2_fill_1 FILLER_0_99_868 ();
 sg13g2_fill_2 FILLER_0_99_914 ();
 sg13g2_fill_1 FILLER_0_99_916 ();
 sg13g2_fill_8 FILLER_0_99_924 ();
 sg13g2_fill_2 FILLER_0_99_932 ();
 sg13g2_decap_8 FILLER_0_99_938 ();
 sg13g2_fill_8 FILLER_0_99_950 ();
 sg13g2_decap_8 FILLER_0_99_989 ();
 sg13g2_fill_1 FILLER_0_99_1005 ();
 sg13g2_fill_1 FILLER_0_99_1042 ();
 sg13g2_fill_8 FILLER_0_99_1103 ();
 sg13g2_fill_8 FILLER_0_99_1111 ();
 sg13g2_fill_8 FILLER_0_99_1119 ();
 sg13g2_fill_8 FILLER_0_99_1127 ();
 sg13g2_fill_8 FILLER_0_99_1135 ();
 sg13g2_fill_8 FILLER_0_99_1143 ();
 sg13g2_fill_8 FILLER_0_99_1151 ();
 sg13g2_fill_8 FILLER_0_99_1159 ();
 sg13g2_fill_8 FILLER_0_99_1167 ();
 sg13g2_fill_8 FILLER_0_99_1175 ();
 sg13g2_fill_8 FILLER_0_99_1183 ();
 sg13g2_fill_8 FILLER_0_99_1191 ();
 sg13g2_fill_8 FILLER_0_99_1199 ();
 sg13g2_fill_8 FILLER_0_99_1207 ();
 sg13g2_fill_8 FILLER_0_99_1215 ();
 sg13g2_fill_4 FILLER_0_99_1223 ();
 sg13g2_fill_1 FILLER_0_99_1227 ();
 sg13g2_decap_8 FILLER_0_100_0 ();
 sg13g2_fill_4 FILLER_0_100_11 ();
 sg13g2_fill_1 FILLER_0_100_15 ();
 sg13g2_decap_8 FILLER_0_100_21 ();
 sg13g2_fill_2 FILLER_0_100_55 ();
 sg13g2_fill_2 FILLER_0_100_135 ();
 sg13g2_fill_1 FILLER_0_100_137 ();
 sg13g2_fill_1 FILLER_0_100_196 ();
 sg13g2_fill_8 FILLER_0_100_202 ();
 sg13g2_fill_4 FILLER_0_100_210 ();
 sg13g2_fill_1 FILLER_0_100_214 ();
 sg13g2_fill_1 FILLER_0_100_219 ();
 sg13g2_fill_8 FILLER_0_100_229 ();
 sg13g2_fill_8 FILLER_0_100_237 ();
 sg13g2_fill_8 FILLER_0_100_245 ();
 sg13g2_fill_4 FILLER_0_100_253 ();
 sg13g2_fill_1 FILLER_0_100_257 ();
 sg13g2_fill_8 FILLER_0_100_284 ();
 sg13g2_decap_8 FILLER_0_100_292 ();
 sg13g2_fill_2 FILLER_0_100_312 ();
 sg13g2_fill_8 FILLER_0_100_328 ();
 sg13g2_fill_8 FILLER_0_100_336 ();
 sg13g2_fill_4 FILLER_0_100_344 ();
 sg13g2_fill_2 FILLER_0_100_348 ();
 sg13g2_fill_2 FILLER_0_100_354 ();
 sg13g2_fill_4 FILLER_0_100_361 ();
 sg13g2_fill_1 FILLER_0_100_365 ();
 sg13g2_fill_8 FILLER_0_100_451 ();
 sg13g2_fill_8 FILLER_0_100_459 ();
 sg13g2_fill_4 FILLER_0_100_467 ();
 sg13g2_fill_1 FILLER_0_100_471 ();
 sg13g2_fill_8 FILLER_0_100_486 ();
 sg13g2_fill_2 FILLER_0_100_494 ();
 sg13g2_fill_1 FILLER_0_100_496 ();
 sg13g2_fill_4 FILLER_0_100_501 ();
 sg13g2_fill_2 FILLER_0_100_505 ();
 sg13g2_fill_2 FILLER_0_100_552 ();
 sg13g2_fill_1 FILLER_0_100_554 ();
 sg13g2_fill_2 FILLER_0_100_560 ();
 sg13g2_fill_1 FILLER_0_100_562 ();
 sg13g2_fill_2 FILLER_0_100_583 ();
 sg13g2_fill_1 FILLER_0_100_585 ();
 sg13g2_fill_8 FILLER_0_100_590 ();
 sg13g2_fill_2 FILLER_0_100_598 ();
 sg13g2_fill_4 FILLER_0_100_641 ();
 sg13g2_fill_2 FILLER_0_100_645 ();
 sg13g2_fill_8 FILLER_0_100_678 ();
 sg13g2_fill_2 FILLER_0_100_686 ();
 sg13g2_fill_1 FILLER_0_100_688 ();
 sg13g2_fill_1 FILLER_0_100_720 ();
 sg13g2_fill_1 FILLER_0_100_747 ();
 sg13g2_fill_4 FILLER_0_100_762 ();
 sg13g2_fill_2 FILLER_0_100_771 ();
 sg13g2_fill_8 FILLER_0_100_777 ();
 sg13g2_fill_8 FILLER_0_100_785 ();
 sg13g2_fill_4 FILLER_0_100_793 ();
 sg13g2_fill_1 FILLER_0_100_797 ();
 sg13g2_fill_8 FILLER_0_100_839 ();
 sg13g2_fill_2 FILLER_0_100_851 ();
 sg13g2_fill_1 FILLER_0_100_892 ();
 sg13g2_fill_1 FILLER_0_100_898 ();
 sg13g2_fill_1 FILLER_0_100_904 ();
 sg13g2_fill_2 FILLER_0_100_909 ();
 sg13g2_fill_1 FILLER_0_100_921 ();
 sg13g2_fill_8 FILLER_0_100_963 ();
 sg13g2_fill_8 FILLER_0_100_971 ();
 sg13g2_decap_8 FILLER_0_100_979 ();
 sg13g2_fill_1 FILLER_0_100_999 ();
 sg13g2_fill_8 FILLER_0_100_1014 ();
 sg13g2_fill_4 FILLER_0_100_1026 ();
 sg13g2_fill_1 FILLER_0_100_1044 ();
 sg13g2_fill_2 FILLER_0_100_1058 ();
 sg13g2_fill_1 FILLER_0_100_1064 ();
 sg13g2_fill_8 FILLER_0_100_1075 ();
 sg13g2_fill_2 FILLER_0_100_1096 ();
 sg13g2_fill_1 FILLER_0_100_1102 ();
 sg13g2_fill_8 FILLER_0_100_1108 ();
 sg13g2_fill_8 FILLER_0_100_1116 ();
 sg13g2_fill_8 FILLER_0_100_1132 ();
 sg13g2_fill_8 FILLER_0_100_1140 ();
 sg13g2_fill_8 FILLER_0_100_1148 ();
 sg13g2_fill_8 FILLER_0_100_1156 ();
 sg13g2_fill_8 FILLER_0_100_1164 ();
 sg13g2_fill_8 FILLER_0_100_1172 ();
 sg13g2_fill_8 FILLER_0_100_1180 ();
 sg13g2_fill_8 FILLER_0_100_1188 ();
 sg13g2_fill_8 FILLER_0_100_1196 ();
 sg13g2_fill_8 FILLER_0_100_1204 ();
 sg13g2_fill_8 FILLER_0_100_1212 ();
 sg13g2_fill_8 FILLER_0_100_1220 ();
 sg13g2_fill_1 FILLER_0_101_0 ();
 sg13g2_fill_1 FILLER_0_101_27 ();
 sg13g2_fill_1 FILLER_0_101_33 ();
 sg13g2_fill_1 FILLER_0_101_44 ();
 sg13g2_fill_4 FILLER_0_101_81 ();
 sg13g2_fill_4 FILLER_0_101_93 ();
 sg13g2_fill_4 FILLER_0_101_101 ();
 sg13g2_fill_8 FILLER_0_101_136 ();
 sg13g2_fill_2 FILLER_0_101_144 ();
 sg13g2_fill_2 FILLER_0_101_191 ();
 sg13g2_fill_1 FILLER_0_101_193 ();
 sg13g2_fill_8 FILLER_0_101_199 ();
 sg13g2_fill_4 FILLER_0_101_207 ();
 sg13g2_fill_1 FILLER_0_101_211 ();
 sg13g2_fill_4 FILLER_0_101_247 ();
 sg13g2_fill_1 FILLER_0_101_251 ();
 sg13g2_fill_1 FILLER_0_101_260 ();
 sg13g2_decap_8 FILLER_0_101_291 ();
 sg13g2_fill_4 FILLER_0_101_302 ();
 sg13g2_fill_2 FILLER_0_101_319 ();
 sg13g2_fill_8 FILLER_0_101_352 ();
 sg13g2_fill_8 FILLER_0_101_360 ();
 sg13g2_fill_1 FILLER_0_101_399 ();
 sg13g2_fill_1 FILLER_0_101_404 ();
 sg13g2_fill_4 FILLER_0_101_415 ();
 sg13g2_fill_2 FILLER_0_101_424 ();
 sg13g2_fill_8 FILLER_0_101_491 ();
 sg13g2_fill_2 FILLER_0_101_499 ();
 sg13g2_fill_1 FILLER_0_101_531 ();
 sg13g2_fill_1 FILLER_0_101_536 ();
 sg13g2_fill_2 FILLER_0_101_563 ();
 sg13g2_fill_2 FILLER_0_101_575 ();
 sg13g2_fill_1 FILLER_0_101_577 ();
 sg13g2_fill_2 FILLER_0_101_604 ();
 sg13g2_fill_4 FILLER_0_101_610 ();
 sg13g2_fill_4 FILLER_0_101_633 ();
 sg13g2_fill_1 FILLER_0_101_647 ();
 sg13g2_fill_1 FILLER_0_101_658 ();
 sg13g2_fill_2 FILLER_0_101_664 ();
 sg13g2_fill_2 FILLER_0_101_692 ();
 sg13g2_fill_1 FILLER_0_101_694 ();
 sg13g2_fill_1 FILLER_0_101_699 ();
 sg13g2_fill_1 FILLER_0_101_728 ();
 sg13g2_fill_8 FILLER_0_101_733 ();
 sg13g2_fill_2 FILLER_0_101_840 ();
 sg13g2_fill_1 FILLER_0_101_896 ();
 sg13g2_fill_2 FILLER_0_101_920 ();
 sg13g2_decap_8 FILLER_0_101_926 ();
 sg13g2_fill_1 FILLER_0_101_942 ();
 sg13g2_fill_8 FILLER_0_101_961 ();
 sg13g2_fill_1 FILLER_0_101_986 ();
 sg13g2_fill_1 FILLER_0_101_998 ();
 sg13g2_fill_2 FILLER_0_101_1009 ();
 sg13g2_fill_1 FILLER_0_101_1011 ();
 sg13g2_fill_2 FILLER_0_101_1017 ();
 sg13g2_fill_1 FILLER_0_101_1026 ();
 sg13g2_fill_4 FILLER_0_101_1031 ();
 sg13g2_decap_8 FILLER_0_101_1038 ();
 sg13g2_fill_1 FILLER_0_101_1059 ();
 sg13g2_fill_1 FILLER_0_101_1065 ();
 sg13g2_fill_4 FILLER_0_101_1076 ();
 sg13g2_fill_1 FILLER_0_101_1093 ();
 sg13g2_fill_1 FILLER_0_101_1107 ();
 sg13g2_fill_1 FILLER_0_101_1116 ();
 sg13g2_decap_8 FILLER_0_101_1136 ();
 sg13g2_fill_2 FILLER_0_101_1147 ();
 sg13g2_fill_4 FILLER_0_101_1177 ();
 sg13g2_fill_1 FILLER_0_101_1181 ();
 sg13g2_fill_8 FILLER_0_101_1187 ();
 sg13g2_fill_8 FILLER_0_101_1195 ();
 sg13g2_fill_8 FILLER_0_101_1203 ();
 sg13g2_fill_8 FILLER_0_101_1211 ();
 sg13g2_fill_8 FILLER_0_101_1219 ();
 sg13g2_fill_1 FILLER_0_101_1227 ();
 sg13g2_fill_8 FILLER_0_102_0 ();
 sg13g2_fill_1 FILLER_0_102_8 ();
 sg13g2_fill_4 FILLER_0_102_64 ();
 sg13g2_fill_2 FILLER_0_102_80 ();
 sg13g2_fill_1 FILLER_0_102_82 ();
 sg13g2_fill_8 FILLER_0_102_105 ();
 sg13g2_fill_4 FILLER_0_102_117 ();
 sg13g2_fill_8 FILLER_0_102_131 ();
 sg13g2_fill_8 FILLER_0_102_139 ();
 sg13g2_fill_8 FILLER_0_102_147 ();
 sg13g2_fill_2 FILLER_0_102_155 ();
 sg13g2_fill_4 FILLER_0_102_162 ();
 sg13g2_fill_1 FILLER_0_102_166 ();
 sg13g2_fill_8 FILLER_0_102_171 ();
 sg13g2_decap_8 FILLER_0_102_179 ();
 sg13g2_fill_1 FILLER_0_102_190 ();
 sg13g2_fill_4 FILLER_0_102_251 ();
 sg13g2_fill_2 FILLER_0_102_255 ();
 sg13g2_fill_8 FILLER_0_102_282 ();
 sg13g2_fill_1 FILLER_0_102_290 ();
 sg13g2_fill_8 FILLER_0_102_353 ();
 sg13g2_fill_8 FILLER_0_102_361 ();
 sg13g2_fill_4 FILLER_0_102_369 ();
 sg13g2_fill_1 FILLER_0_102_373 ();
 sg13g2_fill_8 FILLER_0_102_386 ();
 sg13g2_fill_8 FILLER_0_102_394 ();
 sg13g2_fill_2 FILLER_0_102_402 ();
 sg13g2_decap_8 FILLER_0_102_408 ();
 sg13g2_fill_8 FILLER_0_102_447 ();
 sg13g2_fill_4 FILLER_0_102_455 ();
 sg13g2_fill_2 FILLER_0_102_459 ();
 sg13g2_fill_8 FILLER_0_102_478 ();
 sg13g2_fill_4 FILLER_0_102_486 ();
 sg13g2_fill_2 FILLER_0_102_490 ();
 sg13g2_fill_1 FILLER_0_102_522 ();
 sg13g2_fill_1 FILLER_0_102_533 ();
 sg13g2_fill_1 FILLER_0_102_549 ();
 sg13g2_fill_2 FILLER_0_102_560 ();
 sg13g2_fill_8 FILLER_0_102_588 ();
 sg13g2_fill_4 FILLER_0_102_596 ();
 sg13g2_fill_8 FILLER_0_102_608 ();
 sg13g2_fill_2 FILLER_0_102_616 ();
 sg13g2_fill_1 FILLER_0_102_618 ();
 sg13g2_fill_4 FILLER_0_102_683 ();
 sg13g2_fill_8 FILLER_0_102_713 ();
 sg13g2_fill_2 FILLER_0_102_721 ();
 sg13g2_fill_1 FILLER_0_102_723 ();
 sg13g2_fill_4 FILLER_0_102_729 ();
 sg13g2_fill_1 FILLER_0_102_733 ();
 sg13g2_fill_8 FILLER_0_102_744 ();
 sg13g2_fill_1 FILLER_0_102_791 ();
 sg13g2_fill_1 FILLER_0_102_802 ();
 sg13g2_fill_1 FILLER_0_102_808 ();
 sg13g2_fill_2 FILLER_0_102_813 ();
 sg13g2_decap_8 FILLER_0_102_841 ();
 sg13g2_fill_8 FILLER_0_102_852 ();
 sg13g2_fill_8 FILLER_0_102_860 ();
 sg13g2_fill_1 FILLER_0_102_872 ();
 sg13g2_fill_4 FILLER_0_102_882 ();
 sg13g2_fill_2 FILLER_0_102_886 ();
 sg13g2_fill_1 FILLER_0_102_895 ();
 sg13g2_fill_2 FILLER_0_102_905 ();
 sg13g2_fill_1 FILLER_0_102_911 ();
 sg13g2_fill_1 FILLER_0_102_917 ();
 sg13g2_fill_1 FILLER_0_102_936 ();
 sg13g2_fill_1 FILLER_0_102_942 ();
 sg13g2_fill_1 FILLER_0_102_956 ();
 sg13g2_fill_2 FILLER_0_102_962 ();
 sg13g2_fill_1 FILLER_0_102_964 ();
 sg13g2_fill_4 FILLER_0_102_971 ();
 sg13g2_fill_2 FILLER_0_102_975 ();
 sg13g2_fill_4 FILLER_0_102_983 ();
 sg13g2_fill_1 FILLER_0_102_987 ();
 sg13g2_fill_4 FILLER_0_102_993 ();
 sg13g2_fill_1 FILLER_0_102_997 ();
 sg13g2_fill_2 FILLER_0_102_1038 ();
 sg13g2_fill_1 FILLER_0_102_1040 ();
 sg13g2_fill_2 FILLER_0_102_1074 ();
 sg13g2_fill_4 FILLER_0_102_1081 ();
 sg13g2_fill_1 FILLER_0_102_1085 ();
 sg13g2_fill_4 FILLER_0_102_1095 ();
 sg13g2_fill_1 FILLER_0_102_1103 ();
 sg13g2_fill_1 FILLER_0_102_1179 ();
 sg13g2_fill_8 FILLER_0_102_1196 ();
 sg13g2_fill_8 FILLER_0_102_1204 ();
 sg13g2_fill_8 FILLER_0_102_1212 ();
 sg13g2_fill_8 FILLER_0_102_1220 ();
 sg13g2_fill_4 FILLER_0_103_0 ();
 sg13g2_fill_1 FILLER_0_103_4 ();
 sg13g2_fill_4 FILLER_0_103_36 ();
 sg13g2_fill_8 FILLER_0_103_44 ();
 sg13g2_fill_8 FILLER_0_103_56 ();
 sg13g2_fill_8 FILLER_0_103_64 ();
 sg13g2_fill_1 FILLER_0_103_138 ();
 sg13g2_fill_2 FILLER_0_103_175 ();
 sg13g2_fill_1 FILLER_0_103_177 ();
 sg13g2_fill_2 FILLER_0_103_183 ();
 sg13g2_fill_2 FILLER_0_103_216 ();
 sg13g2_fill_2 FILLER_0_103_228 ();
 sg13g2_fill_1 FILLER_0_103_230 ();
 sg13g2_fill_1 FILLER_0_103_241 ();
 sg13g2_fill_2 FILLER_0_103_252 ();
 sg13g2_fill_1 FILLER_0_103_254 ();
 sg13g2_fill_8 FILLER_0_103_286 ();
 sg13g2_fill_1 FILLER_0_103_339 ();
 sg13g2_fill_2 FILLER_0_103_350 ();
 sg13g2_fill_8 FILLER_0_103_383 ();
 sg13g2_fill_2 FILLER_0_103_391 ();
 sg13g2_fill_1 FILLER_0_103_393 ();
 sg13g2_decap_8 FILLER_0_103_398 ();
 sg13g2_fill_1 FILLER_0_103_410 ();
 sg13g2_fill_1 FILLER_0_103_429 ();
 sg13g2_fill_2 FILLER_0_103_456 ();
 sg13g2_fill_1 FILLER_0_103_458 ();
 sg13g2_fill_2 FILLER_0_103_463 ();
 sg13g2_fill_1 FILLER_0_103_465 ();
 sg13g2_fill_4 FILLER_0_103_476 ();
 sg13g2_fill_1 FILLER_0_103_480 ();
 sg13g2_fill_4 FILLER_0_103_485 ();
 sg13g2_fill_1 FILLER_0_103_489 ();
 sg13g2_fill_2 FILLER_0_103_494 ();
 sg13g2_fill_1 FILLER_0_103_496 ();
 sg13g2_fill_2 FILLER_0_103_501 ();
 sg13g2_fill_8 FILLER_0_103_522 ();
 sg13g2_fill_8 FILLER_0_103_530 ();
 sg13g2_fill_2 FILLER_0_103_538 ();
 sg13g2_fill_1 FILLER_0_103_540 ();
 sg13g2_fill_8 FILLER_0_103_580 ();
 sg13g2_fill_8 FILLER_0_103_588 ();
 sg13g2_fill_8 FILLER_0_103_596 ();
 sg13g2_fill_4 FILLER_0_103_604 ();
 sg13g2_fill_8 FILLER_0_103_612 ();
 sg13g2_fill_4 FILLER_0_103_620 ();
 sg13g2_fill_1 FILLER_0_103_624 ();
 sg13g2_fill_8 FILLER_0_103_629 ();
 sg13g2_fill_8 FILLER_0_103_637 ();
 sg13g2_fill_1 FILLER_0_103_650 ();
 sg13g2_fill_1 FILLER_0_103_656 ();
 sg13g2_fill_8 FILLER_0_103_671 ();
 sg13g2_fill_4 FILLER_0_103_679 ();
 sg13g2_fill_1 FILLER_0_103_683 ();
 sg13g2_fill_4 FILLER_0_103_714 ();
 sg13g2_fill_2 FILLER_0_103_718 ();
 sg13g2_decap_8 FILLER_0_103_750 ();
 sg13g2_fill_4 FILLER_0_103_767 ();
 sg13g2_fill_2 FILLER_0_103_775 ();
 sg13g2_fill_8 FILLER_0_103_787 ();
 sg13g2_fill_4 FILLER_0_103_795 ();
 sg13g2_fill_1 FILLER_0_103_799 ();
 sg13g2_fill_8 FILLER_0_103_882 ();
 sg13g2_fill_1 FILLER_0_103_894 ();
 sg13g2_fill_2 FILLER_0_103_907 ();
 sg13g2_fill_1 FILLER_0_103_929 ();
 sg13g2_fill_1 FILLER_0_103_935 ();
 sg13g2_fill_1 FILLER_0_103_941 ();
 sg13g2_fill_1 FILLER_0_103_951 ();
 sg13g2_fill_2 FILLER_0_103_956 ();
 sg13g2_fill_1 FILLER_0_103_958 ();
 sg13g2_fill_1 FILLER_0_103_964 ();
 sg13g2_fill_1 FILLER_0_103_969 ();
 sg13g2_fill_2 FILLER_0_103_975 ();
 sg13g2_fill_1 FILLER_0_103_985 ();
 sg13g2_fill_4 FILLER_0_103_991 ();
 sg13g2_fill_1 FILLER_0_103_995 ();
 sg13g2_fill_1 FILLER_0_103_1008 ();
 sg13g2_fill_2 FILLER_0_103_1014 ();
 sg13g2_fill_1 FILLER_0_103_1024 ();
 sg13g2_fill_4 FILLER_0_103_1029 ();
 sg13g2_fill_1 FILLER_0_103_1033 ();
 sg13g2_fill_2 FILLER_0_103_1057 ();
 sg13g2_fill_2 FILLER_0_103_1063 ();
 sg13g2_fill_2 FILLER_0_103_1088 ();
 sg13g2_fill_1 FILLER_0_103_1099 ();
 sg13g2_fill_1 FILLER_0_103_1109 ();
 sg13g2_fill_1 FILLER_0_103_1123 ();
 sg13g2_fill_1 FILLER_0_103_1129 ();
 sg13g2_fill_1 FILLER_0_103_1171 ();
 sg13g2_fill_2 FILLER_0_103_1188 ();
 sg13g2_fill_1 FILLER_0_103_1190 ();
 sg13g2_fill_8 FILLER_0_103_1195 ();
 sg13g2_fill_8 FILLER_0_103_1203 ();
 sg13g2_fill_8 FILLER_0_103_1211 ();
 sg13g2_fill_8 FILLER_0_103_1219 ();
 sg13g2_fill_1 FILLER_0_103_1227 ();
 sg13g2_fill_8 FILLER_0_104_0 ();
 sg13g2_fill_2 FILLER_0_104_8 ();
 sg13g2_fill_1 FILLER_0_104_10 ();
 sg13g2_fill_2 FILLER_0_104_29 ();
 sg13g2_fill_2 FILLER_0_104_36 ();
 sg13g2_fill_1 FILLER_0_104_77 ();
 sg13g2_fill_2 FILLER_0_104_152 ();
 sg13g2_fill_8 FILLER_0_104_158 ();
 sg13g2_fill_4 FILLER_0_104_166 ();
 sg13g2_fill_2 FILLER_0_104_170 ();
 sg13g2_fill_2 FILLER_0_104_176 ();
 sg13g2_fill_2 FILLER_0_104_204 ();
 sg13g2_fill_4 FILLER_0_104_210 ();
 sg13g2_fill_8 FILLER_0_104_224 ();
 sg13g2_fill_2 FILLER_0_104_232 ();
 sg13g2_fill_1 FILLER_0_104_234 ();
 sg13g2_fill_2 FILLER_0_104_239 ();
 sg13g2_fill_1 FILLER_0_104_241 ();
 sg13g2_fill_4 FILLER_0_104_252 ();
 sg13g2_fill_1 FILLER_0_104_256 ();
 sg13g2_fill_4 FILLER_0_104_261 ();
 sg13g2_fill_1 FILLER_0_104_265 ();
 sg13g2_fill_2 FILLER_0_104_270 ();
 sg13g2_fill_1 FILLER_0_104_272 ();
 sg13g2_decap_8 FILLER_0_104_283 ();
 sg13g2_fill_4 FILLER_0_104_299 ();
 sg13g2_fill_2 FILLER_0_104_313 ();
 sg13g2_fill_1 FILLER_0_104_325 ();
 sg13g2_fill_2 FILLER_0_104_330 ();
 sg13g2_fill_1 FILLER_0_104_336 ();
 sg13g2_fill_2 FILLER_0_104_341 ();
 sg13g2_fill_1 FILLER_0_104_353 ();
 sg13g2_fill_1 FILLER_0_104_359 ();
 sg13g2_fill_4 FILLER_0_104_386 ();
 sg13g2_fill_1 FILLER_0_104_390 ();
 sg13g2_fill_8 FILLER_0_104_427 ();
 sg13g2_fill_1 FILLER_0_104_435 ();
 sg13g2_fill_1 FILLER_0_104_441 ();
 sg13g2_fill_1 FILLER_0_104_446 ();
 sg13g2_fill_1 FILLER_0_104_473 ();
 sg13g2_fill_1 FILLER_0_104_505 ();
 sg13g2_fill_8 FILLER_0_104_524 ();
 sg13g2_fill_8 FILLER_0_104_536 ();
 sg13g2_fill_8 FILLER_0_104_544 ();
 sg13g2_fill_8 FILLER_0_104_552 ();
 sg13g2_decap_8 FILLER_0_104_560 ();
 sg13g2_fill_4 FILLER_0_104_597 ();
 sg13g2_fill_4 FILLER_0_104_632 ();
 sg13g2_fill_2 FILLER_0_104_636 ();
 sg13g2_fill_2 FILLER_0_104_648 ();
 sg13g2_fill_8 FILLER_0_104_669 ();
 sg13g2_fill_8 FILLER_0_104_677 ();
 sg13g2_fill_2 FILLER_0_104_685 ();
 sg13g2_fill_1 FILLER_0_104_687 ();
 sg13g2_fill_4 FILLER_0_104_745 ();
 sg13g2_fill_2 FILLER_0_104_749 ();
 sg13g2_fill_4 FILLER_0_104_786 ();
 sg13g2_fill_2 FILLER_0_104_800 ();
 sg13g2_decap_8 FILLER_0_104_812 ();
 sg13g2_fill_8 FILLER_0_104_827 ();
 sg13g2_fill_8 FILLER_0_104_835 ();
 sg13g2_fill_8 FILLER_0_104_843 ();
 sg13g2_fill_2 FILLER_0_104_891 ();
 sg13g2_fill_1 FILLER_0_104_893 ();
 sg13g2_fill_1 FILLER_0_104_908 ();
 sg13g2_fill_2 FILLER_0_104_929 ();
 sg13g2_fill_2 FILLER_0_104_940 ();
 sg13g2_fill_1 FILLER_0_104_942 ();
 sg13g2_fill_2 FILLER_0_104_952 ();
 sg13g2_fill_1 FILLER_0_104_954 ();
 sg13g2_fill_1 FILLER_0_104_969 ();
 sg13g2_fill_2 FILLER_0_104_996 ();
 sg13g2_fill_1 FILLER_0_104_1025 ();
 sg13g2_fill_1 FILLER_0_104_1047 ();
 sg13g2_fill_1 FILLER_0_104_1052 ();
 sg13g2_fill_2 FILLER_0_104_1058 ();
 sg13g2_fill_1 FILLER_0_104_1064 ();
 sg13g2_fill_2 FILLER_0_104_1071 ();
 sg13g2_fill_1 FILLER_0_104_1073 ();
 sg13g2_fill_4 FILLER_0_104_1096 ();
 sg13g2_decap_8 FILLER_0_104_1114 ();
 sg13g2_fill_2 FILLER_0_104_1146 ();
 sg13g2_fill_8 FILLER_0_104_1186 ();
 sg13g2_fill_8 FILLER_0_104_1194 ();
 sg13g2_fill_8 FILLER_0_104_1202 ();
 sg13g2_fill_8 FILLER_0_104_1210 ();
 sg13g2_fill_8 FILLER_0_104_1218 ();
 sg13g2_fill_2 FILLER_0_104_1226 ();
 sg13g2_decap_8 FILLER_0_105_0 ();
 sg13g2_fill_8 FILLER_0_105_33 ();
 sg13g2_fill_1 FILLER_0_105_41 ();
 sg13g2_fill_2 FILLER_0_105_88 ();
 sg13g2_fill_8 FILLER_0_105_110 ();
 sg13g2_fill_1 FILLER_0_105_133 ();
 sg13g2_fill_8 FILLER_0_105_209 ();
 sg13g2_fill_4 FILLER_0_105_217 ();
 sg13g2_fill_2 FILLER_0_105_221 ();
 sg13g2_fill_2 FILLER_0_105_280 ();
 sg13g2_fill_2 FILLER_0_105_313 ();
 sg13g2_fill_2 FILLER_0_105_372 ();
 sg13g2_fill_8 FILLER_0_105_378 ();
 sg13g2_fill_4 FILLER_0_105_386 ();
 sg13g2_fill_8 FILLER_0_105_426 ();
 sg13g2_fill_2 FILLER_0_105_434 ();
 sg13g2_fill_1 FILLER_0_105_460 ();
 sg13g2_fill_2 FILLER_0_105_471 ();
 sg13g2_fill_1 FILLER_0_105_478 ();
 sg13g2_fill_2 FILLER_0_105_483 ();
 sg13g2_fill_4 FILLER_0_105_516 ();
 sg13g2_fill_8 FILLER_0_105_551 ();
 sg13g2_decap_8 FILLER_0_105_559 ();
 sg13g2_fill_2 FILLER_0_105_617 ();
 sg13g2_fill_2 FILLER_0_105_645 ();
 sg13g2_fill_8 FILLER_0_105_673 ();
 sg13g2_fill_8 FILLER_0_105_681 ();
 sg13g2_fill_4 FILLER_0_105_689 ();
 sg13g2_fill_1 FILLER_0_105_693 ();
 sg13g2_fill_1 FILLER_0_105_699 ();
 sg13g2_fill_1 FILLER_0_105_710 ();
 sg13g2_fill_1 FILLER_0_105_726 ();
 sg13g2_fill_1 FILLER_0_105_731 ();
 sg13g2_fill_8 FILLER_0_105_742 ();
 sg13g2_fill_1 FILLER_0_105_750 ();
 sg13g2_fill_1 FILLER_0_105_776 ();
 sg13g2_fill_8 FILLER_0_105_827 ();
 sg13g2_fill_8 FILLER_0_105_835 ();
 sg13g2_fill_8 FILLER_0_105_843 ();
 sg13g2_fill_2 FILLER_0_105_851 ();
 sg13g2_decap_8 FILLER_0_105_858 ();
 sg13g2_fill_4 FILLER_0_105_891 ();
 sg13g2_fill_1 FILLER_0_105_905 ();
 sg13g2_fill_2 FILLER_0_105_919 ();
 sg13g2_decap_8 FILLER_0_105_925 ();
 sg13g2_fill_4 FILLER_0_105_937 ();
 sg13g2_fill_4 FILLER_0_105_963 ();
 sg13g2_fill_2 FILLER_0_105_967 ();
 sg13g2_fill_4 FILLER_0_105_973 ();
 sg13g2_fill_4 FILLER_0_105_982 ();
 sg13g2_fill_1 FILLER_0_105_991 ();
 sg13g2_fill_2 FILLER_0_105_997 ();
 sg13g2_fill_1 FILLER_0_105_999 ();
 sg13g2_decap_8 FILLER_0_105_1026 ();
 sg13g2_fill_1 FILLER_0_105_1047 ();
 sg13g2_fill_4 FILLER_0_105_1066 ();
 sg13g2_fill_8 FILLER_0_105_1075 ();
 sg13g2_fill_2 FILLER_0_105_1083 ();
 sg13g2_fill_1 FILLER_0_105_1085 ();
 sg13g2_fill_8 FILLER_0_105_1113 ();
 sg13g2_fill_8 FILLER_0_105_1121 ();
 sg13g2_fill_2 FILLER_0_105_1129 ();
 sg13g2_fill_1 FILLER_0_105_1131 ();
 sg13g2_fill_8 FILLER_0_105_1136 ();
 sg13g2_fill_4 FILLER_0_105_1144 ();
 sg13g2_fill_1 FILLER_0_105_1148 ();
 sg13g2_fill_2 FILLER_0_105_1153 ();
 sg13g2_fill_1 FILLER_0_105_1165 ();
 sg13g2_fill_2 FILLER_0_105_1171 ();
 sg13g2_fill_4 FILLER_0_105_1178 ();
 sg13g2_fill_1 FILLER_0_105_1182 ();
 sg13g2_fill_1 FILLER_0_105_1188 ();
 sg13g2_fill_8 FILLER_0_105_1194 ();
 sg13g2_fill_8 FILLER_0_105_1202 ();
 sg13g2_fill_8 FILLER_0_105_1210 ();
 sg13g2_fill_8 FILLER_0_105_1218 ();
 sg13g2_fill_2 FILLER_0_105_1226 ();
 sg13g2_fill_2 FILLER_0_106_0 ();
 sg13g2_fill_2 FILLER_0_106_37 ();
 sg13g2_fill_1 FILLER_0_106_39 ();
 sg13g2_fill_2 FILLER_0_106_54 ();
 sg13g2_fill_2 FILLER_0_106_66 ();
 sg13g2_fill_1 FILLER_0_106_68 ();
 sg13g2_fill_2 FILLER_0_106_73 ();
 sg13g2_fill_8 FILLER_0_106_109 ();
 sg13g2_decap_8 FILLER_0_106_117 ();
 sg13g2_fill_2 FILLER_0_106_128 ();
 sg13g2_fill_1 FILLER_0_106_130 ();
 sg13g2_fill_1 FILLER_0_106_136 ();
 sg13g2_fill_4 FILLER_0_106_151 ();
 sg13g2_fill_2 FILLER_0_106_155 ();
 sg13g2_fill_1 FILLER_0_106_161 ();
 sg13g2_fill_1 FILLER_0_106_175 ();
 sg13g2_fill_8 FILLER_0_106_196 ();
 sg13g2_fill_2 FILLER_0_106_204 ();
 sg13g2_fill_1 FILLER_0_106_206 ();
 sg13g2_fill_2 FILLER_0_106_248 ();
 sg13g2_fill_1 FILLER_0_106_250 ();
 sg13g2_fill_2 FILLER_0_106_264 ();
 sg13g2_fill_1 FILLER_0_106_266 ();
 sg13g2_fill_8 FILLER_0_106_279 ();
 sg13g2_fill_4 FILLER_0_106_287 ();
 sg13g2_fill_4 FILLER_0_106_295 ();
 sg13g2_fill_2 FILLER_0_106_325 ();
 sg13g2_fill_2 FILLER_0_106_331 ();
 sg13g2_fill_8 FILLER_0_106_368 ();
 sg13g2_decap_8 FILLER_0_106_376 ();
 sg13g2_decap_8 FILLER_0_106_388 ();
 sg13g2_fill_2 FILLER_0_106_399 ();
 sg13g2_fill_1 FILLER_0_106_401 ();
 sg13g2_decap_8 FILLER_0_106_433 ();
 sg13g2_fill_1 FILLER_0_106_455 ();
 sg13g2_fill_4 FILLER_0_106_461 ();
 sg13g2_fill_1 FILLER_0_106_465 ();
 sg13g2_fill_2 FILLER_0_106_471 ();
 sg13g2_fill_1 FILLER_0_106_473 ();
 sg13g2_fill_8 FILLER_0_106_478 ();
 sg13g2_fill_2 FILLER_0_106_486 ();
 sg13g2_fill_8 FILLER_0_106_558 ();
 sg13g2_fill_4 FILLER_0_106_566 ();
 sg13g2_fill_2 FILLER_0_106_604 ();
 sg13g2_fill_1 FILLER_0_106_606 ();
 sg13g2_fill_4 FILLER_0_106_612 ();
 sg13g2_fill_2 FILLER_0_106_646 ();
 sg13g2_fill_8 FILLER_0_106_684 ();
 sg13g2_fill_8 FILLER_0_106_692 ();
 sg13g2_fill_8 FILLER_0_106_704 ();
 sg13g2_fill_8 FILLER_0_106_712 ();
 sg13g2_fill_8 FILLER_0_106_720 ();
 sg13g2_fill_4 FILLER_0_106_728 ();
 sg13g2_fill_8 FILLER_0_106_818 ();
 sg13g2_fill_8 FILLER_0_106_826 ();
 sg13g2_fill_8 FILLER_0_106_895 ();
 sg13g2_fill_2 FILLER_0_106_903 ();
 sg13g2_decap_8 FILLER_0_106_917 ();
 sg13g2_fill_1 FILLER_0_106_936 ();
 sg13g2_fill_1 FILLER_0_106_953 ();
 sg13g2_fill_1 FILLER_0_106_958 ();
 sg13g2_fill_2 FILLER_0_106_964 ();
 sg13g2_fill_4 FILLER_0_106_970 ();
 sg13g2_fill_8 FILLER_0_106_983 ();
 sg13g2_fill_8 FILLER_0_106_991 ();
 sg13g2_fill_8 FILLER_0_106_999 ();
 sg13g2_fill_2 FILLER_0_106_1007 ();
 sg13g2_fill_8 FILLER_0_106_1031 ();
 sg13g2_fill_1 FILLER_0_106_1039 ();
 sg13g2_decap_8 FILLER_0_106_1045 ();
 sg13g2_decap_8 FILLER_0_106_1066 ();
 sg13g2_fill_8 FILLER_0_106_1077 ();
 sg13g2_fill_4 FILLER_0_106_1085 ();
 sg13g2_fill_2 FILLER_0_106_1089 ();
 sg13g2_fill_2 FILLER_0_106_1101 ();
 sg13g2_fill_1 FILLER_0_106_1103 ();
 sg13g2_fill_4 FILLER_0_106_1124 ();
 sg13g2_fill_1 FILLER_0_106_1128 ();
 sg13g2_fill_4 FILLER_0_106_1144 ();
 sg13g2_fill_2 FILLER_0_106_1148 ();
 sg13g2_fill_8 FILLER_0_106_1155 ();
 sg13g2_fill_4 FILLER_0_106_1163 ();
 sg13g2_fill_2 FILLER_0_106_1177 ();
 sg13g2_fill_8 FILLER_0_106_1197 ();
 sg13g2_fill_8 FILLER_0_106_1205 ();
 sg13g2_fill_8 FILLER_0_106_1213 ();
 sg13g2_decap_8 FILLER_0_106_1221 ();
 sg13g2_fill_8 FILLER_0_107_0 ();
 sg13g2_fill_8 FILLER_0_107_8 ();
 sg13g2_fill_2 FILLER_0_107_16 ();
 sg13g2_fill_1 FILLER_0_107_18 ();
 sg13g2_fill_8 FILLER_0_107_29 ();
 sg13g2_fill_8 FILLER_0_107_37 ();
 sg13g2_fill_4 FILLER_0_107_45 ();
 sg13g2_fill_2 FILLER_0_107_49 ();
 sg13g2_fill_8 FILLER_0_107_74 ();
 sg13g2_fill_8 FILLER_0_107_86 ();
 sg13g2_fill_2 FILLER_0_107_94 ();
 sg13g2_fill_8 FILLER_0_107_118 ();
 sg13g2_fill_4 FILLER_0_107_126 ();
 sg13g2_fill_1 FILLER_0_107_130 ();
 sg13g2_fill_8 FILLER_0_107_139 ();
 sg13g2_fill_8 FILLER_0_107_147 ();
 sg13g2_fill_4 FILLER_0_107_155 ();
 sg13g2_fill_4 FILLER_0_107_195 ();
 sg13g2_fill_8 FILLER_0_107_227 ();
 sg13g2_fill_8 FILLER_0_107_235 ();
 sg13g2_fill_8 FILLER_0_107_243 ();
 sg13g2_fill_1 FILLER_0_107_251 ();
 sg13g2_fill_4 FILLER_0_107_256 ();
 sg13g2_fill_1 FILLER_0_107_260 ();
 sg13g2_fill_8 FILLER_0_107_269 ();
 sg13g2_fill_4 FILLER_0_107_277 ();
 sg13g2_fill_2 FILLER_0_107_281 ();
 sg13g2_fill_8 FILLER_0_107_287 ();
 sg13g2_fill_8 FILLER_0_107_295 ();
 sg13g2_fill_2 FILLER_0_107_303 ();
 sg13g2_fill_1 FILLER_0_107_305 ();
 sg13g2_fill_4 FILLER_0_107_310 ();
 sg13g2_fill_1 FILLER_0_107_314 ();
 sg13g2_fill_2 FILLER_0_107_354 ();
 sg13g2_fill_1 FILLER_0_107_356 ();
 sg13g2_fill_2 FILLER_0_107_383 ();
 sg13g2_fill_8 FILLER_0_107_393 ();
 sg13g2_fill_4 FILLER_0_107_401 ();
 sg13g2_fill_1 FILLER_0_107_405 ();
 sg13g2_fill_8 FILLER_0_107_451 ();
 sg13g2_fill_2 FILLER_0_107_464 ();
 sg13g2_fill_8 FILLER_0_107_492 ();
 sg13g2_fill_4 FILLER_0_107_500 ();
 sg13g2_fill_4 FILLER_0_107_519 ();
 sg13g2_fill_4 FILLER_0_107_555 ();
 sg13g2_fill_8 FILLER_0_107_607 ();
 sg13g2_fill_2 FILLER_0_107_615 ();
 sg13g2_fill_1 FILLER_0_107_617 ();
 sg13g2_fill_4 FILLER_0_107_623 ();
 sg13g2_fill_1 FILLER_0_107_627 ();
 sg13g2_fill_1 FILLER_0_107_632 ();
 sg13g2_fill_1 FILLER_0_107_647 ();
 sg13g2_fill_1 FILLER_0_107_665 ();
 sg13g2_fill_8 FILLER_0_107_692 ();
 sg13g2_decap_8 FILLER_0_107_700 ();
 sg13g2_fill_8 FILLER_0_107_717 ();
 sg13g2_fill_8 FILLER_0_107_725 ();
 sg13g2_fill_8 FILLER_0_107_733 ();
 sg13g2_fill_8 FILLER_0_107_745 ();
 sg13g2_fill_8 FILLER_0_107_753 ();
 sg13g2_fill_4 FILLER_0_107_761 ();
 sg13g2_fill_2 FILLER_0_107_765 ();
 sg13g2_fill_4 FILLER_0_107_771 ();
 sg13g2_fill_1 FILLER_0_107_775 ();
 sg13g2_fill_8 FILLER_0_107_812 ();
 sg13g2_fill_8 FILLER_0_107_820 ();
 sg13g2_fill_8 FILLER_0_107_828 ();
 sg13g2_fill_4 FILLER_0_107_836 ();
 sg13g2_fill_4 FILLER_0_107_844 ();
 sg13g2_fill_1 FILLER_0_107_848 ();
 sg13g2_fill_1 FILLER_0_107_853 ();
 sg13g2_fill_8 FILLER_0_107_880 ();
 sg13g2_decap_8 FILLER_0_107_888 ();
 sg13g2_fill_1 FILLER_0_107_909 ();
 sg13g2_fill_8 FILLER_0_107_914 ();
 sg13g2_fill_1 FILLER_0_107_922 ();
 sg13g2_fill_1 FILLER_0_107_927 ();
 sg13g2_fill_2 FILLER_0_107_948 ();
 sg13g2_fill_1 FILLER_0_107_963 ();
 sg13g2_fill_2 FILLER_0_107_975 ();
 sg13g2_fill_1 FILLER_0_107_977 ();
 sg13g2_fill_1 FILLER_0_107_982 ();
 sg13g2_fill_2 FILLER_0_107_990 ();
 sg13g2_fill_1 FILLER_0_107_992 ();
 sg13g2_decap_8 FILLER_0_107_998 ();
 sg13g2_fill_1 FILLER_0_107_1021 ();
 sg13g2_fill_2 FILLER_0_107_1027 ();
 sg13g2_fill_2 FILLER_0_107_1034 ();
 sg13g2_fill_1 FILLER_0_107_1070 ();
 sg13g2_fill_1 FILLER_0_107_1095 ();
 sg13g2_fill_1 FILLER_0_107_1103 ();
 sg13g2_fill_4 FILLER_0_107_1115 ();
 sg13g2_fill_8 FILLER_0_107_1124 ();
 sg13g2_fill_4 FILLER_0_107_1132 ();
 sg13g2_fill_1 FILLER_0_107_1173 ();
 sg13g2_fill_8 FILLER_0_107_1190 ();
 sg13g2_fill_8 FILLER_0_107_1198 ();
 sg13g2_fill_8 FILLER_0_107_1206 ();
 sg13g2_fill_8 FILLER_0_107_1214 ();
 sg13g2_fill_4 FILLER_0_107_1222 ();
 sg13g2_fill_2 FILLER_0_107_1226 ();
 sg13g2_fill_2 FILLER_0_108_0 ();
 sg13g2_fill_1 FILLER_0_108_2 ();
 sg13g2_fill_1 FILLER_0_108_29 ();
 sg13g2_fill_4 FILLER_0_108_43 ();
 sg13g2_fill_1 FILLER_0_108_47 ();
 sg13g2_fill_8 FILLER_0_108_78 ();
 sg13g2_fill_1 FILLER_0_108_86 ();
 sg13g2_fill_1 FILLER_0_108_118 ();
 sg13g2_fill_8 FILLER_0_108_145 ();
 sg13g2_fill_4 FILLER_0_108_153 ();
 sg13g2_fill_2 FILLER_0_108_157 ();
 sg13g2_fill_4 FILLER_0_108_235 ();
 sg13g2_fill_1 FILLER_0_108_239 ();
 sg13g2_fill_1 FILLER_0_108_250 ();
 sg13g2_fill_4 FILLER_0_108_291 ();
 sg13g2_fill_1 FILLER_0_108_295 ();
 sg13g2_fill_8 FILLER_0_108_300 ();
 sg13g2_fill_8 FILLER_0_108_308 ();
 sg13g2_fill_8 FILLER_0_108_316 ();
 sg13g2_fill_2 FILLER_0_108_324 ();
 sg13g2_fill_2 FILLER_0_108_360 ();
 sg13g2_decap_8 FILLER_0_108_411 ();
 sg13g2_fill_1 FILLER_0_108_454 ();
 sg13g2_fill_8 FILLER_0_108_491 ();
 sg13g2_fill_8 FILLER_0_108_499 ();
 sg13g2_fill_1 FILLER_0_108_507 ();
 sg13g2_fill_8 FILLER_0_108_512 ();
 sg13g2_fill_2 FILLER_0_108_520 ();
 sg13g2_fill_1 FILLER_0_108_522 ();
 sg13g2_fill_8 FILLER_0_108_599 ();
 sg13g2_fill_8 FILLER_0_108_607 ();
 sg13g2_fill_4 FILLER_0_108_619 ();
 sg13g2_fill_2 FILLER_0_108_623 ();
 sg13g2_fill_2 FILLER_0_108_651 ();
 sg13g2_fill_8 FILLER_0_108_682 ();
 sg13g2_fill_2 FILLER_0_108_690 ();
 sg13g2_fill_1 FILLER_0_108_692 ();
 sg13g2_fill_1 FILLER_0_108_728 ();
 sg13g2_fill_8 FILLER_0_108_760 ();
 sg13g2_fill_8 FILLER_0_108_768 ();
 sg13g2_decap_8 FILLER_0_108_776 ();
 sg13g2_fill_8 FILLER_0_108_787 ();
 sg13g2_fill_8 FILLER_0_108_795 ();
 sg13g2_fill_8 FILLER_0_108_803 ();
 sg13g2_fill_8 FILLER_0_108_811 ();
 sg13g2_fill_8 FILLER_0_108_819 ();
 sg13g2_fill_8 FILLER_0_108_827 ();
 sg13g2_fill_4 FILLER_0_108_835 ();
 sg13g2_fill_2 FILLER_0_108_865 ();
 sg13g2_fill_8 FILLER_0_108_882 ();
 sg13g2_fill_8 FILLER_0_108_890 ();
 sg13g2_fill_4 FILLER_0_108_898 ();
 sg13g2_fill_2 FILLER_0_108_902 ();
 sg13g2_fill_2 FILLER_0_108_927 ();
 sg13g2_fill_1 FILLER_0_108_929 ();
 sg13g2_fill_2 FILLER_0_108_935 ();
 sg13g2_fill_1 FILLER_0_108_946 ();
 sg13g2_fill_1 FILLER_0_108_953 ();
 sg13g2_fill_2 FILLER_0_108_962 ();
 sg13g2_fill_4 FILLER_0_108_969 ();
 sg13g2_fill_4 FILLER_0_108_993 ();
 sg13g2_fill_2 FILLER_0_108_997 ();
 sg13g2_fill_8 FILLER_0_108_1010 ();
 sg13g2_fill_1 FILLER_0_108_1018 ();
 sg13g2_fill_2 FILLER_0_108_1027 ();
 sg13g2_fill_2 FILLER_0_108_1051 ();
 sg13g2_fill_1 FILLER_0_108_1053 ();
 sg13g2_fill_2 FILLER_0_108_1059 ();
 sg13g2_fill_1 FILLER_0_108_1070 ();
 sg13g2_fill_1 FILLER_0_108_1075 ();
 sg13g2_fill_1 FILLER_0_108_1086 ();
 sg13g2_fill_2 FILLER_0_108_1099 ();
 sg13g2_fill_2 FILLER_0_108_1126 ();
 sg13g2_fill_1 FILLER_0_108_1128 ();
 sg13g2_fill_2 FILLER_0_108_1134 ();
 sg13g2_fill_1 FILLER_0_108_1136 ();
 sg13g2_fill_1 FILLER_0_108_1142 ();
 sg13g2_fill_1 FILLER_0_108_1147 ();
 sg13g2_fill_1 FILLER_0_108_1153 ();
 sg13g2_fill_1 FILLER_0_108_1159 ();
 sg13g2_fill_2 FILLER_0_108_1165 ();
 sg13g2_fill_8 FILLER_0_108_1210 ();
 sg13g2_fill_8 FILLER_0_108_1218 ();
 sg13g2_fill_2 FILLER_0_108_1226 ();
 sg13g2_fill_4 FILLER_0_109_67 ();
 sg13g2_fill_1 FILLER_0_109_71 ();
 sg13g2_fill_2 FILLER_0_109_123 ();
 sg13g2_fill_8 FILLER_0_109_155 ();
 sg13g2_fill_2 FILLER_0_109_163 ();
 sg13g2_fill_1 FILLER_0_109_165 ();
 sg13g2_fill_1 FILLER_0_109_170 ();
 sg13g2_fill_1 FILLER_0_109_197 ();
 sg13g2_fill_1 FILLER_0_109_203 ();
 sg13g2_fill_2 FILLER_0_109_214 ();
 sg13g2_fill_1 FILLER_0_109_242 ();
 sg13g2_fill_1 FILLER_0_109_269 ();
 sg13g2_fill_8 FILLER_0_109_305 ();
 sg13g2_fill_8 FILLER_0_109_313 ();
 sg13g2_fill_8 FILLER_0_109_321 ();
 sg13g2_fill_1 FILLER_0_109_329 ();
 sg13g2_fill_2 FILLER_0_109_339 ();
 sg13g2_fill_1 FILLER_0_109_345 ();
 sg13g2_fill_1 FILLER_0_109_356 ();
 sg13g2_fill_1 FILLER_0_109_367 ();
 sg13g2_fill_2 FILLER_0_109_372 ();
 sg13g2_decap_8 FILLER_0_109_419 ();
 sg13g2_fill_4 FILLER_0_109_430 ();
 sg13g2_fill_8 FILLER_0_109_438 ();
 sg13g2_fill_2 FILLER_0_109_446 ();
 sg13g2_fill_1 FILLER_0_109_458 ();
 sg13g2_fill_4 FILLER_0_109_469 ();
 sg13g2_fill_2 FILLER_0_109_477 ();
 sg13g2_fill_1 FILLER_0_109_479 ();
 sg13g2_fill_8 FILLER_0_109_488 ();
 sg13g2_fill_8 FILLER_0_109_558 ();
 sg13g2_fill_2 FILLER_0_109_566 ();
 sg13g2_fill_1 FILLER_0_109_568 ();
 sg13g2_fill_8 FILLER_0_109_615 ();
 sg13g2_fill_2 FILLER_0_109_623 ();
 sg13g2_fill_8 FILLER_0_109_630 ();
 sg13g2_fill_2 FILLER_0_109_638 ();
 sg13g2_fill_4 FILLER_0_109_681 ();
 sg13g2_fill_2 FILLER_0_109_685 ();
 sg13g2_fill_2 FILLER_0_109_739 ();
 sg13g2_fill_1 FILLER_0_109_741 ();
 sg13g2_fill_2 FILLER_0_109_776 ();
 sg13g2_fill_1 FILLER_0_109_778 ();
 sg13g2_fill_8 FILLER_0_109_783 ();
 sg13g2_fill_8 FILLER_0_109_791 ();
 sg13g2_fill_8 FILLER_0_109_799 ();
 sg13g2_fill_8 FILLER_0_109_807 ();
 sg13g2_fill_8 FILLER_0_109_815 ();
 sg13g2_fill_8 FILLER_0_109_823 ();
 sg13g2_fill_8 FILLER_0_109_831 ();
 sg13g2_decap_8 FILLER_0_109_839 ();
 sg13g2_fill_1 FILLER_0_109_881 ();
 sg13g2_fill_2 FILLER_0_109_887 ();
 sg13g2_fill_1 FILLER_0_109_889 ();
 sg13g2_fill_8 FILLER_0_109_899 ();
 sg13g2_fill_1 FILLER_0_109_907 ();
 sg13g2_fill_2 FILLER_0_109_923 ();
 sg13g2_fill_1 FILLER_0_109_925 ();
 sg13g2_fill_4 FILLER_0_109_934 ();
 sg13g2_fill_2 FILLER_0_109_938 ();
 sg13g2_fill_2 FILLER_0_109_945 ();
 sg13g2_fill_1 FILLER_0_109_947 ();
 sg13g2_fill_2 FILLER_0_109_952 ();
 sg13g2_fill_8 FILLER_0_109_959 ();
 sg13g2_fill_8 FILLER_0_109_967 ();
 sg13g2_fill_8 FILLER_0_109_983 ();
 sg13g2_fill_2 FILLER_0_109_996 ();
 sg13g2_fill_8 FILLER_0_109_1003 ();
 sg13g2_fill_8 FILLER_0_109_1011 ();
 sg13g2_fill_8 FILLER_0_109_1019 ();
 sg13g2_fill_4 FILLER_0_109_1027 ();
 sg13g2_fill_2 FILLER_0_109_1044 ();
 sg13g2_fill_1 FILLER_0_109_1050 ();
 sg13g2_fill_4 FILLER_0_109_1060 ();
 sg13g2_fill_1 FILLER_0_109_1064 ();
 sg13g2_fill_8 FILLER_0_109_1069 ();
 sg13g2_fill_2 FILLER_0_109_1077 ();
 sg13g2_fill_2 FILLER_0_109_1093 ();
 sg13g2_fill_1 FILLER_0_109_1095 ();
 sg13g2_fill_8 FILLER_0_109_1118 ();
 sg13g2_fill_1 FILLER_0_109_1126 ();
 sg13g2_fill_1 FILLER_0_109_1134 ();
 sg13g2_fill_4 FILLER_0_109_1140 ();
 sg13g2_fill_4 FILLER_0_109_1148 ();
 sg13g2_fill_4 FILLER_0_109_1156 ();
 sg13g2_fill_2 FILLER_0_109_1160 ();
 sg13g2_fill_2 FILLER_0_109_1170 ();
 sg13g2_fill_1 FILLER_0_109_1172 ();
 sg13g2_fill_4 FILLER_0_109_1193 ();
 sg13g2_fill_1 FILLER_0_109_1197 ();
 sg13g2_fill_1 FILLER_0_109_1207 ();
 sg13g2_fill_2 FILLER_0_109_1217 ();
 sg13g2_fill_1 FILLER_0_109_1219 ();
 sg13g2_fill_4 FILLER_0_109_1224 ();
 sg13g2_fill_4 FILLER_0_110_0 ();
 sg13g2_fill_1 FILLER_0_110_12 ();
 sg13g2_fill_1 FILLER_0_110_23 ();
 sg13g2_fill_2 FILLER_0_110_50 ();
 sg13g2_fill_1 FILLER_0_110_93 ();
 sg13g2_fill_1 FILLER_0_110_98 ();
 sg13g2_fill_4 FILLER_0_110_109 ();
 sg13g2_fill_2 FILLER_0_110_113 ();
 sg13g2_fill_2 FILLER_0_110_130 ();
 sg13g2_fill_2 FILLER_0_110_140 ();
 sg13g2_fill_1 FILLER_0_110_142 ();
 sg13g2_fill_4 FILLER_0_110_169 ();
 sg13g2_fill_2 FILLER_0_110_173 ();
 sg13g2_fill_1 FILLER_0_110_189 ();
 sg13g2_fill_1 FILLER_0_110_216 ();
 sg13g2_fill_1 FILLER_0_110_227 ();
 sg13g2_fill_1 FILLER_0_110_269 ();
 sg13g2_fill_8 FILLER_0_110_301 ();
 sg13g2_fill_8 FILLER_0_110_309 ();
 sg13g2_fill_8 FILLER_0_110_317 ();
 sg13g2_fill_4 FILLER_0_110_325 ();
 sg13g2_fill_2 FILLER_0_110_333 ();
 sg13g2_fill_1 FILLER_0_110_335 ();
 sg13g2_fill_8 FILLER_0_110_345 ();
 sg13g2_fill_8 FILLER_0_110_353 ();
 sg13g2_fill_8 FILLER_0_110_361 ();
 sg13g2_decap_8 FILLER_0_110_369 ();
 sg13g2_fill_2 FILLER_0_110_380 ();
 sg13g2_fill_1 FILLER_0_110_382 ();
 sg13g2_fill_2 FILLER_0_110_393 ();
 sg13g2_fill_2 FILLER_0_110_404 ();
 sg13g2_fill_1 FILLER_0_110_406 ();
 sg13g2_fill_1 FILLER_0_110_433 ();
 sg13g2_fill_1 FILLER_0_110_447 ();
 sg13g2_decap_8 FILLER_0_110_474 ();
 sg13g2_fill_2 FILLER_0_110_540 ();
 sg13g2_fill_8 FILLER_0_110_546 ();
 sg13g2_fill_8 FILLER_0_110_554 ();
 sg13g2_fill_8 FILLER_0_110_562 ();
 sg13g2_fill_2 FILLER_0_110_570 ();
 sg13g2_fill_8 FILLER_0_110_577 ();
 sg13g2_fill_1 FILLER_0_110_585 ();
 sg13g2_fill_4 FILLER_0_110_590 ();
 sg13g2_fill_1 FILLER_0_110_594 ();
 sg13g2_fill_1 FILLER_0_110_600 ();
 sg13g2_fill_2 FILLER_0_110_627 ();
 sg13g2_fill_4 FILLER_0_110_660 ();
 sg13g2_fill_2 FILLER_0_110_664 ();
 sg13g2_fill_1 FILLER_0_110_697 ();
 sg13g2_fill_1 FILLER_0_110_729 ();
 sg13g2_fill_1 FILLER_0_110_740 ();
 sg13g2_fill_1 FILLER_0_110_756 ();
 sg13g2_fill_4 FILLER_0_110_761 ();
 sg13g2_fill_2 FILLER_0_110_765 ();
 sg13g2_fill_1 FILLER_0_110_808 ();
 sg13g2_fill_8 FILLER_0_110_822 ();
 sg13g2_fill_8 FILLER_0_110_830 ();
 sg13g2_fill_8 FILLER_0_110_838 ();
 sg13g2_fill_8 FILLER_0_110_846 ();
 sg13g2_fill_4 FILLER_0_110_854 ();
 sg13g2_fill_4 FILLER_0_110_862 ();
 sg13g2_fill_1 FILLER_0_110_879 ();
 sg13g2_fill_1 FILLER_0_110_889 ();
 sg13g2_fill_1 FILLER_0_110_895 ();
 sg13g2_fill_1 FILLER_0_110_914 ();
 sg13g2_fill_2 FILLER_0_110_920 ();
 sg13g2_fill_1 FILLER_0_110_927 ();
 sg13g2_fill_2 FILLER_0_110_932 ();
 sg13g2_fill_1 FILLER_0_110_942 ();
 sg13g2_fill_2 FILLER_0_110_948 ();
 sg13g2_fill_1 FILLER_0_110_950 ();
 sg13g2_fill_2 FILLER_0_110_966 ();
 sg13g2_fill_2 FILLER_0_110_978 ();
 sg13g2_fill_1 FILLER_0_110_980 ();
 sg13g2_fill_1 FILLER_0_110_985 ();
 sg13g2_fill_2 FILLER_0_110_1015 ();
 sg13g2_fill_1 FILLER_0_110_1017 ();
 sg13g2_fill_1 FILLER_0_110_1040 ();
 sg13g2_fill_1 FILLER_0_110_1046 ();
 sg13g2_fill_1 FILLER_0_110_1052 ();
 sg13g2_fill_1 FILLER_0_110_1058 ();
 sg13g2_fill_1 FILLER_0_110_1069 ();
 sg13g2_fill_8 FILLER_0_110_1080 ();
 sg13g2_fill_4 FILLER_0_110_1088 ();
 sg13g2_fill_2 FILLER_0_110_1092 ();
 sg13g2_fill_8 FILLER_0_110_1099 ();
 sg13g2_fill_2 FILLER_0_110_1107 ();
 sg13g2_decap_8 FILLER_0_110_1113 ();
 sg13g2_fill_4 FILLER_0_110_1136 ();
 sg13g2_fill_2 FILLER_0_110_1140 ();
 sg13g2_fill_1 FILLER_0_110_1150 ();
 sg13g2_fill_8 FILLER_0_110_1164 ();
 sg13g2_decap_8 FILLER_0_110_1172 ();
 sg13g2_fill_2 FILLER_0_110_1183 ();
 sg13g2_fill_1 FILLER_0_110_1185 ();
 sg13g2_fill_4 FILLER_0_110_1190 ();
 sg13g2_fill_4 FILLER_0_110_1223 ();
 sg13g2_fill_1 FILLER_0_110_1227 ();
 sg13g2_fill_8 FILLER_0_111_0 ();
 sg13g2_fill_4 FILLER_0_111_8 ();
 sg13g2_fill_2 FILLER_0_111_12 ();
 sg13g2_fill_8 FILLER_0_111_19 ();
 sg13g2_fill_4 FILLER_0_111_27 ();
 sg13g2_fill_2 FILLER_0_111_31 ();
 sg13g2_decap_8 FILLER_0_111_37 ();
 sg13g2_fill_1 FILLER_0_111_48 ();
 sg13g2_fill_4 FILLER_0_111_54 ();
 sg13g2_fill_1 FILLER_0_111_58 ();
 sg13g2_fill_1 FILLER_0_111_69 ();
 sg13g2_fill_8 FILLER_0_111_79 ();
 sg13g2_fill_4 FILLER_0_111_87 ();
 sg13g2_fill_2 FILLER_0_111_91 ();
 sg13g2_fill_8 FILLER_0_111_112 ();
 sg13g2_fill_8 FILLER_0_111_120 ();
 sg13g2_fill_4 FILLER_0_111_128 ();
 sg13g2_fill_4 FILLER_0_111_140 ();
 sg13g2_fill_4 FILLER_0_111_148 ();
 sg13g2_fill_8 FILLER_0_111_156 ();
 sg13g2_fill_8 FILLER_0_111_164 ();
 sg13g2_fill_8 FILLER_0_111_172 ();
 sg13g2_fill_1 FILLER_0_111_180 ();
 sg13g2_fill_2 FILLER_0_111_190 ();
 sg13g2_fill_2 FILLER_0_111_197 ();
 sg13g2_fill_8 FILLER_0_111_203 ();
 sg13g2_fill_1 FILLER_0_111_211 ();
 sg13g2_fill_4 FILLER_0_111_217 ();
 sg13g2_fill_1 FILLER_0_111_221 ();
 sg13g2_fill_8 FILLER_0_111_256 ();
 sg13g2_fill_8 FILLER_0_111_264 ();
 sg13g2_fill_8 FILLER_0_111_272 ();
 sg13g2_fill_2 FILLER_0_111_280 ();
 sg13g2_fill_2 FILLER_0_111_296 ();
 sg13g2_fill_2 FILLER_0_111_333 ();
 sg13g2_fill_1 FILLER_0_111_335 ();
 sg13g2_fill_8 FILLER_0_111_362 ();
 sg13g2_fill_8 FILLER_0_111_370 ();
 sg13g2_fill_2 FILLER_0_111_378 ();
 sg13g2_fill_8 FILLER_0_111_407 ();
 sg13g2_fill_8 FILLER_0_111_415 ();
 sg13g2_fill_1 FILLER_0_111_423 ();
 sg13g2_fill_2 FILLER_0_111_459 ();
 sg13g2_fill_2 FILLER_0_111_487 ();
 sg13g2_fill_1 FILLER_0_111_489 ();
 sg13g2_fill_8 FILLER_0_111_525 ();
 sg13g2_fill_8 FILLER_0_111_533 ();
 sg13g2_fill_4 FILLER_0_111_541 ();
 sg13g2_fill_4 FILLER_0_111_550 ();
 sg13g2_fill_1 FILLER_0_111_554 ();
 sg13g2_fill_8 FILLER_0_111_560 ();
 sg13g2_fill_8 FILLER_0_111_568 ();
 sg13g2_fill_8 FILLER_0_111_576 ();
 sg13g2_fill_4 FILLER_0_111_584 ();
 sg13g2_fill_1 FILLER_0_111_588 ();
 sg13g2_fill_1 FILLER_0_111_607 ();
 sg13g2_fill_8 FILLER_0_111_616 ();
 sg13g2_fill_4 FILLER_0_111_624 ();
 sg13g2_fill_1 FILLER_0_111_628 ();
 sg13g2_fill_2 FILLER_0_111_670 ();
 sg13g2_fill_8 FILLER_0_111_676 ();
 sg13g2_fill_8 FILLER_0_111_684 ();
 sg13g2_fill_2 FILLER_0_111_692 ();
 sg13g2_fill_1 FILLER_0_111_694 ();
 sg13g2_fill_4 FILLER_0_111_700 ();
 sg13g2_fill_1 FILLER_0_111_704 ();
 sg13g2_fill_8 FILLER_0_111_719 ();
 sg13g2_fill_8 FILLER_0_111_727 ();
 sg13g2_fill_2 FILLER_0_111_735 ();
 sg13g2_fill_8 FILLER_0_111_742 ();
 sg13g2_fill_2 FILLER_0_111_750 ();
 sg13g2_fill_4 FILLER_0_111_762 ();
 sg13g2_fill_4 FILLER_0_111_807 ();
 sg13g2_fill_4 FILLER_0_111_837 ();
 sg13g2_fill_2 FILLER_0_111_845 ();
 sg13g2_fill_1 FILLER_0_111_847 ();
 sg13g2_fill_2 FILLER_0_111_853 ();
 sg13g2_fill_1 FILLER_0_111_855 ();
 sg13g2_fill_4 FILLER_0_111_905 ();
 sg13g2_fill_1 FILLER_0_111_909 ();
 sg13g2_fill_1 FILLER_0_111_943 ();
 sg13g2_fill_1 FILLER_0_111_952 ();
 sg13g2_fill_2 FILLER_0_111_961 ();
 sg13g2_fill_2 FILLER_0_111_971 ();
 sg13g2_fill_1 FILLER_0_111_986 ();
 sg13g2_fill_1 FILLER_0_111_997 ();
 sg13g2_fill_1 FILLER_0_111_1026 ();
 sg13g2_fill_1 FILLER_0_111_1040 ();
 sg13g2_fill_1 FILLER_0_111_1046 ();
 sg13g2_fill_1 FILLER_0_111_1074 ();
 sg13g2_fill_2 FILLER_0_111_1086 ();
 sg13g2_fill_1 FILLER_0_111_1088 ();
 sg13g2_fill_1 FILLER_0_111_1103 ();
 sg13g2_fill_4 FILLER_0_111_1114 ();
 sg13g2_fill_2 FILLER_0_111_1118 ();
 sg13g2_fill_8 FILLER_0_111_1124 ();
 sg13g2_fill_8 FILLER_0_111_1132 ();
 sg13g2_fill_4 FILLER_0_111_1140 ();
 sg13g2_decap_8 FILLER_0_111_1161 ();
 sg13g2_fill_4 FILLER_0_111_1179 ();
 sg13g2_fill_1 FILLER_0_111_1196 ();
 sg13g2_fill_4 FILLER_0_111_1224 ();
 sg13g2_fill_8 FILLER_0_112_0 ();
 sg13g2_fill_8 FILLER_0_112_8 ();
 sg13g2_fill_8 FILLER_0_112_16 ();
 sg13g2_fill_8 FILLER_0_112_24 ();
 sg13g2_fill_8 FILLER_0_112_32 ();
 sg13g2_fill_8 FILLER_0_112_40 ();
 sg13g2_fill_8 FILLER_0_112_48 ();
 sg13g2_fill_8 FILLER_0_112_56 ();
 sg13g2_fill_8 FILLER_0_112_64 ();
 sg13g2_fill_8 FILLER_0_112_72 ();
 sg13g2_fill_1 FILLER_0_112_80 ();
 sg13g2_fill_8 FILLER_0_112_122 ();
 sg13g2_fill_4 FILLER_0_112_130 ();
 sg13g2_fill_2 FILLER_0_112_134 ();
 sg13g2_fill_1 FILLER_0_112_158 ();
 sg13g2_fill_2 FILLER_0_112_182 ();
 sg13g2_fill_1 FILLER_0_112_184 ();
 sg13g2_fill_8 FILLER_0_112_193 ();
 sg13g2_fill_8 FILLER_0_112_201 ();
 sg13g2_fill_1 FILLER_0_112_239 ();
 sg13g2_fill_8 FILLER_0_112_244 ();
 sg13g2_decap_8 FILLER_0_112_252 ();
 sg13g2_fill_1 FILLER_0_112_285 ();
 sg13g2_fill_8 FILLER_0_112_296 ();
 sg13g2_fill_2 FILLER_0_112_304 ();
 sg13g2_fill_1 FILLER_0_112_306 ();
 sg13g2_fill_1 FILLER_0_112_322 ();
 sg13g2_fill_1 FILLER_0_112_349 ();
 sg13g2_fill_2 FILLER_0_112_376 ();
 sg13g2_fill_2 FILLER_0_112_388 ();
 sg13g2_fill_1 FILLER_0_112_390 ();
 sg13g2_fill_1 FILLER_0_112_401 ();
 sg13g2_fill_2 FILLER_0_112_428 ();
 sg13g2_fill_1 FILLER_0_112_430 ();
 sg13g2_fill_1 FILLER_0_112_461 ();
 sg13g2_fill_1 FILLER_0_112_467 ();
 sg13g2_fill_1 FILLER_0_112_503 ();
 sg13g2_decap_8 FILLER_0_112_519 ();
 sg13g2_fill_1 FILLER_0_112_552 ();
 sg13g2_fill_4 FILLER_0_112_594 ();
 sg13g2_fill_1 FILLER_0_112_598 ();
 sg13g2_fill_4 FILLER_0_112_630 ();
 sg13g2_fill_8 FILLER_0_112_639 ();
 sg13g2_fill_8 FILLER_0_112_647 ();
 sg13g2_fill_8 FILLER_0_112_655 ();
 sg13g2_fill_8 FILLER_0_112_663 ();
 sg13g2_fill_8 FILLER_0_112_679 ();
 sg13g2_fill_2 FILLER_0_112_687 ();
 sg13g2_fill_2 FILLER_0_112_725 ();
 sg13g2_fill_1 FILLER_0_112_727 ();
 sg13g2_fill_1 FILLER_0_112_732 ();
 sg13g2_fill_1 FILLER_0_112_759 ();
 sg13g2_fill_2 FILLER_0_112_795 ();
 sg13g2_fill_1 FILLER_0_112_797 ();
 sg13g2_fill_1 FILLER_0_112_808 ();
 sg13g2_fill_1 FILLER_0_112_835 ();
 sg13g2_fill_4 FILLER_0_112_866 ();
 sg13g2_fill_4 FILLER_0_112_879 ();
 sg13g2_fill_4 FILLER_0_112_914 ();
 sg13g2_fill_2 FILLER_0_112_928 ();
 sg13g2_fill_2 FILLER_0_112_940 ();
 sg13g2_fill_2 FILLER_0_112_957 ();
 sg13g2_decap_8 FILLER_0_112_964 ();
 sg13g2_fill_1 FILLER_0_112_986 ();
 sg13g2_fill_1 FILLER_0_112_992 ();
 sg13g2_fill_1 FILLER_0_112_999 ();
 sg13g2_fill_4 FILLER_0_112_1008 ();
 sg13g2_fill_2 FILLER_0_112_1023 ();
 sg13g2_fill_1 FILLER_0_112_1025 ();
 sg13g2_fill_2 FILLER_0_112_1031 ();
 sg13g2_fill_8 FILLER_0_112_1041 ();
 sg13g2_fill_2 FILLER_0_112_1049 ();
 sg13g2_fill_1 FILLER_0_112_1051 ();
 sg13g2_fill_2 FILLER_0_112_1057 ();
 sg13g2_fill_1 FILLER_0_112_1059 ();
 sg13g2_fill_2 FILLER_0_112_1068 ();
 sg13g2_fill_1 FILLER_0_112_1070 ();
 sg13g2_fill_2 FILLER_0_112_1088 ();
 sg13g2_fill_2 FILLER_0_112_1120 ();
 sg13g2_fill_1 FILLER_0_112_1122 ();
 sg13g2_fill_2 FILLER_0_112_1127 ();
 sg13g2_fill_1 FILLER_0_112_1129 ();
 sg13g2_fill_1 FILLER_0_112_1154 ();
 sg13g2_fill_1 FILLER_0_112_1161 ();
 sg13g2_fill_8 FILLER_0_112_1166 ();
 sg13g2_fill_8 FILLER_0_112_1174 ();
 sg13g2_fill_4 FILLER_0_112_1182 ();
 sg13g2_fill_1 FILLER_0_112_1186 ();
 sg13g2_fill_2 FILLER_0_112_1196 ();
 sg13g2_fill_1 FILLER_0_112_1198 ();
 sg13g2_fill_4 FILLER_0_112_1222 ();
 sg13g2_fill_2 FILLER_0_112_1226 ();
 sg13g2_fill_8 FILLER_0_113_0 ();
 sg13g2_fill_8 FILLER_0_113_8 ();
 sg13g2_fill_8 FILLER_0_113_16 ();
 sg13g2_fill_8 FILLER_0_113_24 ();
 sg13g2_fill_8 FILLER_0_113_32 ();
 sg13g2_fill_8 FILLER_0_113_40 ();
 sg13g2_fill_8 FILLER_0_113_48 ();
 sg13g2_fill_8 FILLER_0_113_56 ();
 sg13g2_fill_8 FILLER_0_113_64 ();
 sg13g2_fill_4 FILLER_0_113_72 ();
 sg13g2_fill_2 FILLER_0_113_76 ();
 sg13g2_fill_2 FILLER_0_113_104 ();
 sg13g2_fill_1 FILLER_0_113_106 ();
 sg13g2_fill_4 FILLER_0_113_117 ();
 sg13g2_fill_1 FILLER_0_113_121 ();
 sg13g2_fill_1 FILLER_0_113_127 ();
 sg13g2_fill_2 FILLER_0_113_142 ();
 sg13g2_fill_1 FILLER_0_113_144 ();
 sg13g2_fill_1 FILLER_0_113_171 ();
 sg13g2_fill_1 FILLER_0_113_198 ();
 sg13g2_decap_8 FILLER_0_113_203 ();
 sg13g2_fill_8 FILLER_0_113_220 ();
 sg13g2_fill_8 FILLER_0_113_228 ();
 sg13g2_fill_8 FILLER_0_113_236 ();
 sg13g2_fill_4 FILLER_0_113_244 ();
 sg13g2_fill_8 FILLER_0_113_252 ();
 sg13g2_fill_2 FILLER_0_113_260 ();
 sg13g2_fill_4 FILLER_0_113_324 ();
 sg13g2_fill_2 FILLER_0_113_338 ();
 sg13g2_fill_2 FILLER_0_113_386 ();
 sg13g2_fill_8 FILLER_0_113_423 ();
 sg13g2_fill_4 FILLER_0_113_431 ();
 sg13g2_fill_2 FILLER_0_113_435 ();
 sg13g2_fill_1 FILLER_0_113_446 ();
 sg13g2_fill_2 FILLER_0_113_457 ();
 sg13g2_fill_8 FILLER_0_113_469 ();
 sg13g2_fill_1 FILLER_0_113_477 ();
 sg13g2_fill_1 FILLER_0_113_497 ();
 sg13g2_fill_8 FILLER_0_113_506 ();
 sg13g2_fill_8 FILLER_0_113_514 ();
 sg13g2_fill_4 FILLER_0_113_522 ();
 sg13g2_fill_1 FILLER_0_113_567 ();
 sg13g2_fill_8 FILLER_0_113_604 ();
 sg13g2_fill_2 FILLER_0_113_612 ();
 sg13g2_fill_1 FILLER_0_113_618 ();
 sg13g2_fill_1 FILLER_0_113_623 ();
 sg13g2_fill_2 FILLER_0_113_629 ();
 sg13g2_fill_8 FILLER_0_113_645 ();
 sg13g2_fill_1 FILLER_0_113_653 ();
 sg13g2_fill_4 FILLER_0_113_724 ();
 sg13g2_fill_1 FILLER_0_113_728 ();
 sg13g2_fill_1 FILLER_0_113_737 ();
 sg13g2_fill_2 FILLER_0_113_774 ();
 sg13g2_fill_8 FILLER_0_113_786 ();
 sg13g2_fill_2 FILLER_0_113_804 ();
 sg13g2_fill_1 FILLER_0_113_806 ();
 sg13g2_fill_2 FILLER_0_113_812 ();
 sg13g2_fill_1 FILLER_0_113_814 ();
 sg13g2_fill_2 FILLER_0_113_819 ();
 sg13g2_fill_1 FILLER_0_113_821 ();
 sg13g2_fill_8 FILLER_0_113_826 ();
 sg13g2_fill_2 FILLER_0_113_838 ();
 sg13g2_decap_8 FILLER_0_113_866 ();
 sg13g2_fill_8 FILLER_0_113_878 ();
 sg13g2_fill_4 FILLER_0_113_886 ();
 sg13g2_fill_1 FILLER_0_113_890 ();
 sg13g2_fill_4 FILLER_0_113_899 ();
 sg13g2_fill_8 FILLER_0_113_922 ();
 sg13g2_fill_1 FILLER_0_113_930 ();
 sg13g2_fill_8 FILLER_0_113_934 ();
 sg13g2_fill_4 FILLER_0_113_942 ();
 sg13g2_fill_1 FILLER_0_113_946 ();
 sg13g2_fill_1 FILLER_0_113_959 ();
 sg13g2_fill_8 FILLER_0_113_965 ();
 sg13g2_fill_2 FILLER_0_113_973 ();
 sg13g2_fill_8 FILLER_0_113_980 ();
 sg13g2_fill_2 FILLER_0_113_988 ();
 sg13g2_fill_1 FILLER_0_113_990 ();
 sg13g2_fill_8 FILLER_0_113_1000 ();
 sg13g2_fill_8 FILLER_0_113_1008 ();
 sg13g2_fill_8 FILLER_0_113_1035 ();
 sg13g2_fill_8 FILLER_0_113_1043 ();
 sg13g2_fill_4 FILLER_0_113_1051 ();
 sg13g2_fill_4 FILLER_0_113_1058 ();
 sg13g2_fill_2 FILLER_0_113_1062 ();
 sg13g2_fill_2 FILLER_0_113_1068 ();
 sg13g2_fill_1 FILLER_0_113_1091 ();
 sg13g2_fill_4 FILLER_0_113_1101 ();
 sg13g2_fill_2 FILLER_0_113_1121 ();
 sg13g2_fill_8 FILLER_0_113_1131 ();
 sg13g2_fill_1 FILLER_0_113_1159 ();
 sg13g2_fill_1 FILLER_0_113_1165 ();
 sg13g2_fill_1 FILLER_0_113_1171 ();
 sg13g2_fill_1 FILLER_0_113_1200 ();
 sg13g2_fill_8 FILLER_0_113_1208 ();
 sg13g2_fill_8 FILLER_0_113_1216 ();
 sg13g2_fill_4 FILLER_0_113_1224 ();
 sg13g2_fill_8 FILLER_0_114_0 ();
 sg13g2_fill_8 FILLER_0_114_8 ();
 sg13g2_fill_8 FILLER_0_114_16 ();
 sg13g2_fill_8 FILLER_0_114_24 ();
 sg13g2_fill_8 FILLER_0_114_32 ();
 sg13g2_fill_8 FILLER_0_114_40 ();
 sg13g2_fill_8 FILLER_0_114_48 ();
 sg13g2_fill_8 FILLER_0_114_56 ();
 sg13g2_fill_8 FILLER_0_114_64 ();
 sg13g2_fill_1 FILLER_0_114_72 ();
 sg13g2_fill_1 FILLER_0_114_179 ();
 sg13g2_fill_1 FILLER_0_114_190 ();
 sg13g2_fill_2 FILLER_0_114_222 ();
 sg13g2_fill_1 FILLER_0_114_224 ();
 sg13g2_fill_1 FILLER_0_114_235 ();
 sg13g2_fill_2 FILLER_0_114_240 ();
 sg13g2_decap_8 FILLER_0_114_257 ();
 sg13g2_fill_4 FILLER_0_114_294 ();
 sg13g2_fill_2 FILLER_0_114_298 ();
 sg13g2_fill_1 FILLER_0_114_351 ();
 sg13g2_fill_2 FILLER_0_114_402 ();
 sg13g2_fill_8 FILLER_0_114_408 ();
 sg13g2_fill_8 FILLER_0_114_416 ();
 sg13g2_decap_8 FILLER_0_114_424 ();
 sg13g2_fill_8 FILLER_0_114_441 ();
 sg13g2_fill_8 FILLER_0_114_449 ();
 sg13g2_fill_8 FILLER_0_114_457 ();
 sg13g2_fill_4 FILLER_0_114_465 ();
 sg13g2_fill_2 FILLER_0_114_469 ();
 sg13g2_fill_8 FILLER_0_114_481 ();
 sg13g2_fill_8 FILLER_0_114_489 ();
 sg13g2_fill_8 FILLER_0_114_497 ();
 sg13g2_fill_8 FILLER_0_114_505 ();
 sg13g2_fill_8 FILLER_0_114_513 ();
 sg13g2_fill_2 FILLER_0_114_521 ();
 sg13g2_fill_1 FILLER_0_114_553 ();
 sg13g2_fill_1 FILLER_0_114_564 ();
 sg13g2_fill_1 FILLER_0_114_621 ();
 sg13g2_fill_8 FILLER_0_114_648 ();
 sg13g2_fill_1 FILLER_0_114_656 ();
 sg13g2_fill_1 FILLER_0_114_661 ();
 sg13g2_fill_1 FILLER_0_114_667 ();
 sg13g2_fill_2 FILLER_0_114_678 ();
 sg13g2_fill_1 FILLER_0_114_680 ();
 sg13g2_fill_8 FILLER_0_114_691 ();
 sg13g2_decap_8 FILLER_0_114_699 ();
 sg13g2_fill_2 FILLER_0_114_710 ();
 sg13g2_fill_1 FILLER_0_114_712 ();
 sg13g2_fill_1 FILLER_0_114_731 ();
 sg13g2_fill_2 FILLER_0_114_751 ();
 sg13g2_fill_1 FILLER_0_114_753 ();
 sg13g2_fill_4 FILLER_0_114_764 ();
 sg13g2_fill_1 FILLER_0_114_768 ();
 sg13g2_fill_8 FILLER_0_114_773 ();
 sg13g2_fill_8 FILLER_0_114_781 ();
 sg13g2_fill_8 FILLER_0_114_789 ();
 sg13g2_fill_8 FILLER_0_114_828 ();
 sg13g2_fill_2 FILLER_0_114_871 ();
 sg13g2_fill_1 FILLER_0_114_877 ();
 sg13g2_fill_4 FILLER_0_114_883 ();
 sg13g2_decap_8 FILLER_0_114_916 ();
 sg13g2_fill_1 FILLER_0_114_927 ();
 sg13g2_fill_4 FILLER_0_114_931 ();
 sg13g2_fill_2 FILLER_0_114_935 ();
 sg13g2_fill_4 FILLER_0_114_950 ();
 sg13g2_fill_2 FILLER_0_114_954 ();
 sg13g2_fill_1 FILLER_0_114_961 ();
 sg13g2_fill_2 FILLER_0_114_967 ();
 sg13g2_fill_4 FILLER_0_114_974 ();
 sg13g2_fill_8 FILLER_0_114_982 ();
 sg13g2_fill_8 FILLER_0_114_990 ();
 sg13g2_fill_8 FILLER_0_114_998 ();
 sg13g2_fill_8 FILLER_0_114_1006 ();
 sg13g2_fill_4 FILLER_0_114_1014 ();
 sg13g2_fill_1 FILLER_0_114_1018 ();
 sg13g2_fill_1 FILLER_0_114_1027 ();
 sg13g2_fill_1 FILLER_0_114_1037 ();
 sg13g2_fill_8 FILLER_0_114_1043 ();
 sg13g2_decap_8 FILLER_0_114_1051 ();
 sg13g2_fill_8 FILLER_0_114_1069 ();
 sg13g2_fill_8 FILLER_0_114_1077 ();
 sg13g2_fill_1 FILLER_0_114_1085 ();
 sg13g2_fill_1 FILLER_0_114_1095 ();
 sg13g2_fill_4 FILLER_0_114_1102 ();
 sg13g2_fill_1 FILLER_0_114_1114 ();
 sg13g2_fill_1 FILLER_0_114_1122 ();
 sg13g2_fill_4 FILLER_0_114_1128 ();
 sg13g2_fill_1 FILLER_0_114_1132 ();
 sg13g2_fill_2 FILLER_0_114_1138 ();
 sg13g2_fill_1 FILLER_0_114_1140 ();
 sg13g2_fill_2 FILLER_0_114_1146 ();
 sg13g2_fill_1 FILLER_0_114_1148 ();
 sg13g2_fill_2 FILLER_0_114_1167 ();
 sg13g2_fill_2 FILLER_0_114_1179 ();
 sg13g2_fill_1 FILLER_0_114_1181 ();
 sg13g2_fill_1 FILLER_0_114_1190 ();
 sg13g2_fill_1 FILLER_0_114_1211 ();
 sg13g2_fill_8 FILLER_0_114_1217 ();
 sg13g2_fill_2 FILLER_0_114_1225 ();
 sg13g2_fill_1 FILLER_0_114_1227 ();
 sg13g2_fill_8 FILLER_0_115_0 ();
 sg13g2_fill_8 FILLER_0_115_8 ();
 sg13g2_fill_8 FILLER_0_115_16 ();
 sg13g2_fill_8 FILLER_0_115_24 ();
 sg13g2_fill_8 FILLER_0_115_32 ();
 sg13g2_fill_8 FILLER_0_115_40 ();
 sg13g2_fill_8 FILLER_0_115_48 ();
 sg13g2_fill_8 FILLER_0_115_56 ();
 sg13g2_fill_8 FILLER_0_115_64 ();
 sg13g2_fill_8 FILLER_0_115_72 ();
 sg13g2_fill_1 FILLER_0_115_84 ();
 sg13g2_fill_1 FILLER_0_115_89 ();
 sg13g2_fill_2 FILLER_0_115_117 ();
 sg13g2_fill_1 FILLER_0_115_145 ();
 sg13g2_fill_1 FILLER_0_115_156 ();
 sg13g2_fill_2 FILLER_0_115_183 ();
 sg13g2_fill_2 FILLER_0_115_189 ();
 sg13g2_fill_2 FILLER_0_115_195 ();
 sg13g2_fill_1 FILLER_0_115_197 ();
 sg13g2_fill_2 FILLER_0_115_202 ();
 sg13g2_fill_4 FILLER_0_115_300 ();
 sg13g2_fill_1 FILLER_0_115_304 ();
 sg13g2_fill_8 FILLER_0_115_331 ();
 sg13g2_fill_8 FILLER_0_115_339 ();
 sg13g2_fill_8 FILLER_0_115_347 ();
 sg13g2_fill_4 FILLER_0_115_355 ();
 sg13g2_fill_1 FILLER_0_115_359 ();
 sg13g2_fill_2 FILLER_0_115_365 ();
 sg13g2_fill_4 FILLER_0_115_371 ();
 sg13g2_fill_2 FILLER_0_115_375 ();
 sg13g2_decap_8 FILLER_0_115_390 ();
 sg13g2_fill_8 FILLER_0_115_401 ();
 sg13g2_fill_4 FILLER_0_115_409 ();
 sg13g2_fill_2 FILLER_0_115_413 ();
 sg13g2_fill_2 FILLER_0_115_420 ();
 sg13g2_fill_1 FILLER_0_115_422 ();
 sg13g2_fill_8 FILLER_0_115_464 ();
 sg13g2_fill_4 FILLER_0_115_472 ();
 sg13g2_fill_8 FILLER_0_115_502 ();
 sg13g2_fill_8 FILLER_0_115_510 ();
 sg13g2_fill_2 FILLER_0_115_518 ();
 sg13g2_fill_1 FILLER_0_115_520 ();
 sg13g2_fill_8 FILLER_0_115_525 ();
 sg13g2_fill_8 FILLER_0_115_533 ();
 sg13g2_fill_8 FILLER_0_115_541 ();
 sg13g2_fill_8 FILLER_0_115_549 ();
 sg13g2_fill_4 FILLER_0_115_557 ();
 sg13g2_fill_1 FILLER_0_115_561 ();
 sg13g2_fill_8 FILLER_0_115_566 ();
 sg13g2_fill_1 FILLER_0_115_583 ();
 sg13g2_fill_2 FILLER_0_115_611 ();
 sg13g2_fill_1 FILLER_0_115_618 ();
 sg13g2_fill_8 FILLER_0_115_633 ();
 sg13g2_fill_4 FILLER_0_115_641 ();
 sg13g2_fill_8 FILLER_0_115_745 ();
 sg13g2_fill_2 FILLER_0_115_753 ();
 sg13g2_fill_1 FILLER_0_115_755 ();
 sg13g2_fill_4 FILLER_0_115_760 ();
 sg13g2_fill_2 FILLER_0_115_764 ();
 sg13g2_fill_1 FILLER_0_115_801 ();
 sg13g2_fill_2 FILLER_0_115_806 ();
 sg13g2_fill_1 FILLER_0_115_808 ();
 sg13g2_fill_8 FILLER_0_115_813 ();
 sg13g2_fill_8 FILLER_0_115_821 ();
 sg13g2_fill_8 FILLER_0_115_829 ();
 sg13g2_fill_8 FILLER_0_115_837 ();
 sg13g2_decap_8 FILLER_0_115_845 ();
 sg13g2_decap_8 FILLER_0_115_856 ();
 sg13g2_fill_1 FILLER_0_115_887 ();
 sg13g2_fill_8 FILLER_0_115_898 ();
 sg13g2_fill_1 FILLER_0_115_906 ();
 sg13g2_fill_4 FILLER_0_115_916 ();
 sg13g2_fill_2 FILLER_0_115_920 ();
 sg13g2_fill_2 FILLER_0_115_925 ();
 sg13g2_fill_1 FILLER_0_115_953 ();
 sg13g2_fill_2 FILLER_0_115_965 ();
 sg13g2_fill_2 FILLER_0_115_972 ();
 sg13g2_fill_2 FILLER_0_115_984 ();
 sg13g2_fill_1 FILLER_0_115_991 ();
 sg13g2_fill_2 FILLER_0_115_997 ();
 sg13g2_decap_8 FILLER_0_115_1004 ();
 sg13g2_fill_4 FILLER_0_115_1027 ();
 sg13g2_fill_2 FILLER_0_115_1046 ();
 sg13g2_fill_4 FILLER_0_115_1053 ();
 sg13g2_fill_1 FILLER_0_115_1057 ();
 sg13g2_fill_8 FILLER_0_115_1072 ();
 sg13g2_fill_2 FILLER_0_115_1080 ();
 sg13g2_fill_1 FILLER_0_115_1109 ();
 sg13g2_fill_2 FILLER_0_115_1114 ();
 sg13g2_decap_8 FILLER_0_115_1120 ();
 sg13g2_fill_1 FILLER_0_115_1148 ();
 sg13g2_fill_2 FILLER_0_115_1176 ();
 sg13g2_fill_1 FILLER_0_115_1183 ();
 sg13g2_fill_1 FILLER_0_115_1220 ();
 sg13g2_fill_2 FILLER_0_115_1225 ();
 sg13g2_fill_1 FILLER_0_115_1227 ();
 sg13g2_fill_8 FILLER_0_116_0 ();
 sg13g2_fill_8 FILLER_0_116_8 ();
 sg13g2_fill_8 FILLER_0_116_16 ();
 sg13g2_fill_8 FILLER_0_116_24 ();
 sg13g2_fill_8 FILLER_0_116_32 ();
 sg13g2_fill_8 FILLER_0_116_40 ();
 sg13g2_fill_8 FILLER_0_116_48 ();
 sg13g2_fill_8 FILLER_0_116_56 ();
 sg13g2_fill_8 FILLER_0_116_64 ();
 sg13g2_fill_8 FILLER_0_116_72 ();
 sg13g2_fill_8 FILLER_0_116_80 ();
 sg13g2_fill_8 FILLER_0_116_88 ();
 sg13g2_fill_8 FILLER_0_116_96 ();
 sg13g2_fill_8 FILLER_0_116_104 ();
 sg13g2_fill_1 FILLER_0_116_112 ();
 sg13g2_fill_8 FILLER_0_116_118 ();
 sg13g2_fill_2 FILLER_0_116_126 ();
 sg13g2_fill_8 FILLER_0_116_132 ();
 sg13g2_fill_8 FILLER_0_116_140 ();
 sg13g2_fill_4 FILLER_0_116_148 ();
 sg13g2_fill_4 FILLER_0_116_156 ();
 sg13g2_fill_2 FILLER_0_116_179 ();
 sg13g2_fill_2 FILLER_0_116_189 ();
 sg13g2_fill_1 FILLER_0_116_191 ();
 sg13g2_fill_2 FILLER_0_116_249 ();
 sg13g2_fill_2 FILLER_0_116_261 ();
 sg13g2_fill_8 FILLER_0_116_292 ();
 sg13g2_fill_8 FILLER_0_116_300 ();
 sg13g2_fill_8 FILLER_0_116_353 ();
 sg13g2_fill_8 FILLER_0_116_361 ();
 sg13g2_fill_8 FILLER_0_116_369 ();
 sg13g2_fill_8 FILLER_0_116_377 ();
 sg13g2_fill_8 FILLER_0_116_385 ();
 sg13g2_fill_8 FILLER_0_116_393 ();
 sg13g2_fill_4 FILLER_0_116_401 ();
 sg13g2_fill_1 FILLER_0_116_410 ();
 sg13g2_fill_2 FILLER_0_116_416 ();
 sg13g2_fill_2 FILLER_0_116_444 ();
 sg13g2_fill_1 FILLER_0_116_446 ();
 sg13g2_fill_8 FILLER_0_116_499 ();
 sg13g2_fill_2 FILLER_0_116_507 ();
 sg13g2_fill_1 FILLER_0_116_509 ();
 sg13g2_fill_8 FILLER_0_116_551 ();
 sg13g2_decap_8 FILLER_0_116_559 ();
 sg13g2_fill_8 FILLER_0_116_578 ();
 sg13g2_fill_8 FILLER_0_116_586 ();
 sg13g2_fill_4 FILLER_0_116_594 ();
 sg13g2_fill_2 FILLER_0_116_598 ();
 sg13g2_fill_8 FILLER_0_116_604 ();
 sg13g2_fill_8 FILLER_0_116_638 ();
 sg13g2_fill_8 FILLER_0_116_646 ();
 sg13g2_fill_1 FILLER_0_116_654 ();
 sg13g2_fill_4 FILLER_0_116_659 ();
 sg13g2_fill_1 FILLER_0_116_663 ();
 sg13g2_fill_1 FILLER_0_116_686 ();
 sg13g2_fill_8 FILLER_0_116_691 ();
 sg13g2_fill_8 FILLER_0_116_699 ();
 sg13g2_decap_8 FILLER_0_116_707 ();
 sg13g2_fill_2 FILLER_0_116_724 ();
 sg13g2_fill_8 FILLER_0_116_730 ();
 sg13g2_fill_8 FILLER_0_116_738 ();
 sg13g2_decap_8 FILLER_0_116_746 ();
 sg13g2_fill_2 FILLER_0_116_757 ();
 sg13g2_fill_8 FILLER_0_116_816 ();
 sg13g2_fill_8 FILLER_0_116_824 ();
 sg13g2_fill_8 FILLER_0_116_832 ();
 sg13g2_decap_8 FILLER_0_116_840 ();
 sg13g2_fill_4 FILLER_0_116_856 ();
 sg13g2_fill_2 FILLER_0_116_860 ();
 sg13g2_fill_1 FILLER_0_116_871 ();
 sg13g2_fill_2 FILLER_0_116_905 ();
 sg13g2_fill_1 FILLER_0_116_907 ();
 sg13g2_fill_2 FILLER_0_116_920 ();
 sg13g2_fill_1 FILLER_0_116_922 ();
 sg13g2_fill_2 FILLER_0_116_934 ();
 sg13g2_fill_2 FILLER_0_116_940 ();
 sg13g2_fill_2 FILLER_0_116_960 ();
 sg13g2_fill_1 FILLER_0_116_962 ();
 sg13g2_fill_1 FILLER_0_116_977 ();
 sg13g2_fill_1 FILLER_0_116_1007 ();
 sg13g2_fill_8 FILLER_0_116_1016 ();
 sg13g2_fill_1 FILLER_0_116_1024 ();
 sg13g2_fill_1 FILLER_0_116_1034 ();
 sg13g2_fill_2 FILLER_0_116_1039 ();
 sg13g2_fill_1 FILLER_0_116_1046 ();
 sg13g2_fill_1 FILLER_0_116_1055 ();
 sg13g2_fill_1 FILLER_0_116_1060 ();
 sg13g2_fill_2 FILLER_0_116_1066 ();
 sg13g2_fill_4 FILLER_0_116_1081 ();
 sg13g2_fill_1 FILLER_0_116_1085 ();
 sg13g2_fill_1 FILLER_0_116_1097 ();
 sg13g2_fill_1 FILLER_0_116_1102 ();
 sg13g2_fill_1 FILLER_0_116_1110 ();
 sg13g2_fill_1 FILLER_0_116_1124 ();
 sg13g2_fill_2 FILLER_0_116_1130 ();
 sg13g2_fill_2 FILLER_0_116_1142 ();
 sg13g2_fill_1 FILLER_0_116_1144 ();
 sg13g2_fill_4 FILLER_0_116_1182 ();
 sg13g2_fill_1 FILLER_0_116_1186 ();
 sg13g2_fill_1 FILLER_0_116_1191 ();
 sg13g2_decap_8 FILLER_0_116_1196 ();
 sg13g2_fill_1 FILLER_0_116_1210 ();
 sg13g2_fill_8 FILLER_0_116_1219 ();
 sg13g2_fill_1 FILLER_0_116_1227 ();
 sg13g2_fill_8 FILLER_0_117_0 ();
 sg13g2_fill_8 FILLER_0_117_8 ();
 sg13g2_fill_8 FILLER_0_117_16 ();
 sg13g2_fill_8 FILLER_0_117_24 ();
 sg13g2_fill_8 FILLER_0_117_32 ();
 sg13g2_fill_8 FILLER_0_117_40 ();
 sg13g2_fill_8 FILLER_0_117_48 ();
 sg13g2_fill_8 FILLER_0_117_56 ();
 sg13g2_fill_8 FILLER_0_117_64 ();
 sg13g2_fill_8 FILLER_0_117_72 ();
 sg13g2_fill_8 FILLER_0_117_80 ();
 sg13g2_fill_8 FILLER_0_117_88 ();
 sg13g2_fill_8 FILLER_0_117_96 ();
 sg13g2_fill_8 FILLER_0_117_104 ();
 sg13g2_fill_4 FILLER_0_117_112 ();
 sg13g2_fill_2 FILLER_0_117_116 ();
 sg13g2_fill_4 FILLER_0_117_154 ();
 sg13g2_fill_1 FILLER_0_117_158 ();
 sg13g2_fill_4 FILLER_0_117_185 ();
 sg13g2_fill_2 FILLER_0_117_189 ();
 sg13g2_fill_8 FILLER_0_117_196 ();
 sg13g2_fill_1 FILLER_0_117_204 ();
 sg13g2_fill_4 FILLER_0_117_209 ();
 sg13g2_fill_2 FILLER_0_117_213 ();
 sg13g2_fill_8 FILLER_0_117_219 ();
 sg13g2_fill_8 FILLER_0_117_227 ();
 sg13g2_fill_8 FILLER_0_117_300 ();
 sg13g2_fill_8 FILLER_0_117_308 ();
 sg13g2_decap_8 FILLER_0_117_316 ();
 sg13g2_fill_1 FILLER_0_117_338 ();
 sg13g2_fill_2 FILLER_0_117_365 ();
 sg13g2_fill_1 FILLER_0_117_372 ();
 sg13g2_fill_2 FILLER_0_117_383 ();
 sg13g2_fill_1 FILLER_0_117_411 ();
 sg13g2_fill_1 FILLER_0_117_438 ();
 sg13g2_fill_1 FILLER_0_117_443 ();
 sg13g2_fill_1 FILLER_0_117_454 ();
 sg13g2_fill_1 FILLER_0_117_459 ();
 sg13g2_fill_1 FILLER_0_117_470 ();
 sg13g2_fill_1 FILLER_0_117_481 ();
 sg13g2_fill_1 FILLER_0_117_486 ();
 sg13g2_fill_8 FILLER_0_117_491 ();
 sg13g2_fill_8 FILLER_0_117_499 ();
 sg13g2_fill_8 FILLER_0_117_507 ();
 sg13g2_fill_8 FILLER_0_117_515 ();
 sg13g2_fill_8 FILLER_0_117_523 ();
 sg13g2_fill_2 FILLER_0_117_531 ();
 sg13g2_fill_8 FILLER_0_117_543 ();
 sg13g2_fill_8 FILLER_0_117_551 ();
 sg13g2_fill_8 FILLER_0_117_559 ();
 sg13g2_fill_8 FILLER_0_117_603 ();
 sg13g2_fill_2 FILLER_0_117_611 ();
 sg13g2_fill_1 FILLER_0_117_613 ();
 sg13g2_fill_1 FILLER_0_117_622 ();
 sg13g2_fill_8 FILLER_0_117_637 ();
 sg13g2_fill_2 FILLER_0_117_671 ();
 sg13g2_fill_2 FILLER_0_117_678 ();
 sg13g2_fill_1 FILLER_0_117_680 ();
 sg13g2_fill_2 FILLER_0_117_707 ();
 sg13g2_fill_1 FILLER_0_117_709 ();
 sg13g2_fill_2 FILLER_0_117_779 ();
 sg13g2_fill_2 FILLER_0_117_789 ();
 sg13g2_fill_8 FILLER_0_117_817 ();
 sg13g2_decap_8 FILLER_0_117_825 ();
 sg13g2_fill_2 FILLER_0_117_845 ();
 sg13g2_fill_2 FILLER_0_117_862 ();
 sg13g2_fill_1 FILLER_0_117_864 ();
 sg13g2_fill_2 FILLER_0_117_878 ();
 sg13g2_fill_1 FILLER_0_117_880 ();
 sg13g2_fill_2 FILLER_0_117_886 ();
 sg13g2_fill_4 FILLER_0_117_924 ();
 sg13g2_fill_1 FILLER_0_117_934 ();
 sg13g2_fill_2 FILLER_0_117_939 ();
 sg13g2_fill_1 FILLER_0_117_946 ();
 sg13g2_fill_1 FILLER_0_117_957 ();
 sg13g2_fill_1 FILLER_0_117_962 ();
 sg13g2_fill_1 FILLER_0_117_967 ();
 sg13g2_fill_2 FILLER_0_117_972 ();
 sg13g2_fill_2 FILLER_0_117_981 ();
 sg13g2_fill_1 FILLER_0_117_983 ();
 sg13g2_fill_2 FILLER_0_117_997 ();
 sg13g2_fill_2 FILLER_0_117_1003 ();
 sg13g2_fill_2 FILLER_0_117_1037 ();
 sg13g2_fill_1 FILLER_0_117_1039 ();
 sg13g2_fill_1 FILLER_0_117_1102 ();
 sg13g2_fill_1 FILLER_0_117_1108 ();
 sg13g2_fill_8 FILLER_0_117_1122 ();
 sg13g2_fill_8 FILLER_0_117_1130 ();
 sg13g2_fill_8 FILLER_0_117_1138 ();
 sg13g2_fill_4 FILLER_0_117_1146 ();
 sg13g2_fill_1 FILLER_0_117_1150 ();
 sg13g2_fill_2 FILLER_0_117_1176 ();
 sg13g2_decap_8 FILLER_0_117_1183 ();
 sg13g2_fill_2 FILLER_0_117_1194 ();
 sg13g2_fill_8 FILLER_0_117_1201 ();
 sg13g2_fill_8 FILLER_0_117_1209 ();
 sg13g2_fill_8 FILLER_0_117_1217 ();
 sg13g2_fill_2 FILLER_0_117_1225 ();
 sg13g2_fill_1 FILLER_0_117_1227 ();
 sg13g2_fill_8 FILLER_0_118_0 ();
 sg13g2_fill_8 FILLER_0_118_8 ();
 sg13g2_fill_8 FILLER_0_118_16 ();
 sg13g2_fill_8 FILLER_0_118_24 ();
 sg13g2_fill_8 FILLER_0_118_32 ();
 sg13g2_fill_8 FILLER_0_118_40 ();
 sg13g2_fill_8 FILLER_0_118_48 ();
 sg13g2_fill_8 FILLER_0_118_56 ();
 sg13g2_fill_8 FILLER_0_118_64 ();
 sg13g2_fill_8 FILLER_0_118_72 ();
 sg13g2_fill_8 FILLER_0_118_80 ();
 sg13g2_fill_8 FILLER_0_118_88 ();
 sg13g2_fill_8 FILLER_0_118_96 ();
 sg13g2_fill_8 FILLER_0_118_104 ();
 sg13g2_fill_8 FILLER_0_118_112 ();
 sg13g2_fill_4 FILLER_0_118_120 ();
 sg13g2_fill_1 FILLER_0_118_124 ();
 sg13g2_fill_1 FILLER_0_118_170 ();
 sg13g2_fill_4 FILLER_0_118_207 ();
 sg13g2_fill_2 FILLER_0_118_211 ();
 sg13g2_fill_8 FILLER_0_118_228 ();
 sg13g2_fill_1 FILLER_0_118_236 ();
 sg13g2_fill_2 FILLER_0_118_287 ();
 sg13g2_fill_8 FILLER_0_118_293 ();
 sg13g2_fill_8 FILLER_0_118_301 ();
 sg13g2_fill_1 FILLER_0_118_314 ();
 sg13g2_decap_8 FILLER_0_118_349 ();
 sg13g2_fill_2 FILLER_0_118_382 ();
 sg13g2_fill_8 FILLER_0_118_434 ();
 sg13g2_fill_1 FILLER_0_118_442 ();
 sg13g2_fill_8 FILLER_0_118_456 ();
 sg13g2_fill_4 FILLER_0_118_464 ();
 sg13g2_fill_2 FILLER_0_118_468 ();
 sg13g2_fill_8 FILLER_0_118_480 ();
 sg13g2_fill_4 FILLER_0_118_488 ();
 sg13g2_fill_8 FILLER_0_118_496 ();
 sg13g2_fill_2 FILLER_0_118_504 ();
 sg13g2_fill_1 FILLER_0_118_506 ();
 sg13g2_fill_8 FILLER_0_118_515 ();
 sg13g2_fill_4 FILLER_0_118_523 ();
 sg13g2_fill_2 FILLER_0_118_527 ();
 sg13g2_fill_2 FILLER_0_118_575 ();
 sg13g2_fill_1 FILLER_0_118_577 ();
 sg13g2_fill_1 FILLER_0_118_609 ();
 sg13g2_fill_1 FILLER_0_118_649 ();
 sg13g2_fill_2 FILLER_0_118_680 ();
 sg13g2_fill_1 FILLER_0_118_682 ();
 sg13g2_fill_2 FILLER_0_118_728 ();
 sg13g2_fill_1 FILLER_0_118_745 ();
 sg13g2_fill_8 FILLER_0_118_751 ();
 sg13g2_fill_1 FILLER_0_118_759 ();
 sg13g2_fill_4 FILLER_0_118_770 ();
 sg13g2_fill_1 FILLER_0_118_774 ();
 sg13g2_fill_2 FILLER_0_118_872 ();
 sg13g2_fill_1 FILLER_0_118_874 ();
 sg13g2_fill_1 FILLER_0_118_897 ();
 sg13g2_fill_8 FILLER_0_118_908 ();
 sg13g2_fill_2 FILLER_0_118_916 ();
 sg13g2_fill_1 FILLER_0_118_918 ();
 sg13g2_fill_1 FILLER_0_118_937 ();
 sg13g2_fill_4 FILLER_0_118_950 ();
 sg13g2_fill_8 FILLER_0_118_958 ();
 sg13g2_fill_8 FILLER_0_118_966 ();
 sg13g2_fill_8 FILLER_0_118_974 ();
 sg13g2_fill_4 FILLER_0_118_982 ();
 sg13g2_fill_1 FILLER_0_118_986 ();
 sg13g2_fill_2 FILLER_0_118_1018 ();
 sg13g2_fill_1 FILLER_0_118_1020 ();
 sg13g2_fill_4 FILLER_0_118_1030 ();
 sg13g2_fill_2 FILLER_0_118_1034 ();
 sg13g2_fill_1 FILLER_0_118_1065 ();
 sg13g2_fill_4 FILLER_0_118_1083 ();
 sg13g2_fill_2 FILLER_0_118_1092 ();
 sg13g2_fill_2 FILLER_0_118_1098 ();
 sg13g2_fill_4 FILLER_0_118_1115 ();
 sg13g2_fill_8 FILLER_0_118_1126 ();
 sg13g2_fill_8 FILLER_0_118_1134 ();
 sg13g2_decap_8 FILLER_0_118_1142 ();
 sg13g2_fill_2 FILLER_0_118_1166 ();
 sg13g2_fill_1 FILLER_0_118_1168 ();
 sg13g2_fill_4 FILLER_0_118_1174 ();
 sg13g2_fill_2 FILLER_0_118_1183 ();
 sg13g2_fill_1 FILLER_0_118_1185 ();
 sg13g2_fill_1 FILLER_0_118_1200 ();
 sg13g2_fill_2 FILLER_0_118_1205 ();
 sg13g2_fill_8 FILLER_0_118_1219 ();
 sg13g2_fill_1 FILLER_0_118_1227 ();
 sg13g2_fill_8 FILLER_0_119_0 ();
 sg13g2_fill_8 FILLER_0_119_8 ();
 sg13g2_fill_8 FILLER_0_119_16 ();
 sg13g2_fill_8 FILLER_0_119_24 ();
 sg13g2_fill_8 FILLER_0_119_32 ();
 sg13g2_fill_8 FILLER_0_119_40 ();
 sg13g2_fill_8 FILLER_0_119_48 ();
 sg13g2_fill_8 FILLER_0_119_56 ();
 sg13g2_fill_8 FILLER_0_119_64 ();
 sg13g2_fill_8 FILLER_0_119_72 ();
 sg13g2_fill_8 FILLER_0_119_80 ();
 sg13g2_fill_8 FILLER_0_119_88 ();
 sg13g2_fill_8 FILLER_0_119_96 ();
 sg13g2_fill_8 FILLER_0_119_104 ();
 sg13g2_decap_8 FILLER_0_119_112 ();
 sg13g2_fill_2 FILLER_0_119_155 ();
 sg13g2_fill_2 FILLER_0_119_162 ();
 sg13g2_fill_1 FILLER_0_119_164 ();
 sg13g2_fill_1 FILLER_0_119_234 ();
 sg13g2_fill_2 FILLER_0_119_265 ();
 sg13g2_fill_1 FILLER_0_119_267 ();
 sg13g2_fill_2 FILLER_0_119_335 ();
 sg13g2_fill_8 FILLER_0_119_342 ();
 sg13g2_fill_2 FILLER_0_119_399 ();
 sg13g2_decap_8 FILLER_0_119_409 ();
 sg13g2_fill_2 FILLER_0_119_424 ();
 sg13g2_decap_8 FILLER_0_119_440 ();
 sg13g2_fill_8 FILLER_0_119_452 ();
 sg13g2_fill_1 FILLER_0_119_460 ();
 sg13g2_fill_1 FILLER_0_119_486 ();
 sg13g2_fill_8 FILLER_0_119_513 ();
 sg13g2_fill_2 FILLER_0_119_521 ();
 sg13g2_fill_4 FILLER_0_119_527 ();
 sg13g2_fill_4 FILLER_0_119_562 ();
 sg13g2_fill_4 FILLER_0_119_576 ();
 sg13g2_fill_1 FILLER_0_119_580 ();
 sg13g2_fill_1 FILLER_0_119_585 ();
 sg13g2_fill_2 FILLER_0_119_596 ();
 sg13g2_fill_1 FILLER_0_119_632 ();
 sg13g2_fill_1 FILLER_0_119_707 ();
 sg13g2_fill_8 FILLER_0_119_712 ();
 sg13g2_fill_2 FILLER_0_119_772 ();
 sg13g2_fill_1 FILLER_0_119_774 ();
 sg13g2_fill_1 FILLER_0_119_785 ();
 sg13g2_fill_4 FILLER_0_119_806 ();
 sg13g2_fill_1 FILLER_0_119_810 ();
 sg13g2_fill_8 FILLER_0_119_815 ();
 sg13g2_fill_4 FILLER_0_119_823 ();
 sg13g2_fill_2 FILLER_0_119_827 ();
 sg13g2_fill_2 FILLER_0_119_833 ();
 sg13g2_fill_1 FILLER_0_119_835 ();
 sg13g2_fill_2 FILLER_0_119_862 ();
 sg13g2_fill_4 FILLER_0_119_869 ();
 sg13g2_fill_1 FILLER_0_119_873 ();
 sg13g2_fill_4 FILLER_0_119_878 ();
 sg13g2_fill_2 FILLER_0_119_882 ();
 sg13g2_fill_2 FILLER_0_119_887 ();
 sg13g2_fill_1 FILLER_0_119_889 ();
 sg13g2_fill_2 FILLER_0_119_907 ();
 sg13g2_fill_4 FILLER_0_119_917 ();
 sg13g2_fill_1 FILLER_0_119_921 ();
 sg13g2_fill_1 FILLER_0_119_926 ();
 sg13g2_fill_8 FILLER_0_119_957 ();
 sg13g2_fill_2 FILLER_0_119_965 ();
 sg13g2_fill_8 FILLER_0_119_981 ();
 sg13g2_fill_2 FILLER_0_119_989 ();
 sg13g2_fill_1 FILLER_0_119_991 ();
 sg13g2_fill_1 FILLER_0_119_997 ();
 sg13g2_fill_1 FILLER_0_119_1007 ();
 sg13g2_fill_2 FILLER_0_119_1013 ();
 sg13g2_fill_2 FILLER_0_119_1020 ();
 sg13g2_fill_1 FILLER_0_119_1032 ();
 sg13g2_fill_8 FILLER_0_119_1042 ();
 sg13g2_fill_4 FILLER_0_119_1054 ();
 sg13g2_fill_8 FILLER_0_119_1065 ();
 sg13g2_fill_2 FILLER_0_119_1073 ();
 sg13g2_fill_1 FILLER_0_119_1075 ();
 sg13g2_fill_8 FILLER_0_119_1080 ();
 sg13g2_fill_8 FILLER_0_119_1088 ();
 sg13g2_fill_8 FILLER_0_119_1096 ();
 sg13g2_fill_8 FILLER_0_119_1104 ();
 sg13g2_fill_8 FILLER_0_119_1112 ();
 sg13g2_fill_2 FILLER_0_119_1120 ();
 sg13g2_fill_2 FILLER_0_119_1136 ();
 sg13g2_fill_4 FILLER_0_119_1151 ();
 sg13g2_fill_1 FILLER_0_119_1155 ();
 sg13g2_fill_1 FILLER_0_119_1169 ();
 sg13g2_fill_1 FILLER_0_119_1193 ();
 sg13g2_fill_1 FILLER_0_119_1199 ();
 sg13g2_fill_2 FILLER_0_119_1217 ();
 sg13g2_fill_2 FILLER_0_119_1225 ();
 sg13g2_fill_1 FILLER_0_119_1227 ();
 sg13g2_fill_8 FILLER_0_120_0 ();
 sg13g2_fill_8 FILLER_0_120_8 ();
 sg13g2_fill_8 FILLER_0_120_16 ();
 sg13g2_fill_8 FILLER_0_120_24 ();
 sg13g2_fill_8 FILLER_0_120_32 ();
 sg13g2_fill_8 FILLER_0_120_40 ();
 sg13g2_fill_8 FILLER_0_120_48 ();
 sg13g2_fill_8 FILLER_0_120_56 ();
 sg13g2_fill_8 FILLER_0_120_64 ();
 sg13g2_fill_8 FILLER_0_120_72 ();
 sg13g2_fill_8 FILLER_0_120_80 ();
 sg13g2_fill_8 FILLER_0_120_88 ();
 sg13g2_fill_8 FILLER_0_120_96 ();
 sg13g2_fill_8 FILLER_0_120_104 ();
 sg13g2_fill_8 FILLER_0_120_112 ();
 sg13g2_fill_4 FILLER_0_120_120 ();
 sg13g2_fill_2 FILLER_0_120_124 ();
 sg13g2_fill_1 FILLER_0_120_135 ();
 sg13g2_fill_8 FILLER_0_120_155 ();
 sg13g2_fill_2 FILLER_0_120_163 ();
 sg13g2_fill_8 FILLER_0_120_169 ();
 sg13g2_fill_2 FILLER_0_120_177 ();
 sg13g2_fill_1 FILLER_0_120_179 ();
 sg13g2_fill_4 FILLER_0_120_204 ();
 sg13g2_fill_2 FILLER_0_120_208 ();
 sg13g2_fill_2 FILLER_0_120_214 ();
 sg13g2_decap_8 FILLER_0_120_220 ();
 sg13g2_fill_2 FILLER_0_120_235 ();
 sg13g2_fill_1 FILLER_0_120_237 ();
 sg13g2_fill_2 FILLER_0_120_269 ();
 sg13g2_decap_8 FILLER_0_120_297 ();
 sg13g2_fill_2 FILLER_0_120_326 ();
 sg13g2_fill_1 FILLER_0_120_328 ();
 sg13g2_fill_8 FILLER_0_120_334 ();
 sg13g2_fill_8 FILLER_0_120_342 ();
 sg13g2_fill_8 FILLER_0_120_350 ();
 sg13g2_decap_8 FILLER_0_120_358 ();
 sg13g2_fill_1 FILLER_0_120_383 ();
 sg13g2_fill_1 FILLER_0_120_394 ();
 sg13g2_fill_8 FILLER_0_120_399 ();
 sg13g2_fill_2 FILLER_0_120_407 ();
 sg13g2_fill_1 FILLER_0_120_409 ();
 sg13g2_fill_4 FILLER_0_120_441 ();
 sg13g2_fill_1 FILLER_0_120_476 ();
 sg13g2_fill_8 FILLER_0_120_481 ();
 sg13g2_fill_8 FILLER_0_120_489 ();
 sg13g2_fill_8 FILLER_0_120_497 ();
 sg13g2_fill_8 FILLER_0_120_505 ();
 sg13g2_fill_4 FILLER_0_120_513 ();
 sg13g2_fill_1 FILLER_0_120_548 ();
 sg13g2_fill_2 FILLER_0_120_563 ();
 sg13g2_fill_4 FILLER_0_120_570 ();
 sg13g2_fill_4 FILLER_0_120_578 ();
 sg13g2_fill_2 FILLER_0_120_592 ();
 sg13g2_fill_2 FILLER_0_120_599 ();
 sg13g2_fill_1 FILLER_0_120_633 ();
 sg13g2_fill_8 FILLER_0_120_649 ();
 sg13g2_fill_4 FILLER_0_120_657 ();
 sg13g2_fill_4 FILLER_0_120_665 ();
 sg13g2_fill_2 FILLER_0_120_669 ();
 sg13g2_fill_8 FILLER_0_120_676 ();
 sg13g2_fill_1 FILLER_0_120_684 ();
 sg13g2_fill_8 FILLER_0_120_730 ();
 sg13g2_fill_4 FILLER_0_120_738 ();
 sg13g2_fill_2 FILLER_0_120_742 ();
 sg13g2_fill_1 FILLER_0_120_752 ();
 sg13g2_decap_8 FILLER_0_120_834 ();
 sg13g2_fill_2 FILLER_0_120_845 ();
 sg13g2_fill_2 FILLER_0_120_861 ();
 sg13g2_fill_1 FILLER_0_120_863 ();
 sg13g2_fill_1 FILLER_0_120_869 ();
 sg13g2_fill_1 FILLER_0_120_875 ();
 sg13g2_fill_1 FILLER_0_120_902 ();
 sg13g2_fill_1 FILLER_0_120_908 ();
 sg13g2_fill_2 FILLER_0_120_917 ();
 sg13g2_fill_2 FILLER_0_120_937 ();
 sg13g2_fill_1 FILLER_0_120_939 ();
 sg13g2_fill_2 FILLER_0_120_950 ();
 sg13g2_decap_8 FILLER_0_120_962 ();
 sg13g2_fill_2 FILLER_0_120_977 ();
 sg13g2_fill_4 FILLER_0_120_984 ();
 sg13g2_fill_1 FILLER_0_120_992 ();
 sg13g2_fill_4 FILLER_0_120_1011 ();
 sg13g2_fill_2 FILLER_0_120_1015 ();
 sg13g2_fill_1 FILLER_0_120_1027 ();
 sg13g2_fill_8 FILLER_0_120_1043 ();
 sg13g2_fill_2 FILLER_0_120_1051 ();
 sg13g2_fill_1 FILLER_0_120_1053 ();
 sg13g2_fill_8 FILLER_0_120_1058 ();
 sg13g2_decap_8 FILLER_0_120_1066 ();
 sg13g2_fill_4 FILLER_0_120_1078 ();
 sg13g2_fill_1 FILLER_0_120_1082 ();
 sg13g2_fill_2 FILLER_0_120_1098 ();
 sg13g2_fill_1 FILLER_0_120_1104 ();
 sg13g2_fill_1 FILLER_0_120_1109 ();
 sg13g2_fill_2 FILLER_0_120_1115 ();
 sg13g2_fill_1 FILLER_0_120_1117 ();
 sg13g2_fill_1 FILLER_0_120_1124 ();
 sg13g2_fill_2 FILLER_0_120_1130 ();
 sg13g2_fill_1 FILLER_0_120_1132 ();
 sg13g2_fill_4 FILLER_0_120_1161 ();
 sg13g2_fill_2 FILLER_0_120_1165 ();
 sg13g2_fill_1 FILLER_0_120_1172 ();
 sg13g2_fill_1 FILLER_0_120_1177 ();
 sg13g2_fill_4 FILLER_0_120_1214 ();
 sg13g2_fill_8 FILLER_0_121_0 ();
 sg13g2_fill_8 FILLER_0_121_8 ();
 sg13g2_fill_8 FILLER_0_121_16 ();
 sg13g2_fill_8 FILLER_0_121_24 ();
 sg13g2_fill_8 FILLER_0_121_32 ();
 sg13g2_fill_8 FILLER_0_121_40 ();
 sg13g2_fill_8 FILLER_0_121_48 ();
 sg13g2_fill_8 FILLER_0_121_56 ();
 sg13g2_fill_8 FILLER_0_121_64 ();
 sg13g2_fill_8 FILLER_0_121_72 ();
 sg13g2_fill_4 FILLER_0_121_80 ();
 sg13g2_fill_8 FILLER_0_121_89 ();
 sg13g2_fill_8 FILLER_0_121_97 ();
 sg13g2_fill_8 FILLER_0_121_105 ();
 sg13g2_fill_8 FILLER_0_121_113 ();
 sg13g2_fill_8 FILLER_0_121_121 ();
 sg13g2_fill_8 FILLER_0_121_129 ();
 sg13g2_fill_4 FILLER_0_121_137 ();
 sg13g2_fill_2 FILLER_0_121_141 ();
 sg13g2_decap_8 FILLER_0_121_153 ();
 sg13g2_fill_4 FILLER_0_121_170 ();
 sg13g2_fill_2 FILLER_0_121_174 ();
 sg13g2_fill_8 FILLER_0_121_186 ();
 sg13g2_fill_4 FILLER_0_121_194 ();
 sg13g2_fill_8 FILLER_0_121_229 ();
 sg13g2_fill_8 FILLER_0_121_237 ();
 sg13g2_fill_8 FILLER_0_121_249 ();
 sg13g2_fill_8 FILLER_0_121_257 ();
 sg13g2_fill_8 FILLER_0_121_265 ();
 sg13g2_fill_4 FILLER_0_121_273 ();
 sg13g2_fill_1 FILLER_0_121_277 ();
 sg13g2_fill_1 FILLER_0_121_318 ();
 sg13g2_fill_2 FILLER_0_121_327 ();
 sg13g2_fill_1 FILLER_0_121_329 ();
 sg13g2_fill_8 FILLER_0_121_335 ();
 sg13g2_fill_8 FILLER_0_121_343 ();
 sg13g2_fill_8 FILLER_0_121_361 ();
 sg13g2_fill_4 FILLER_0_121_369 ();
 sg13g2_fill_1 FILLER_0_121_383 ();
 sg13g2_fill_1 FILLER_0_121_410 ();
 sg13g2_fill_2 FILLER_0_121_437 ();
 sg13g2_fill_1 FILLER_0_121_439 ();
 sg13g2_fill_8 FILLER_0_121_480 ();
 sg13g2_fill_8 FILLER_0_121_488 ();
 sg13g2_fill_8 FILLER_0_121_496 ();
 sg13g2_fill_8 FILLER_0_121_504 ();
 sg13g2_fill_8 FILLER_0_121_512 ();
 sg13g2_fill_8 FILLER_0_121_520 ();
 sg13g2_fill_8 FILLER_0_121_528 ();
 sg13g2_fill_8 FILLER_0_121_536 ();
 sg13g2_fill_8 FILLER_0_121_548 ();
 sg13g2_fill_8 FILLER_0_121_556 ();
 sg13g2_fill_2 FILLER_0_121_564 ();
 sg13g2_decap_8 FILLER_0_121_592 ();
 sg13g2_fill_8 FILLER_0_121_603 ();
 sg13g2_fill_4 FILLER_0_121_611 ();
 sg13g2_fill_1 FILLER_0_121_615 ();
 sg13g2_fill_8 FILLER_0_121_656 ();
 sg13g2_fill_8 FILLER_0_121_664 ();
 sg13g2_fill_2 FILLER_0_121_672 ();
 sg13g2_fill_8 FILLER_0_121_697 ();
 sg13g2_fill_2 FILLER_0_121_705 ();
 sg13g2_fill_8 FILLER_0_121_711 ();
 sg13g2_fill_8 FILLER_0_121_719 ();
 sg13g2_decap_8 FILLER_0_121_727 ();
 sg13g2_fill_4 FILLER_0_121_753 ();
 sg13g2_fill_2 FILLER_0_121_792 ();
 sg13g2_fill_8 FILLER_0_121_804 ();
 sg13g2_fill_2 FILLER_0_121_812 ();
 sg13g2_fill_8 FILLER_0_121_818 ();
 sg13g2_fill_8 FILLER_0_121_826 ();
 sg13g2_fill_8 FILLER_0_121_834 ();
 sg13g2_fill_8 FILLER_0_121_842 ();
 sg13g2_fill_4 FILLER_0_121_850 ();
 sg13g2_fill_2 FILLER_0_121_859 ();
 sg13g2_fill_4 FILLER_0_121_870 ();
 sg13g2_fill_2 FILLER_0_121_878 ();
 sg13g2_fill_2 FILLER_0_121_906 ();
 sg13g2_fill_2 FILLER_0_121_947 ();
 sg13g2_fill_1 FILLER_0_121_954 ();
 sg13g2_fill_1 FILLER_0_121_965 ();
 sg13g2_fill_2 FILLER_0_121_992 ();
 sg13g2_fill_1 FILLER_0_121_999 ();
 sg13g2_fill_2 FILLER_0_121_1009 ();
 sg13g2_fill_1 FILLER_0_121_1011 ();
 sg13g2_fill_1 FILLER_0_121_1017 ();
 sg13g2_fill_2 FILLER_0_121_1045 ();
 sg13g2_fill_1 FILLER_0_121_1047 ();
 sg13g2_fill_4 FILLER_0_121_1084 ();
 sg13g2_fill_4 FILLER_0_121_1112 ();
 sg13g2_fill_8 FILLER_0_121_1122 ();
 sg13g2_fill_2 FILLER_0_121_1130 ();
 sg13g2_fill_1 FILLER_0_121_1132 ();
 sg13g2_fill_1 FILLER_0_121_1159 ();
 sg13g2_fill_4 FILLER_0_121_1165 ();
 sg13g2_fill_1 FILLER_0_121_1169 ();
 sg13g2_fill_2 FILLER_0_121_1190 ();
 sg13g2_fill_1 FILLER_0_121_1192 ();
 sg13g2_fill_8 FILLER_0_121_1215 ();
 sg13g2_fill_4 FILLER_0_121_1223 ();
 sg13g2_fill_1 FILLER_0_121_1227 ();
 sg13g2_fill_8 FILLER_0_122_0 ();
 sg13g2_fill_8 FILLER_0_122_8 ();
 sg13g2_fill_8 FILLER_0_122_16 ();
 sg13g2_fill_8 FILLER_0_122_24 ();
 sg13g2_fill_8 FILLER_0_122_32 ();
 sg13g2_fill_8 FILLER_0_122_40 ();
 sg13g2_fill_8 FILLER_0_122_48 ();
 sg13g2_fill_8 FILLER_0_122_56 ();
 sg13g2_fill_8 FILLER_0_122_64 ();
 sg13g2_fill_8 FILLER_0_122_72 ();
 sg13g2_fill_8 FILLER_0_122_80 ();
 sg13g2_fill_8 FILLER_0_122_88 ();
 sg13g2_fill_8 FILLER_0_122_96 ();
 sg13g2_fill_8 FILLER_0_122_104 ();
 sg13g2_fill_8 FILLER_0_122_112 ();
 sg13g2_fill_2 FILLER_0_122_120 ();
 sg13g2_fill_1 FILLER_0_122_122 ();
 sg13g2_fill_1 FILLER_0_122_154 ();
 sg13g2_fill_8 FILLER_0_122_236 ();
 sg13g2_fill_8 FILLER_0_122_244 ();
 sg13g2_fill_8 FILLER_0_122_252 ();
 sg13g2_fill_8 FILLER_0_122_260 ();
 sg13g2_fill_8 FILLER_0_122_268 ();
 sg13g2_fill_8 FILLER_0_122_276 ();
 sg13g2_fill_2 FILLER_0_122_293 ();
 sg13g2_fill_2 FILLER_0_122_326 ();
 sg13g2_fill_2 FILLER_0_122_358 ();
 sg13g2_fill_1 FILLER_0_122_380 ();
 sg13g2_fill_1 FILLER_0_122_391 ();
 sg13g2_fill_1 FILLER_0_122_397 ();
 sg13g2_fill_8 FILLER_0_122_402 ();
 sg13g2_fill_4 FILLER_0_122_410 ();
 sg13g2_fill_2 FILLER_0_122_414 ();
 sg13g2_fill_2 FILLER_0_122_420 ();
 sg13g2_fill_1 FILLER_0_122_426 ();
 sg13g2_fill_2 FILLER_0_122_435 ();
 sg13g2_fill_1 FILLER_0_122_437 ();
 sg13g2_fill_2 FILLER_0_122_443 ();
 sg13g2_fill_8 FILLER_0_122_476 ();
 sg13g2_fill_8 FILLER_0_122_484 ();
 sg13g2_fill_8 FILLER_0_122_492 ();
 sg13g2_fill_8 FILLER_0_122_500 ();
 sg13g2_fill_8 FILLER_0_122_508 ();
 sg13g2_fill_8 FILLER_0_122_516 ();
 sg13g2_fill_4 FILLER_0_122_524 ();
 sg13g2_fill_2 FILLER_0_122_528 ();
 sg13g2_fill_4 FILLER_0_122_556 ();
 sg13g2_fill_2 FILLER_0_122_560 ();
 sg13g2_fill_4 FILLER_0_122_598 ();
 sg13g2_fill_1 FILLER_0_122_602 ();
 sg13g2_fill_2 FILLER_0_122_608 ();
 sg13g2_fill_1 FILLER_0_122_610 ();
 sg13g2_fill_2 FILLER_0_122_662 ();
 sg13g2_fill_8 FILLER_0_122_668 ();
 sg13g2_fill_4 FILLER_0_122_720 ();
 sg13g2_fill_2 FILLER_0_122_724 ();
 sg13g2_fill_1 FILLER_0_122_760 ();
 sg13g2_fill_4 FILLER_0_122_769 ();
 sg13g2_fill_4 FILLER_0_122_781 ();
 sg13g2_fill_1 FILLER_0_122_785 ();
 sg13g2_fill_2 FILLER_0_122_790 ();
 sg13g2_fill_1 FILLER_0_122_792 ();
 sg13g2_fill_8 FILLER_0_122_819 ();
 sg13g2_fill_8 FILLER_0_122_827 ();
 sg13g2_fill_2 FILLER_0_122_835 ();
 sg13g2_fill_1 FILLER_0_122_837 ();
 sg13g2_fill_2 FILLER_0_122_880 ();
 sg13g2_fill_2 FILLER_0_122_887 ();
 sg13g2_fill_1 FILLER_0_122_889 ();
 sg13g2_fill_2 FILLER_0_122_894 ();
 sg13g2_fill_1 FILLER_0_122_896 ();
 sg13g2_fill_2 FILLER_0_122_902 ();
 sg13g2_fill_1 FILLER_0_122_904 ();
 sg13g2_fill_4 FILLER_0_122_915 ();
 sg13g2_fill_1 FILLER_0_122_919 ();
 sg13g2_fill_4 FILLER_0_122_928 ();
 sg13g2_fill_4 FILLER_0_122_939 ();
 sg13g2_fill_1 FILLER_0_122_966 ();
 sg13g2_fill_2 FILLER_0_122_972 ();
 sg13g2_fill_1 FILLER_0_122_974 ();
 sg13g2_fill_1 FILLER_0_122_980 ();
 sg13g2_fill_2 FILLER_0_122_1007 ();
 sg13g2_fill_1 FILLER_0_122_1009 ();
 sg13g2_fill_1 FILLER_0_122_1030 ();
 sg13g2_fill_2 FILLER_0_122_1035 ();
 sg13g2_fill_1 FILLER_0_122_1057 ();
 sg13g2_fill_8 FILLER_0_122_1070 ();
 sg13g2_fill_8 FILLER_0_122_1078 ();
 sg13g2_fill_8 FILLER_0_122_1086 ();
 sg13g2_fill_4 FILLER_0_122_1094 ();
 sg13g2_fill_2 FILLER_0_122_1098 ();
 sg13g2_fill_8 FILLER_0_122_1109 ();
 sg13g2_fill_1 FILLER_0_122_1117 ();
 sg13g2_fill_1 FILLER_0_122_1129 ();
 sg13g2_fill_1 FILLER_0_122_1135 ();
 sg13g2_fill_1 FILLER_0_122_1144 ();
 sg13g2_fill_8 FILLER_0_122_1150 ();
 sg13g2_fill_8 FILLER_0_122_1158 ();
 sg13g2_fill_8 FILLER_0_122_1166 ();
 sg13g2_fill_2 FILLER_0_122_1174 ();
 sg13g2_fill_8 FILLER_0_122_1214 ();
 sg13g2_fill_4 FILLER_0_122_1222 ();
 sg13g2_fill_2 FILLER_0_122_1226 ();
 sg13g2_fill_8 FILLER_0_123_0 ();
 sg13g2_fill_8 FILLER_0_123_8 ();
 sg13g2_fill_8 FILLER_0_123_16 ();
 sg13g2_fill_8 FILLER_0_123_24 ();
 sg13g2_fill_8 FILLER_0_123_32 ();
 sg13g2_fill_8 FILLER_0_123_40 ();
 sg13g2_fill_8 FILLER_0_123_48 ();
 sg13g2_fill_8 FILLER_0_123_56 ();
 sg13g2_fill_8 FILLER_0_123_64 ();
 sg13g2_fill_8 FILLER_0_123_72 ();
 sg13g2_fill_8 FILLER_0_123_80 ();
 sg13g2_fill_8 FILLER_0_123_88 ();
 sg13g2_fill_8 FILLER_0_123_96 ();
 sg13g2_fill_8 FILLER_0_123_104 ();
 sg13g2_fill_8 FILLER_0_123_112 ();
 sg13g2_fill_8 FILLER_0_123_120 ();
 sg13g2_fill_8 FILLER_0_123_132 ();
 sg13g2_fill_8 FILLER_0_123_140 ();
 sg13g2_fill_1 FILLER_0_123_148 ();
 sg13g2_fill_2 FILLER_0_123_184 ();
 sg13g2_fill_1 FILLER_0_123_186 ();
 sg13g2_fill_8 FILLER_0_123_205 ();
 sg13g2_fill_8 FILLER_0_123_213 ();
 sg13g2_fill_8 FILLER_0_123_221 ();
 sg13g2_fill_8 FILLER_0_123_229 ();
 sg13g2_fill_8 FILLER_0_123_237 ();
 sg13g2_fill_8 FILLER_0_123_245 ();
 sg13g2_fill_8 FILLER_0_123_253 ();
 sg13g2_fill_8 FILLER_0_123_261 ();
 sg13g2_fill_8 FILLER_0_123_269 ();
 sg13g2_fill_8 FILLER_0_123_277 ();
 sg13g2_fill_8 FILLER_0_123_285 ();
 sg13g2_fill_4 FILLER_0_123_293 ();
 sg13g2_fill_1 FILLER_0_123_297 ();
 sg13g2_fill_1 FILLER_0_123_307 ();
 sg13g2_fill_1 FILLER_0_123_334 ();
 sg13g2_fill_2 FILLER_0_123_376 ();
 sg13g2_fill_2 FILLER_0_123_404 ();
 sg13g2_fill_8 FILLER_0_123_414 ();
 sg13g2_fill_4 FILLER_0_123_448 ();
 sg13g2_fill_1 FILLER_0_123_452 ();
 sg13g2_fill_2 FILLER_0_123_462 ();
 sg13g2_fill_4 FILLER_0_123_474 ();
 sg13g2_fill_1 FILLER_0_123_504 ();
 sg13g2_fill_8 FILLER_0_123_510 ();
 sg13g2_fill_1 FILLER_0_123_518 ();
 sg13g2_fill_1 FILLER_0_123_528 ();
 sg13g2_fill_4 FILLER_0_123_534 ();
 sg13g2_fill_2 FILLER_0_123_538 ();
 sg13g2_fill_8 FILLER_0_123_545 ();
 sg13g2_fill_8 FILLER_0_123_553 ();
 sg13g2_fill_1 FILLER_0_123_561 ();
 sg13g2_fill_4 FILLER_0_123_576 ();
 sg13g2_fill_2 FILLER_0_123_580 ();
 sg13g2_fill_1 FILLER_0_123_592 ();
 sg13g2_fill_2 FILLER_0_123_603 ();
 sg13g2_fill_4 FILLER_0_123_675 ();
 sg13g2_fill_8 FILLER_0_123_710 ();
 sg13g2_fill_2 FILLER_0_123_718 ();
 sg13g2_fill_1 FILLER_0_123_720 ();
 sg13g2_fill_1 FILLER_0_123_730 ();
 sg13g2_fill_8 FILLER_0_123_745 ();
 sg13g2_fill_1 FILLER_0_123_758 ();
 sg13g2_fill_2 FILLER_0_123_764 ();
 sg13g2_fill_1 FILLER_0_123_766 ();
 sg13g2_fill_2 FILLER_0_123_771 ();
 sg13g2_fill_1 FILLER_0_123_773 ();
 sg13g2_fill_2 FILLER_0_123_784 ();
 sg13g2_fill_1 FILLER_0_123_791 ();
 sg13g2_fill_1 FILLER_0_123_802 ();
 sg13g2_decap_8 FILLER_0_123_829 ();
 sg13g2_fill_2 FILLER_0_123_862 ();
 sg13g2_fill_8 FILLER_0_123_869 ();
 sg13g2_fill_1 FILLER_0_123_877 ();
 sg13g2_fill_8 FILLER_0_123_883 ();
 sg13g2_decap_8 FILLER_0_123_891 ();
 sg13g2_fill_8 FILLER_0_123_903 ();
 sg13g2_fill_8 FILLER_0_123_931 ();
 sg13g2_fill_8 FILLER_0_123_939 ();
 sg13g2_fill_1 FILLER_0_123_962 ();
 sg13g2_fill_2 FILLER_0_123_968 ();
 sg13g2_fill_8 FILLER_0_123_979 ();
 sg13g2_fill_1 FILLER_0_123_987 ();
 sg13g2_fill_2 FILLER_0_123_1001 ();
 sg13g2_fill_1 FILLER_0_123_1021 ();
 sg13g2_fill_2 FILLER_0_123_1027 ();
 sg13g2_fill_1 FILLER_0_123_1034 ();
 sg13g2_fill_1 FILLER_0_123_1041 ();
 sg13g2_decap_8 FILLER_0_123_1047 ();
 sg13g2_fill_4 FILLER_0_123_1083 ();
 sg13g2_fill_2 FILLER_0_123_1092 ();
 sg13g2_fill_2 FILLER_0_123_1102 ();
 sg13g2_fill_8 FILLER_0_123_1114 ();
 sg13g2_fill_4 FILLER_0_123_1122 ();
 sg13g2_fill_1 FILLER_0_123_1143 ();
 sg13g2_fill_1 FILLER_0_123_1156 ();
 sg13g2_fill_8 FILLER_0_123_1172 ();
 sg13g2_fill_8 FILLER_0_123_1180 ();
 sg13g2_fill_8 FILLER_0_123_1188 ();
 sg13g2_fill_1 FILLER_0_123_1196 ();
 sg13g2_fill_8 FILLER_0_123_1204 ();
 sg13g2_fill_8 FILLER_0_123_1212 ();
 sg13g2_fill_8 FILLER_0_123_1220 ();
 sg13g2_fill_8 FILLER_0_124_0 ();
 sg13g2_fill_8 FILLER_0_124_8 ();
 sg13g2_fill_8 FILLER_0_124_16 ();
 sg13g2_fill_8 FILLER_0_124_24 ();
 sg13g2_fill_8 FILLER_0_124_32 ();
 sg13g2_fill_8 FILLER_0_124_40 ();
 sg13g2_fill_8 FILLER_0_124_48 ();
 sg13g2_fill_8 FILLER_0_124_56 ();
 sg13g2_fill_8 FILLER_0_124_64 ();
 sg13g2_fill_8 FILLER_0_124_72 ();
 sg13g2_fill_8 FILLER_0_124_80 ();
 sg13g2_fill_8 FILLER_0_124_88 ();
 sg13g2_fill_8 FILLER_0_124_96 ();
 sg13g2_fill_8 FILLER_0_124_104 ();
 sg13g2_fill_8 FILLER_0_124_112 ();
 sg13g2_fill_8 FILLER_0_124_120 ();
 sg13g2_fill_8 FILLER_0_124_128 ();
 sg13g2_fill_8 FILLER_0_124_136 ();
 sg13g2_fill_8 FILLER_0_124_144 ();
 sg13g2_fill_2 FILLER_0_124_152 ();
 sg13g2_fill_1 FILLER_0_124_154 ();
 sg13g2_fill_2 FILLER_0_124_186 ();
 sg13g2_fill_2 FILLER_0_124_203 ();
 sg13g2_fill_4 FILLER_0_124_210 ();
 sg13g2_fill_1 FILLER_0_124_240 ();
 sg13g2_fill_4 FILLER_0_124_272 ();
 sg13g2_fill_2 FILLER_0_124_276 ();
 sg13g2_fill_8 FILLER_0_124_288 ();
 sg13g2_fill_8 FILLER_0_124_296 ();
 sg13g2_fill_4 FILLER_0_124_304 ();
 sg13g2_fill_2 FILLER_0_124_308 ();
 sg13g2_fill_1 FILLER_0_124_334 ();
 sg13g2_fill_2 FILLER_0_124_383 ();
 sg13g2_fill_8 FILLER_0_124_389 ();
 sg13g2_fill_8 FILLER_0_124_397 ();
 sg13g2_fill_1 FILLER_0_124_405 ();
 sg13g2_fill_8 FILLER_0_124_433 ();
 sg13g2_fill_2 FILLER_0_124_441 ();
 sg13g2_fill_1 FILLER_0_124_443 ();
 sg13g2_fill_8 FILLER_0_124_457 ();
 sg13g2_fill_2 FILLER_0_124_465 ();
 sg13g2_fill_2 FILLER_0_124_482 ();
 sg13g2_fill_1 FILLER_0_124_484 ();
 sg13g2_fill_2 FILLER_0_124_619 ();
 sg13g2_fill_2 FILLER_0_124_631 ();
 sg13g2_fill_1 FILLER_0_124_633 ();
 sg13g2_fill_2 FILLER_0_124_657 ();
 sg13g2_fill_1 FILLER_0_124_659 ();
 sg13g2_fill_2 FILLER_0_124_672 ();
 sg13g2_fill_4 FILLER_0_124_689 ();
 sg13g2_fill_8 FILLER_0_124_697 ();
 sg13g2_fill_8 FILLER_0_124_705 ();
 sg13g2_fill_2 FILLER_0_124_713 ();
 sg13g2_fill_4 FILLER_0_124_745 ();
 sg13g2_fill_2 FILLER_0_124_757 ();
 sg13g2_fill_1 FILLER_0_124_759 ();
 sg13g2_fill_4 FILLER_0_124_786 ();
 sg13g2_fill_1 FILLER_0_124_790 ();
 sg13g2_fill_8 FILLER_0_124_806 ();
 sg13g2_fill_8 FILLER_0_124_818 ();
 sg13g2_fill_8 FILLER_0_124_826 ();
 sg13g2_fill_2 FILLER_0_124_834 ();
 sg13g2_fill_4 FILLER_0_124_852 ();
 sg13g2_fill_1 FILLER_0_124_856 ();
 sg13g2_fill_2 FILLER_0_124_862 ();
 sg13g2_fill_1 FILLER_0_124_864 ();
 sg13g2_fill_4 FILLER_0_124_874 ();
 sg13g2_fill_1 FILLER_0_124_878 ();
 sg13g2_fill_1 FILLER_0_124_891 ();
 sg13g2_fill_1 FILLER_0_124_907 ();
 sg13g2_fill_1 FILLER_0_124_918 ();
 sg13g2_fill_2 FILLER_0_124_927 ();
 sg13g2_fill_2 FILLER_0_124_934 ();
 sg13g2_fill_1 FILLER_0_124_936 ();
 sg13g2_fill_1 FILLER_0_124_947 ();
 sg13g2_decap_8 FILLER_0_124_973 ();
 sg13g2_decap_8 FILLER_0_124_985 ();
 sg13g2_fill_8 FILLER_0_124_997 ();
 sg13g2_fill_8 FILLER_0_124_1005 ();
 sg13g2_fill_8 FILLER_0_124_1013 ();
 sg13g2_fill_2 FILLER_0_124_1021 ();
 sg13g2_fill_1 FILLER_0_124_1023 ();
 sg13g2_fill_2 FILLER_0_124_1036 ();
 sg13g2_fill_1 FILLER_0_124_1042 ();
 sg13g2_fill_2 FILLER_0_124_1049 ();
 sg13g2_fill_1 FILLER_0_124_1063 ();
 sg13g2_fill_1 FILLER_0_124_1076 ();
 sg13g2_fill_8 FILLER_0_124_1109 ();
 sg13g2_fill_8 FILLER_0_124_1117 ();
 sg13g2_fill_2 FILLER_0_124_1125 ();
 sg13g2_fill_1 FILLER_0_124_1127 ();
 sg13g2_fill_1 FILLER_0_124_1134 ();
 sg13g2_fill_2 FILLER_0_124_1166 ();
 sg13g2_fill_1 FILLER_0_124_1171 ();
 sg13g2_fill_8 FILLER_0_124_1180 ();
 sg13g2_fill_8 FILLER_0_124_1188 ();
 sg13g2_fill_8 FILLER_0_124_1196 ();
 sg13g2_fill_8 FILLER_0_124_1204 ();
 sg13g2_fill_8 FILLER_0_124_1212 ();
 sg13g2_fill_8 FILLER_0_124_1220 ();
 sg13g2_fill_8 FILLER_0_125_0 ();
 sg13g2_fill_8 FILLER_0_125_8 ();
 sg13g2_fill_8 FILLER_0_125_16 ();
 sg13g2_fill_8 FILLER_0_125_24 ();
 sg13g2_fill_8 FILLER_0_125_32 ();
 sg13g2_fill_8 FILLER_0_125_40 ();
 sg13g2_fill_8 FILLER_0_125_48 ();
 sg13g2_fill_8 FILLER_0_125_56 ();
 sg13g2_fill_8 FILLER_0_125_64 ();
 sg13g2_fill_8 FILLER_0_125_72 ();
 sg13g2_fill_8 FILLER_0_125_80 ();
 sg13g2_fill_8 FILLER_0_125_88 ();
 sg13g2_fill_8 FILLER_0_125_96 ();
 sg13g2_fill_8 FILLER_0_125_104 ();
 sg13g2_fill_4 FILLER_0_125_112 ();
 sg13g2_fill_1 FILLER_0_125_116 ();
 sg13g2_fill_8 FILLER_0_125_122 ();
 sg13g2_fill_8 FILLER_0_125_130 ();
 sg13g2_fill_8 FILLER_0_125_138 ();
 sg13g2_fill_8 FILLER_0_125_146 ();
 sg13g2_fill_8 FILLER_0_125_154 ();
 sg13g2_fill_4 FILLER_0_125_162 ();
 sg13g2_fill_1 FILLER_0_125_166 ();
 sg13g2_fill_2 FILLER_0_125_185 ();
 sg13g2_fill_4 FILLER_0_125_213 ();
 sg13g2_fill_8 FILLER_0_125_221 ();
 sg13g2_fill_8 FILLER_0_125_229 ();
 sg13g2_fill_8 FILLER_0_125_237 ();
 sg13g2_fill_2 FILLER_0_125_245 ();
 sg13g2_fill_1 FILLER_0_125_247 ();
 sg13g2_fill_8 FILLER_0_125_252 ();
 sg13g2_fill_8 FILLER_0_125_260 ();
 sg13g2_fill_2 FILLER_0_125_268 ();
 sg13g2_fill_1 FILLER_0_125_270 ();
 sg13g2_fill_8 FILLER_0_125_276 ();
 sg13g2_fill_8 FILLER_0_125_284 ();
 sg13g2_fill_8 FILLER_0_125_292 ();
 sg13g2_fill_8 FILLER_0_125_300 ();
 sg13g2_fill_8 FILLER_0_125_308 ();
 sg13g2_fill_2 FILLER_0_125_316 ();
 sg13g2_fill_1 FILLER_0_125_318 ();
 sg13g2_fill_8 FILLER_0_125_323 ();
 sg13g2_fill_8 FILLER_0_125_331 ();
 sg13g2_fill_4 FILLER_0_125_339 ();
 sg13g2_fill_1 FILLER_0_125_371 ();
 sg13g2_fill_4 FILLER_0_125_398 ();
 sg13g2_fill_1 FILLER_0_125_402 ();
 sg13g2_fill_1 FILLER_0_125_429 ();
 sg13g2_fill_1 FILLER_0_125_456 ();
 sg13g2_fill_2 FILLER_0_125_483 ();
 sg13g2_fill_2 FILLER_0_125_489 ();
 sg13g2_fill_2 FILLER_0_125_495 ();
 sg13g2_fill_2 FILLER_0_125_507 ();
 sg13g2_fill_4 FILLER_0_125_548 ();
 sg13g2_fill_2 FILLER_0_125_552 ();
 sg13g2_fill_4 FILLER_0_125_564 ();
 sg13g2_fill_2 FILLER_0_125_568 ();
 sg13g2_fill_8 FILLER_0_125_582 ();
 sg13g2_fill_2 FILLER_0_125_590 ();
 sg13g2_fill_1 FILLER_0_125_596 ();
 sg13g2_fill_1 FILLER_0_125_602 ();
 sg13g2_fill_1 FILLER_0_125_613 ();
 sg13g2_fill_1 FILLER_0_125_640 ();
 sg13g2_fill_2 FILLER_0_125_646 ();
 sg13g2_fill_4 FILLER_0_125_658 ();
 sg13g2_fill_2 FILLER_0_125_662 ();
 sg13g2_fill_8 FILLER_0_125_690 ();
 sg13g2_fill_8 FILLER_0_125_698 ();
 sg13g2_fill_4 FILLER_0_125_706 ();
 sg13g2_fill_1 FILLER_0_125_710 ();
 sg13g2_fill_1 FILLER_0_125_751 ();
 sg13g2_fill_8 FILLER_0_125_790 ();
 sg13g2_decap_8 FILLER_0_125_829 ();
 sg13g2_fill_2 FILLER_0_125_869 ();
 sg13g2_fill_1 FILLER_0_125_871 ();
 sg13g2_fill_2 FILLER_0_125_932 ();
 sg13g2_fill_1 FILLER_0_125_934 ();
 sg13g2_fill_4 FILLER_0_125_960 ();
 sg13g2_fill_1 FILLER_0_125_964 ();
 sg13g2_fill_4 FILLER_0_125_981 ();
 sg13g2_fill_2 FILLER_0_125_1001 ();
 sg13g2_fill_1 FILLER_0_125_1003 ();
 sg13g2_fill_1 FILLER_0_125_1019 ();
 sg13g2_fill_2 FILLER_0_125_1033 ();
 sg13g2_fill_1 FILLER_0_125_1039 ();
 sg13g2_fill_2 FILLER_0_125_1044 ();
 sg13g2_fill_1 FILLER_0_125_1046 ();
 sg13g2_fill_4 FILLER_0_125_1107 ();
 sg13g2_fill_2 FILLER_0_125_1120 ();
 sg13g2_fill_8 FILLER_0_125_1126 ();
 sg13g2_fill_1 FILLER_0_125_1146 ();
 sg13g2_fill_2 FILLER_0_125_1159 ();
 sg13g2_fill_1 FILLER_0_125_1178 ();
 sg13g2_fill_8 FILLER_0_125_1184 ();
 sg13g2_fill_8 FILLER_0_125_1192 ();
 sg13g2_fill_8 FILLER_0_125_1200 ();
 sg13g2_fill_8 FILLER_0_125_1208 ();
 sg13g2_fill_8 FILLER_0_125_1216 ();
 sg13g2_fill_4 FILLER_0_125_1224 ();
 sg13g2_fill_8 FILLER_0_126_0 ();
 sg13g2_fill_8 FILLER_0_126_8 ();
 sg13g2_fill_8 FILLER_0_126_16 ();
 sg13g2_fill_8 FILLER_0_126_24 ();
 sg13g2_fill_8 FILLER_0_126_32 ();
 sg13g2_fill_8 FILLER_0_126_40 ();
 sg13g2_fill_8 FILLER_0_126_48 ();
 sg13g2_fill_8 FILLER_0_126_56 ();
 sg13g2_fill_8 FILLER_0_126_64 ();
 sg13g2_fill_8 FILLER_0_126_72 ();
 sg13g2_fill_8 FILLER_0_126_80 ();
 sg13g2_fill_8 FILLER_0_126_88 ();
 sg13g2_fill_8 FILLER_0_126_96 ();
 sg13g2_fill_8 FILLER_0_126_104 ();
 sg13g2_fill_8 FILLER_0_126_112 ();
 sg13g2_fill_8 FILLER_0_126_120 ();
 sg13g2_fill_8 FILLER_0_126_128 ();
 sg13g2_fill_8 FILLER_0_126_136 ();
 sg13g2_fill_8 FILLER_0_126_144 ();
 sg13g2_fill_8 FILLER_0_126_152 ();
 sg13g2_fill_8 FILLER_0_126_160 ();
 sg13g2_fill_8 FILLER_0_126_168 ();
 sg13g2_fill_8 FILLER_0_126_176 ();
 sg13g2_fill_8 FILLER_0_126_184 ();
 sg13g2_fill_2 FILLER_0_126_192 ();
 sg13g2_fill_8 FILLER_0_126_198 ();
 sg13g2_fill_8 FILLER_0_126_206 ();
 sg13g2_fill_8 FILLER_0_126_214 ();
 sg13g2_fill_8 FILLER_0_126_222 ();
 sg13g2_fill_8 FILLER_0_126_230 ();
 sg13g2_fill_8 FILLER_0_126_238 ();
 sg13g2_fill_8 FILLER_0_126_246 ();
 sg13g2_decap_8 FILLER_0_126_254 ();
 sg13g2_fill_4 FILLER_0_126_302 ();
 sg13g2_fill_1 FILLER_0_126_306 ();
 sg13g2_fill_1 FILLER_0_126_311 ();
 sg13g2_fill_8 FILLER_0_126_338 ();
 sg13g2_fill_1 FILLER_0_126_346 ();
 sg13g2_fill_8 FILLER_0_126_352 ();
 sg13g2_fill_8 FILLER_0_126_360 ();
 sg13g2_fill_8 FILLER_0_126_368 ();
 sg13g2_fill_8 FILLER_0_126_376 ();
 sg13g2_fill_8 FILLER_0_126_384 ();
 sg13g2_fill_4 FILLER_0_126_392 ();
 sg13g2_fill_2 FILLER_0_126_396 ();
 sg13g2_fill_1 FILLER_0_126_450 ();
 sg13g2_fill_8 FILLER_0_126_487 ();
 sg13g2_fill_4 FILLER_0_126_533 ();
 sg13g2_fill_2 FILLER_0_126_541 ();
 sg13g2_fill_8 FILLER_0_126_573 ();
 sg13g2_fill_8 FILLER_0_126_581 ();
 sg13g2_fill_8 FILLER_0_126_589 ();
 sg13g2_fill_8 FILLER_0_126_597 ();
 sg13g2_fill_8 FILLER_0_126_605 ();
 sg13g2_fill_4 FILLER_0_126_613 ();
 sg13g2_fill_1 FILLER_0_126_617 ();
 sg13g2_fill_2 FILLER_0_126_630 ();
 sg13g2_fill_1 FILLER_0_126_632 ();
 sg13g2_fill_1 FILLER_0_126_679 ();
 sg13g2_fill_8 FILLER_0_126_695 ();
 sg13g2_fill_8 FILLER_0_126_703 ();
 sg13g2_fill_2 FILLER_0_126_719 ();
 sg13g2_fill_1 FILLER_0_126_721 ();
 sg13g2_fill_4 FILLER_0_126_727 ();
 sg13g2_fill_8 FILLER_0_126_741 ();
 sg13g2_fill_8 FILLER_0_126_749 ();
 sg13g2_fill_1 FILLER_0_126_757 ();
 sg13g2_fill_8 FILLER_0_126_788 ();
 sg13g2_fill_2 FILLER_0_126_796 ();
 sg13g2_fill_1 FILLER_0_126_798 ();
 sg13g2_fill_8 FILLER_0_126_818 ();
 sg13g2_fill_8 FILLER_0_126_826 ();
 sg13g2_fill_8 FILLER_0_126_834 ();
 sg13g2_fill_1 FILLER_0_126_846 ();
 sg13g2_fill_1 FILLER_0_126_851 ();
 sg13g2_fill_4 FILLER_0_126_871 ();
 sg13g2_fill_2 FILLER_0_126_875 ();
 sg13g2_fill_1 FILLER_0_126_889 ();
 sg13g2_fill_1 FILLER_0_126_895 ();
 sg13g2_fill_2 FILLER_0_126_914 ();
 sg13g2_fill_1 FILLER_0_126_938 ();
 sg13g2_fill_1 FILLER_0_126_947 ();
 sg13g2_fill_1 FILLER_0_126_956 ();
 sg13g2_fill_1 FILLER_0_126_977 ();
 sg13g2_fill_2 FILLER_0_126_1002 ();
 sg13g2_fill_1 FILLER_0_126_1004 ();
 sg13g2_fill_1 FILLER_0_126_1010 ();
 sg13g2_fill_1 FILLER_0_126_1038 ();
 sg13g2_fill_1 FILLER_0_126_1084 ();
 sg13g2_fill_2 FILLER_0_126_1098 ();
 sg13g2_fill_1 FILLER_0_126_1100 ();
 sg13g2_fill_2 FILLER_0_126_1113 ();
 sg13g2_fill_1 FILLER_0_126_1119 ();
 sg13g2_fill_8 FILLER_0_126_1184 ();
 sg13g2_fill_8 FILLER_0_126_1192 ();
 sg13g2_fill_8 FILLER_0_126_1200 ();
 sg13g2_fill_8 FILLER_0_126_1208 ();
 sg13g2_fill_8 FILLER_0_126_1216 ();
 sg13g2_fill_4 FILLER_0_126_1224 ();
 sg13g2_fill_8 FILLER_0_127_0 ();
 sg13g2_fill_8 FILLER_0_127_8 ();
 sg13g2_fill_8 FILLER_0_127_16 ();
 sg13g2_fill_8 FILLER_0_127_24 ();
 sg13g2_fill_8 FILLER_0_127_32 ();
 sg13g2_fill_8 FILLER_0_127_40 ();
 sg13g2_fill_8 FILLER_0_127_48 ();
 sg13g2_fill_8 FILLER_0_127_56 ();
 sg13g2_fill_8 FILLER_0_127_64 ();
 sg13g2_fill_8 FILLER_0_127_72 ();
 sg13g2_fill_8 FILLER_0_127_80 ();
 sg13g2_fill_8 FILLER_0_127_88 ();
 sg13g2_fill_8 FILLER_0_127_96 ();
 sg13g2_fill_8 FILLER_0_127_104 ();
 sg13g2_fill_8 FILLER_0_127_112 ();
 sg13g2_fill_8 FILLER_0_127_120 ();
 sg13g2_fill_8 FILLER_0_127_128 ();
 sg13g2_fill_8 FILLER_0_127_136 ();
 sg13g2_fill_8 FILLER_0_127_144 ();
 sg13g2_fill_8 FILLER_0_127_152 ();
 sg13g2_fill_8 FILLER_0_127_160 ();
 sg13g2_fill_8 FILLER_0_127_168 ();
 sg13g2_fill_8 FILLER_0_127_176 ();
 sg13g2_fill_8 FILLER_0_127_184 ();
 sg13g2_fill_8 FILLER_0_127_192 ();
 sg13g2_fill_8 FILLER_0_127_200 ();
 sg13g2_fill_8 FILLER_0_127_208 ();
 sg13g2_fill_8 FILLER_0_127_216 ();
 sg13g2_fill_8 FILLER_0_127_224 ();
 sg13g2_fill_8 FILLER_0_127_232 ();
 sg13g2_fill_2 FILLER_0_127_240 ();
 sg13g2_fill_1 FILLER_0_127_242 ();
 sg13g2_fill_2 FILLER_0_127_303 ();
 sg13g2_fill_2 FILLER_0_127_331 ();
 sg13g2_fill_2 FILLER_0_127_337 ();
 sg13g2_fill_1 FILLER_0_127_339 ();
 sg13g2_fill_2 FILLER_0_127_371 ();
 sg13g2_fill_1 FILLER_0_127_373 ();
 sg13g2_fill_8 FILLER_0_127_393 ();
 sg13g2_fill_4 FILLER_0_127_401 ();
 sg13g2_fill_2 FILLER_0_127_405 ();
 sg13g2_fill_2 FILLER_0_127_436 ();
 sg13g2_fill_1 FILLER_0_127_442 ();
 sg13g2_fill_1 FILLER_0_127_453 ();
 sg13g2_fill_8 FILLER_0_127_482 ();
 sg13g2_fill_8 FILLER_0_127_490 ();
 sg13g2_fill_4 FILLER_0_127_498 ();
 sg13g2_fill_1 FILLER_0_127_502 ();
 sg13g2_fill_4 FILLER_0_127_523 ();
 sg13g2_fill_1 FILLER_0_127_527 ();
 sg13g2_fill_8 FILLER_0_127_533 ();
 sg13g2_fill_2 FILLER_0_127_541 ();
 sg13g2_fill_2 FILLER_0_127_548 ();
 sg13g2_fill_1 FILLER_0_127_550 ();
 sg13g2_fill_4 FILLER_0_127_561 ();
 sg13g2_fill_1 FILLER_0_127_565 ();
 sg13g2_fill_2 FILLER_0_127_592 ();
 sg13g2_fill_4 FILLER_0_127_604 ();
 sg13g2_fill_1 FILLER_0_127_608 ();
 sg13g2_fill_8 FILLER_0_127_613 ();
 sg13g2_fill_8 FILLER_0_127_621 ();
 sg13g2_fill_4 FILLER_0_127_629 ();
 sg13g2_fill_2 FILLER_0_127_664 ();
 sg13g2_fill_1 FILLER_0_127_666 ();
 sg13g2_fill_1 FILLER_0_127_672 ();
 sg13g2_fill_8 FILLER_0_127_703 ();
 sg13g2_fill_2 FILLER_0_127_711 ();
 sg13g2_fill_1 FILLER_0_127_713 ();
 sg13g2_fill_2 FILLER_0_127_719 ();
 sg13g2_fill_2 FILLER_0_127_731 ();
 sg13g2_fill_1 FILLER_0_127_733 ();
 sg13g2_decap_8 FILLER_0_127_753 ();
 sg13g2_fill_2 FILLER_0_127_790 ();
 sg13g2_fill_2 FILLER_0_127_797 ();
 sg13g2_fill_2 FILLER_0_127_809 ();
 sg13g2_fill_1 FILLER_0_127_811 ();
 sg13g2_fill_2 FILLER_0_127_838 ();
 sg13g2_fill_2 FILLER_0_127_875 ();
 sg13g2_fill_1 FILLER_0_127_877 ();
 sg13g2_fill_1 FILLER_0_127_906 ();
 sg13g2_fill_1 FILLER_0_127_966 ();
 sg13g2_fill_2 FILLER_0_127_975 ();
 sg13g2_decap_8 FILLER_0_127_987 ();
 sg13g2_fill_1 FILLER_0_127_1007 ();
 sg13g2_fill_1 FILLER_0_127_1012 ();
 sg13g2_fill_2 FILLER_0_127_1026 ();
 sg13g2_fill_1 FILLER_0_127_1043 ();
 sg13g2_fill_2 FILLER_0_127_1048 ();
 sg13g2_fill_2 FILLER_0_127_1069 ();
 sg13g2_fill_1 FILLER_0_127_1071 ();
 sg13g2_fill_2 FILLER_0_127_1118 ();
 sg13g2_fill_1 FILLER_0_127_1120 ();
 sg13g2_fill_2 FILLER_0_127_1128 ();
 sg13g2_fill_8 FILLER_0_127_1185 ();
 sg13g2_fill_8 FILLER_0_127_1193 ();
 sg13g2_fill_8 FILLER_0_127_1201 ();
 sg13g2_fill_8 FILLER_0_127_1209 ();
 sg13g2_fill_8 FILLER_0_127_1217 ();
 sg13g2_fill_2 FILLER_0_127_1225 ();
 sg13g2_fill_1 FILLER_0_127_1227 ();
 sg13g2_fill_8 FILLER_0_128_0 ();
 sg13g2_fill_8 FILLER_0_128_8 ();
 sg13g2_fill_8 FILLER_0_128_16 ();
 sg13g2_fill_8 FILLER_0_128_24 ();
 sg13g2_fill_8 FILLER_0_128_32 ();
 sg13g2_fill_8 FILLER_0_128_40 ();
 sg13g2_fill_8 FILLER_0_128_48 ();
 sg13g2_fill_8 FILLER_0_128_56 ();
 sg13g2_fill_8 FILLER_0_128_64 ();
 sg13g2_fill_8 FILLER_0_128_72 ();
 sg13g2_fill_8 FILLER_0_128_80 ();
 sg13g2_fill_8 FILLER_0_128_88 ();
 sg13g2_fill_8 FILLER_0_128_96 ();
 sg13g2_fill_8 FILLER_0_128_104 ();
 sg13g2_fill_8 FILLER_0_128_112 ();
 sg13g2_fill_8 FILLER_0_128_120 ();
 sg13g2_fill_8 FILLER_0_128_128 ();
 sg13g2_fill_8 FILLER_0_128_136 ();
 sg13g2_fill_8 FILLER_0_128_144 ();
 sg13g2_fill_8 FILLER_0_128_152 ();
 sg13g2_fill_8 FILLER_0_128_160 ();
 sg13g2_fill_8 FILLER_0_128_168 ();
 sg13g2_fill_8 FILLER_0_128_176 ();
 sg13g2_fill_8 FILLER_0_128_184 ();
 sg13g2_fill_8 FILLER_0_128_192 ();
 sg13g2_fill_8 FILLER_0_128_200 ();
 sg13g2_fill_8 FILLER_0_128_208 ();
 sg13g2_fill_8 FILLER_0_128_216 ();
 sg13g2_fill_8 FILLER_0_128_224 ();
 sg13g2_fill_8 FILLER_0_128_232 ();
 sg13g2_fill_2 FILLER_0_128_240 ();
 sg13g2_fill_4 FILLER_0_128_247 ();
 sg13g2_fill_2 FILLER_0_128_255 ();
 sg13g2_fill_2 FILLER_0_128_307 ();
 sg13g2_fill_8 FILLER_0_128_402 ();
 sg13g2_fill_4 FILLER_0_128_410 ();
 sg13g2_fill_2 FILLER_0_128_432 ();
 sg13g2_fill_2 FILLER_0_128_438 ();
 sg13g2_fill_8 FILLER_0_128_444 ();
 sg13g2_fill_8 FILLER_0_128_452 ();
 sg13g2_fill_8 FILLER_0_128_460 ();
 sg13g2_fill_8 FILLER_0_128_468 ();
 sg13g2_fill_8 FILLER_0_128_476 ();
 sg13g2_fill_4 FILLER_0_128_484 ();
 sg13g2_fill_2 FILLER_0_128_528 ();
 sg13g2_fill_4 FILLER_0_128_566 ();
 sg13g2_fill_1 FILLER_0_128_596 ();
 sg13g2_fill_1 FILLER_0_128_697 ();
 sg13g2_fill_2 FILLER_0_128_733 ();
 sg13g2_fill_1 FILLER_0_128_766 ();
 sg13g2_fill_1 FILLER_0_128_793 ();
 sg13g2_fill_8 FILLER_0_128_824 ();
 sg13g2_fill_4 FILLER_0_128_832 ();
 sg13g2_fill_2 FILLER_0_128_836 ();
 sg13g2_fill_8 FILLER_0_128_869 ();
 sg13g2_fill_8 FILLER_0_128_877 ();
 sg13g2_fill_2 FILLER_0_128_885 ();
 sg13g2_fill_4 FILLER_0_128_892 ();
 sg13g2_fill_1 FILLER_0_128_932 ();
 sg13g2_fill_4 FILLER_0_128_941 ();
 sg13g2_fill_2 FILLER_0_128_954 ();
 sg13g2_fill_1 FILLER_0_128_956 ();
 sg13g2_fill_8 FILLER_0_128_961 ();
 sg13g2_fill_4 FILLER_0_128_969 ();
 sg13g2_fill_2 FILLER_0_128_973 ();
 sg13g2_fill_8 FILLER_0_128_980 ();
 sg13g2_fill_8 FILLER_0_128_988 ();
 sg13g2_fill_2 FILLER_0_128_996 ();
 sg13g2_fill_4 FILLER_0_128_1007 ();
 sg13g2_fill_2 FILLER_0_128_1011 ();
 sg13g2_fill_4 FILLER_0_128_1017 ();
 sg13g2_fill_8 FILLER_0_128_1026 ();
 sg13g2_fill_2 FILLER_0_128_1034 ();
 sg13g2_fill_1 FILLER_0_128_1036 ();
 sg13g2_fill_1 FILLER_0_128_1041 ();
 sg13g2_fill_2 FILLER_0_128_1047 ();
 sg13g2_fill_4 FILLER_0_128_1057 ();
 sg13g2_fill_4 FILLER_0_128_1066 ();
 sg13g2_fill_1 FILLER_0_128_1070 ();
 sg13g2_fill_2 FILLER_0_128_1075 ();
 sg13g2_fill_2 FILLER_0_128_1086 ();
 sg13g2_fill_1 FILLER_0_128_1093 ();
 sg13g2_fill_1 FILLER_0_128_1098 ();
 sg13g2_fill_2 FILLER_0_128_1104 ();
 sg13g2_fill_2 FILLER_0_128_1120 ();
 sg13g2_fill_2 FILLER_0_128_1127 ();
 sg13g2_fill_2 FILLER_0_128_1133 ();
 sg13g2_fill_1 FILLER_0_128_1135 ();
 sg13g2_fill_1 FILLER_0_128_1141 ();
 sg13g2_fill_1 FILLER_0_128_1147 ();
 sg13g2_fill_1 FILLER_0_128_1163 ();
 sg13g2_fill_8 FILLER_0_128_1169 ();
 sg13g2_fill_8 FILLER_0_128_1177 ();
 sg13g2_fill_8 FILLER_0_128_1185 ();
 sg13g2_fill_8 FILLER_0_128_1193 ();
 sg13g2_fill_8 FILLER_0_128_1201 ();
 sg13g2_fill_8 FILLER_0_128_1209 ();
 sg13g2_fill_8 FILLER_0_128_1217 ();
 sg13g2_fill_2 FILLER_0_128_1225 ();
 sg13g2_fill_1 FILLER_0_128_1227 ();
 sg13g2_fill_8 FILLER_0_129_0 ();
 sg13g2_fill_8 FILLER_0_129_8 ();
 sg13g2_fill_8 FILLER_0_129_16 ();
 sg13g2_fill_8 FILLER_0_129_24 ();
 sg13g2_fill_8 FILLER_0_129_32 ();
 sg13g2_fill_8 FILLER_0_129_40 ();
 sg13g2_fill_8 FILLER_0_129_48 ();
 sg13g2_fill_8 FILLER_0_129_56 ();
 sg13g2_fill_8 FILLER_0_129_64 ();
 sg13g2_fill_8 FILLER_0_129_72 ();
 sg13g2_fill_8 FILLER_0_129_80 ();
 sg13g2_fill_8 FILLER_0_129_88 ();
 sg13g2_fill_8 FILLER_0_129_96 ();
 sg13g2_fill_8 FILLER_0_129_104 ();
 sg13g2_fill_8 FILLER_0_129_112 ();
 sg13g2_fill_8 FILLER_0_129_120 ();
 sg13g2_fill_8 FILLER_0_129_128 ();
 sg13g2_fill_8 FILLER_0_129_136 ();
 sg13g2_fill_8 FILLER_0_129_144 ();
 sg13g2_fill_8 FILLER_0_129_152 ();
 sg13g2_fill_8 FILLER_0_129_160 ();
 sg13g2_fill_8 FILLER_0_129_168 ();
 sg13g2_fill_8 FILLER_0_129_176 ();
 sg13g2_fill_8 FILLER_0_129_184 ();
 sg13g2_fill_8 FILLER_0_129_192 ();
 sg13g2_fill_8 FILLER_0_129_200 ();
 sg13g2_fill_8 FILLER_0_129_208 ();
 sg13g2_fill_8 FILLER_0_129_216 ();
 sg13g2_fill_8 FILLER_0_129_224 ();
 sg13g2_fill_4 FILLER_0_129_232 ();
 sg13g2_fill_1 FILLER_0_129_277 ();
 sg13g2_fill_2 FILLER_0_129_282 ();
 sg13g2_fill_2 FILLER_0_129_303 ();
 sg13g2_fill_1 FILLER_0_129_305 ();
 sg13g2_fill_2 FILLER_0_129_322 ();
 sg13g2_fill_2 FILLER_0_129_329 ();
 sg13g2_fill_1 FILLER_0_129_341 ();
 sg13g2_fill_2 FILLER_0_129_370 ();
 sg13g2_fill_1 FILLER_0_129_382 ();
 sg13g2_fill_4 FILLER_0_129_409 ();
 sg13g2_fill_1 FILLER_0_129_413 ();
 sg13g2_fill_4 FILLER_0_129_449 ();
 sg13g2_fill_1 FILLER_0_129_453 ();
 sg13g2_fill_2 FILLER_0_129_485 ();
 sg13g2_fill_8 FILLER_0_129_517 ();
 sg13g2_fill_2 FILLER_0_129_525 ();
 sg13g2_fill_2 FILLER_0_129_535 ();
 sg13g2_fill_4 FILLER_0_129_563 ();
 sg13g2_fill_1 FILLER_0_129_567 ();
 sg13g2_fill_1 FILLER_0_129_572 ();
 sg13g2_fill_1 FILLER_0_129_592 ();
 sg13g2_fill_1 FILLER_0_129_608 ();
 sg13g2_fill_8 FILLER_0_129_635 ();
 sg13g2_fill_8 FILLER_0_129_643 ();
 sg13g2_fill_2 FILLER_0_129_651 ();
 sg13g2_fill_1 FILLER_0_129_653 ();
 sg13g2_fill_8 FILLER_0_129_658 ();
 sg13g2_fill_8 FILLER_0_129_666 ();
 sg13g2_fill_2 FILLER_0_129_674 ();
 sg13g2_fill_8 FILLER_0_129_680 ();
 sg13g2_fill_8 FILLER_0_129_688 ();
 sg13g2_fill_2 FILLER_0_129_736 ();
 sg13g2_fill_1 FILLER_0_129_738 ();
 sg13g2_fill_4 FILLER_0_129_769 ();
 sg13g2_fill_8 FILLER_0_129_792 ();
 sg13g2_fill_1 FILLER_0_129_800 ();
 sg13g2_fill_2 FILLER_0_129_805 ();
 sg13g2_decap_8 FILLER_0_129_815 ();
 sg13g2_fill_8 FILLER_0_129_826 ();
 sg13g2_fill_8 FILLER_0_129_834 ();
 sg13g2_fill_2 FILLER_0_129_842 ();
 sg13g2_fill_1 FILLER_0_129_844 ();
 sg13g2_fill_2 FILLER_0_129_854 ();
 sg13g2_fill_2 FILLER_0_129_866 ();
 sg13g2_fill_1 FILLER_0_129_868 ();
 sg13g2_fill_1 FILLER_0_129_949 ();
 sg13g2_fill_4 FILLER_0_129_960 ();
 sg13g2_fill_8 FILLER_0_129_969 ();
 sg13g2_fill_8 FILLER_0_129_977 ();
 sg13g2_fill_2 FILLER_0_129_985 ();
 sg13g2_fill_1 FILLER_0_129_1003 ();
 sg13g2_fill_2 FILLER_0_129_1019 ();
 sg13g2_fill_1 FILLER_0_129_1074 ();
 sg13g2_fill_1 FILLER_0_129_1080 ();
 sg13g2_fill_1 FILLER_0_129_1085 ();
 sg13g2_fill_2 FILLER_0_129_1092 ();
 sg13g2_fill_2 FILLER_0_129_1108 ();
 sg13g2_fill_1 FILLER_0_129_1110 ();
 sg13g2_fill_2 FILLER_0_129_1115 ();
 sg13g2_fill_8 FILLER_0_129_1122 ();
 sg13g2_fill_8 FILLER_0_129_1130 ();
 sg13g2_fill_8 FILLER_0_129_1138 ();
 sg13g2_fill_4 FILLER_0_129_1146 ();
 sg13g2_fill_1 FILLER_0_129_1150 ();
 sg13g2_fill_8 FILLER_0_129_1163 ();
 sg13g2_fill_8 FILLER_0_129_1171 ();
 sg13g2_fill_8 FILLER_0_129_1179 ();
 sg13g2_fill_8 FILLER_0_129_1187 ();
 sg13g2_fill_8 FILLER_0_129_1195 ();
 sg13g2_fill_8 FILLER_0_129_1203 ();
 sg13g2_fill_8 FILLER_0_129_1211 ();
 sg13g2_fill_8 FILLER_0_129_1219 ();
 sg13g2_fill_1 FILLER_0_129_1227 ();
 sg13g2_fill_8 FILLER_0_130_0 ();
 sg13g2_fill_8 FILLER_0_130_8 ();
 sg13g2_fill_8 FILLER_0_130_16 ();
 sg13g2_fill_8 FILLER_0_130_24 ();
 sg13g2_fill_8 FILLER_0_130_32 ();
 sg13g2_fill_8 FILLER_0_130_40 ();
 sg13g2_fill_8 FILLER_0_130_48 ();
 sg13g2_fill_8 FILLER_0_130_56 ();
 sg13g2_fill_8 FILLER_0_130_64 ();
 sg13g2_fill_8 FILLER_0_130_72 ();
 sg13g2_fill_8 FILLER_0_130_80 ();
 sg13g2_fill_8 FILLER_0_130_88 ();
 sg13g2_fill_8 FILLER_0_130_96 ();
 sg13g2_fill_8 FILLER_0_130_104 ();
 sg13g2_fill_8 FILLER_0_130_112 ();
 sg13g2_fill_8 FILLER_0_130_120 ();
 sg13g2_fill_8 FILLER_0_130_128 ();
 sg13g2_fill_8 FILLER_0_130_136 ();
 sg13g2_fill_8 FILLER_0_130_144 ();
 sg13g2_fill_8 FILLER_0_130_152 ();
 sg13g2_fill_8 FILLER_0_130_160 ();
 sg13g2_fill_8 FILLER_0_130_168 ();
 sg13g2_fill_8 FILLER_0_130_176 ();
 sg13g2_fill_8 FILLER_0_130_184 ();
 sg13g2_fill_8 FILLER_0_130_192 ();
 sg13g2_fill_8 FILLER_0_130_200 ();
 sg13g2_fill_8 FILLER_0_130_208 ();
 sg13g2_fill_8 FILLER_0_130_216 ();
 sg13g2_fill_8 FILLER_0_130_224 ();
 sg13g2_fill_8 FILLER_0_130_232 ();
 sg13g2_fill_8 FILLER_0_130_240 ();
 sg13g2_fill_1 FILLER_0_130_248 ();
 sg13g2_fill_8 FILLER_0_130_253 ();
 sg13g2_fill_8 FILLER_0_130_261 ();
 sg13g2_fill_8 FILLER_0_130_269 ();
 sg13g2_fill_2 FILLER_0_130_277 ();
 sg13g2_fill_1 FILLER_0_130_305 ();
 sg13g2_fill_8 FILLER_0_130_329 ();
 sg13g2_fill_2 FILLER_0_130_337 ();
 sg13g2_fill_8 FILLER_0_130_347 ();
 sg13g2_fill_4 FILLER_0_130_355 ();
 sg13g2_fill_1 FILLER_0_130_359 ();
 sg13g2_fill_4 FILLER_0_130_364 ();
 sg13g2_fill_1 FILLER_0_130_387 ();
 sg13g2_fill_1 FILLER_0_130_393 ();
 sg13g2_fill_2 FILLER_0_130_398 ();
 sg13g2_fill_8 FILLER_0_130_466 ();
 sg13g2_fill_8 FILLER_0_130_474 ();
 sg13g2_fill_8 FILLER_0_130_518 ();
 sg13g2_fill_8 FILLER_0_130_526 ();
 sg13g2_decap_8 FILLER_0_130_534 ();
 sg13g2_fill_4 FILLER_0_130_546 ();
 sg13g2_fill_2 FILLER_0_130_550 ();
 sg13g2_fill_4 FILLER_0_130_562 ();
 sg13g2_fill_2 FILLER_0_130_566 ();
 sg13g2_fill_1 FILLER_0_130_598 ();
 sg13g2_fill_8 FILLER_0_130_629 ();
 sg13g2_fill_8 FILLER_0_130_637 ();
 sg13g2_decap_8 FILLER_0_130_645 ();
 sg13g2_fill_8 FILLER_0_130_662 ();
 sg13g2_fill_8 FILLER_0_130_670 ();
 sg13g2_fill_8 FILLER_0_130_678 ();
 sg13g2_fill_8 FILLER_0_130_686 ();
 sg13g2_decap_8 FILLER_0_130_694 ();
 sg13g2_fill_8 FILLER_0_130_745 ();
 sg13g2_fill_8 FILLER_0_130_753 ();
 sg13g2_fill_8 FILLER_0_130_761 ();
 sg13g2_fill_8 FILLER_0_130_769 ();
 sg13g2_fill_8 FILLER_0_130_777 ();
 sg13g2_fill_8 FILLER_0_130_785 ();
 sg13g2_fill_8 FILLER_0_130_793 ();
 sg13g2_fill_4 FILLER_0_130_801 ();
 sg13g2_fill_8 FILLER_0_130_841 ();
 sg13g2_fill_8 FILLER_0_130_849 ();
 sg13g2_fill_1 FILLER_0_130_857 ();
 sg13g2_fill_4 FILLER_0_130_871 ();
 sg13g2_fill_2 FILLER_0_130_879 ();
 sg13g2_fill_4 FILLER_0_130_901 ();
 sg13g2_fill_1 FILLER_0_130_905 ();
 sg13g2_fill_8 FILLER_0_130_910 ();
 sg13g2_fill_8 FILLER_0_130_918 ();
 sg13g2_fill_2 FILLER_0_130_926 ();
 sg13g2_fill_2 FILLER_0_130_940 ();
 sg13g2_fill_2 FILLER_0_130_951 ();
 sg13g2_fill_2 FILLER_0_130_973 ();
 sg13g2_fill_1 FILLER_0_130_1008 ();
 sg13g2_fill_2 FILLER_0_130_1013 ();
 sg13g2_fill_1 FILLER_0_130_1019 ();
 sg13g2_fill_1 FILLER_0_130_1024 ();
 sg13g2_fill_1 FILLER_0_130_1034 ();
 sg13g2_fill_1 FILLER_0_130_1039 ();
 sg13g2_fill_4 FILLER_0_130_1044 ();
 sg13g2_fill_2 FILLER_0_130_1052 ();
 sg13g2_fill_8 FILLER_0_130_1107 ();
 sg13g2_fill_8 FILLER_0_130_1115 ();
 sg13g2_fill_8 FILLER_0_130_1123 ();
 sg13g2_fill_8 FILLER_0_130_1131 ();
 sg13g2_fill_8 FILLER_0_130_1139 ();
 sg13g2_fill_8 FILLER_0_130_1147 ();
 sg13g2_fill_8 FILLER_0_130_1155 ();
 sg13g2_fill_8 FILLER_0_130_1163 ();
 sg13g2_fill_8 FILLER_0_130_1171 ();
 sg13g2_fill_8 FILLER_0_130_1179 ();
 sg13g2_fill_8 FILLER_0_130_1187 ();
 sg13g2_fill_8 FILLER_0_130_1195 ();
 sg13g2_fill_8 FILLER_0_130_1203 ();
 sg13g2_fill_8 FILLER_0_130_1211 ();
 sg13g2_fill_8 FILLER_0_130_1219 ();
 sg13g2_fill_1 FILLER_0_130_1227 ();
 sg13g2_fill_8 FILLER_0_131_0 ();
 sg13g2_fill_8 FILLER_0_131_8 ();
 sg13g2_fill_8 FILLER_0_131_16 ();
 sg13g2_fill_8 FILLER_0_131_24 ();
 sg13g2_fill_8 FILLER_0_131_32 ();
 sg13g2_fill_8 FILLER_0_131_40 ();
 sg13g2_fill_8 FILLER_0_131_48 ();
 sg13g2_fill_8 FILLER_0_131_56 ();
 sg13g2_fill_8 FILLER_0_131_64 ();
 sg13g2_fill_8 FILLER_0_131_72 ();
 sg13g2_fill_2 FILLER_0_131_80 ();
 sg13g2_fill_8 FILLER_0_131_116 ();
 sg13g2_fill_8 FILLER_0_131_124 ();
 sg13g2_fill_8 FILLER_0_131_132 ();
 sg13g2_fill_8 FILLER_0_131_140 ();
 sg13g2_fill_8 FILLER_0_131_148 ();
 sg13g2_fill_8 FILLER_0_131_156 ();
 sg13g2_fill_8 FILLER_0_131_164 ();
 sg13g2_fill_8 FILLER_0_131_172 ();
 sg13g2_fill_8 FILLER_0_131_180 ();
 sg13g2_fill_8 FILLER_0_131_188 ();
 sg13g2_fill_8 FILLER_0_131_196 ();
 sg13g2_fill_8 FILLER_0_131_204 ();
 sg13g2_fill_8 FILLER_0_131_212 ();
 sg13g2_fill_8 FILLER_0_131_220 ();
 sg13g2_fill_8 FILLER_0_131_228 ();
 sg13g2_fill_4 FILLER_0_131_236 ();
 sg13g2_fill_2 FILLER_0_131_240 ();
 sg13g2_decap_8 FILLER_0_131_272 ();
 sg13g2_fill_8 FILLER_0_131_320 ();
 sg13g2_fill_2 FILLER_0_131_328 ();
 sg13g2_fill_1 FILLER_0_131_330 ();
 sg13g2_fill_4 FILLER_0_131_336 ();
 sg13g2_fill_1 FILLER_0_131_340 ();
 sg13g2_fill_8 FILLER_0_131_346 ();
 sg13g2_fill_8 FILLER_0_131_354 ();
 sg13g2_fill_2 FILLER_0_131_362 ();
 sg13g2_fill_1 FILLER_0_131_364 ();
 sg13g2_fill_2 FILLER_0_131_396 ();
 sg13g2_fill_1 FILLER_0_131_398 ();
 sg13g2_fill_8 FILLER_0_131_407 ();
 sg13g2_decap_8 FILLER_0_131_415 ();
 sg13g2_fill_2 FILLER_0_131_447 ();
 sg13g2_fill_2 FILLER_0_131_485 ();
 sg13g2_fill_1 FILLER_0_131_487 ();
 sg13g2_fill_1 FILLER_0_131_512 ();
 sg13g2_fill_8 FILLER_0_131_518 ();
 sg13g2_fill_4 FILLER_0_131_526 ();
 sg13g2_fill_4 FILLER_0_131_538 ();
 sg13g2_fill_2 FILLER_0_131_546 ();
 sg13g2_fill_4 FILLER_0_131_563 ();
 sg13g2_fill_1 FILLER_0_131_567 ();
 sg13g2_fill_1 FILLER_0_131_607 ();
 sg13g2_fill_8 FILLER_0_131_618 ();
 sg13g2_fill_8 FILLER_0_131_626 ();
 sg13g2_fill_2 FILLER_0_131_664 ();
 sg13g2_fill_1 FILLER_0_131_666 ();
 sg13g2_fill_8 FILLER_0_131_698 ();
 sg13g2_fill_1 FILLER_0_131_706 ();
 sg13g2_fill_2 FILLER_0_131_716 ();
 sg13g2_fill_1 FILLER_0_131_718 ();
 sg13g2_fill_4 FILLER_0_131_760 ();
 sg13g2_fill_1 FILLER_0_131_774 ();
 sg13g2_fill_8 FILLER_0_131_779 ();
 sg13g2_fill_8 FILLER_0_131_787 ();
 sg13g2_fill_1 FILLER_0_131_795 ();
 sg13g2_fill_2 FILLER_0_131_822 ();
 sg13g2_decap_8 FILLER_0_131_854 ();
 sg13g2_fill_4 FILLER_0_131_900 ();
 sg13g2_fill_1 FILLER_0_131_916 ();
 sg13g2_fill_4 FILLER_0_131_922 ();
 sg13g2_fill_1 FILLER_0_131_951 ();
 sg13g2_fill_2 FILLER_0_131_978 ();
 sg13g2_fill_1 FILLER_0_131_984 ();
 sg13g2_fill_2 FILLER_0_131_989 ();
 sg13g2_fill_1 FILLER_0_131_991 ();
 sg13g2_fill_2 FILLER_0_131_997 ();
 sg13g2_fill_1 FILLER_0_131_999 ();
 sg13g2_fill_1 FILLER_0_131_1005 ();
 sg13g2_fill_2 FILLER_0_131_1011 ();
 sg13g2_fill_1 FILLER_0_131_1013 ();
 sg13g2_fill_1 FILLER_0_131_1059 ();
 sg13g2_fill_2 FILLER_0_131_1065 ();
 sg13g2_fill_1 FILLER_0_131_1067 ();
 sg13g2_fill_1 FILLER_0_131_1071 ();
 sg13g2_fill_1 FILLER_0_131_1076 ();
 sg13g2_fill_1 FILLER_0_131_1082 ();
 sg13g2_fill_2 FILLER_0_131_1087 ();
 sg13g2_fill_4 FILLER_0_131_1099 ();
 sg13g2_fill_1 FILLER_0_131_1103 ();
 sg13g2_fill_8 FILLER_0_131_1111 ();
 sg13g2_fill_8 FILLER_0_131_1119 ();
 sg13g2_fill_8 FILLER_0_131_1127 ();
 sg13g2_fill_8 FILLER_0_131_1135 ();
 sg13g2_fill_8 FILLER_0_131_1143 ();
 sg13g2_fill_8 FILLER_0_131_1151 ();
 sg13g2_fill_8 FILLER_0_131_1159 ();
 sg13g2_fill_8 FILLER_0_131_1167 ();
 sg13g2_fill_8 FILLER_0_131_1175 ();
 sg13g2_fill_8 FILLER_0_131_1183 ();
 sg13g2_fill_8 FILLER_0_131_1191 ();
 sg13g2_fill_8 FILLER_0_131_1199 ();
 sg13g2_fill_8 FILLER_0_131_1207 ();
 sg13g2_fill_8 FILLER_0_131_1215 ();
 sg13g2_fill_4 FILLER_0_131_1223 ();
 sg13g2_fill_1 FILLER_0_131_1227 ();
 sg13g2_fill_8 FILLER_0_132_0 ();
 sg13g2_fill_8 FILLER_0_132_8 ();
 sg13g2_fill_8 FILLER_0_132_16 ();
 sg13g2_fill_8 FILLER_0_132_24 ();
 sg13g2_fill_8 FILLER_0_132_32 ();
 sg13g2_fill_8 FILLER_0_132_40 ();
 sg13g2_fill_8 FILLER_0_132_48 ();
 sg13g2_fill_8 FILLER_0_132_56 ();
 sg13g2_fill_4 FILLER_0_132_64 ();
 sg13g2_fill_8 FILLER_0_132_146 ();
 sg13g2_fill_8 FILLER_0_132_154 ();
 sg13g2_fill_8 FILLER_0_132_162 ();
 sg13g2_fill_8 FILLER_0_132_170 ();
 sg13g2_fill_8 FILLER_0_132_178 ();
 sg13g2_fill_8 FILLER_0_132_186 ();
 sg13g2_fill_8 FILLER_0_132_194 ();
 sg13g2_fill_8 FILLER_0_132_202 ();
 sg13g2_fill_8 FILLER_0_132_210 ();
 sg13g2_fill_8 FILLER_0_132_218 ();
 sg13g2_fill_8 FILLER_0_132_226 ();
 sg13g2_fill_8 FILLER_0_132_234 ();
 sg13g2_fill_4 FILLER_0_132_242 ();
 sg13g2_fill_8 FILLER_0_132_275 ();
 sg13g2_fill_1 FILLER_0_132_327 ();
 sg13g2_fill_1 FILLER_0_132_364 ();
 sg13g2_fill_2 FILLER_0_132_391 ();
 sg13g2_fill_1 FILLER_0_132_419 ();
 sg13g2_fill_2 FILLER_0_132_425 ();
 sg13g2_fill_2 FILLER_0_132_431 ();
 sg13g2_fill_1 FILLER_0_132_433 ();
 sg13g2_fill_2 FILLER_0_132_438 ();
 sg13g2_fill_1 FILLER_0_132_440 ();
 sg13g2_fill_2 FILLER_0_132_464 ();
 sg13g2_fill_1 FILLER_0_132_466 ();
 sg13g2_fill_8 FILLER_0_132_475 ();
 sg13g2_fill_8 FILLER_0_132_483 ();
 sg13g2_fill_1 FILLER_0_132_491 ();
 sg13g2_fill_1 FILLER_0_132_496 ();
 sg13g2_fill_1 FILLER_0_132_523 ();
 sg13g2_fill_2 FILLER_0_132_528 ();
 sg13g2_fill_2 FILLER_0_132_534 ();
 sg13g2_fill_1 FILLER_0_132_536 ();
 sg13g2_fill_1 FILLER_0_132_541 ();
 sg13g2_decap_8 FILLER_0_132_568 ();
 sg13g2_fill_4 FILLER_0_132_579 ();
 sg13g2_fill_2 FILLER_0_132_583 ();
 sg13g2_fill_1 FILLER_0_132_593 ();
 sg13g2_fill_1 FILLER_0_132_598 ();
 sg13g2_fill_1 FILLER_0_132_618 ();
 sg13g2_fill_1 FILLER_0_132_623 ();
 sg13g2_decap_8 FILLER_0_132_650 ();
 sg13g2_fill_8 FILLER_0_132_698 ();
 sg13g2_fill_8 FILLER_0_132_706 ();
 sg13g2_fill_2 FILLER_0_132_714 ();
 sg13g2_fill_1 FILLER_0_132_757 ();
 sg13g2_fill_1 FILLER_0_132_763 ();
 sg13g2_fill_1 FILLER_0_132_816 ();
 sg13g2_fill_1 FILLER_0_132_827 ();
 sg13g2_fill_1 FILLER_0_132_842 ();
 sg13g2_fill_8 FILLER_0_132_861 ();
 sg13g2_fill_8 FILLER_0_132_869 ();
 sg13g2_fill_8 FILLER_0_132_877 ();
 sg13g2_fill_2 FILLER_0_132_885 ();
 sg13g2_decap_8 FILLER_0_132_892 ();
 sg13g2_fill_4 FILLER_0_132_927 ();
 sg13g2_fill_1 FILLER_0_132_931 ();
 sg13g2_fill_8 FILLER_0_132_942 ();
 sg13g2_fill_4 FILLER_0_132_950 ();
 sg13g2_fill_1 FILLER_0_132_954 ();
 sg13g2_fill_1 FILLER_0_132_963 ();
 sg13g2_fill_1 FILLER_0_132_973 ();
 sg13g2_fill_1 FILLER_0_132_984 ();
 sg13g2_fill_1 FILLER_0_132_994 ();
 sg13g2_fill_2 FILLER_0_132_1000 ();
 sg13g2_fill_4 FILLER_0_132_1007 ();
 sg13g2_fill_1 FILLER_0_132_1011 ();
 sg13g2_fill_2 FILLER_0_132_1017 ();
 sg13g2_fill_1 FILLER_0_132_1019 ();
 sg13g2_fill_4 FILLER_0_132_1025 ();
 sg13g2_fill_8 FILLER_0_132_1039 ();
 sg13g2_fill_4 FILLER_0_132_1047 ();
 sg13g2_fill_2 FILLER_0_132_1051 ();
 sg13g2_fill_2 FILLER_0_132_1068 ();
 sg13g2_fill_4 FILLER_0_132_1075 ();
 sg13g2_fill_2 FILLER_0_132_1079 ();
 sg13g2_fill_8 FILLER_0_132_1111 ();
 sg13g2_fill_8 FILLER_0_132_1119 ();
 sg13g2_fill_8 FILLER_0_132_1127 ();
 sg13g2_fill_8 FILLER_0_132_1135 ();
 sg13g2_fill_8 FILLER_0_132_1143 ();
 sg13g2_fill_8 FILLER_0_132_1151 ();
 sg13g2_fill_8 FILLER_0_132_1159 ();
 sg13g2_fill_8 FILLER_0_132_1167 ();
 sg13g2_fill_8 FILLER_0_132_1175 ();
 sg13g2_fill_8 FILLER_0_132_1183 ();
 sg13g2_fill_8 FILLER_0_132_1191 ();
 sg13g2_fill_8 FILLER_0_132_1199 ();
 sg13g2_fill_8 FILLER_0_132_1207 ();
 sg13g2_fill_8 FILLER_0_132_1215 ();
 sg13g2_fill_4 FILLER_0_132_1223 ();
 sg13g2_fill_1 FILLER_0_132_1227 ();
 sg13g2_fill_8 FILLER_0_133_0 ();
 sg13g2_fill_8 FILLER_0_133_8 ();
 sg13g2_fill_8 FILLER_0_133_16 ();
 sg13g2_fill_8 FILLER_0_133_24 ();
 sg13g2_fill_8 FILLER_0_133_32 ();
 sg13g2_fill_8 FILLER_0_133_40 ();
 sg13g2_fill_8 FILLER_0_133_48 ();
 sg13g2_fill_4 FILLER_0_133_56 ();
 sg13g2_fill_1 FILLER_0_133_90 ();
 sg13g2_fill_1 FILLER_0_133_96 ();
 sg13g2_fill_1 FILLER_0_133_135 ();
 sg13g2_fill_8 FILLER_0_133_162 ();
 sg13g2_fill_8 FILLER_0_133_170 ();
 sg13g2_fill_8 FILLER_0_133_178 ();
 sg13g2_fill_8 FILLER_0_133_186 ();
 sg13g2_fill_8 FILLER_0_133_194 ();
 sg13g2_fill_8 FILLER_0_133_202 ();
 sg13g2_fill_8 FILLER_0_133_210 ();
 sg13g2_fill_8 FILLER_0_133_218 ();
 sg13g2_fill_8 FILLER_0_133_226 ();
 sg13g2_fill_8 FILLER_0_133_234 ();
 sg13g2_fill_4 FILLER_0_133_242 ();
 sg13g2_fill_2 FILLER_0_133_246 ();
 sg13g2_decap_8 FILLER_0_133_283 ();
 sg13g2_fill_2 FILLER_0_133_300 ();
 sg13g2_fill_1 FILLER_0_133_306 ();
 sg13g2_fill_2 FILLER_0_133_317 ();
 sg13g2_fill_2 FILLER_0_133_323 ();
 sg13g2_fill_2 FILLER_0_133_330 ();
 sg13g2_fill_1 FILLER_0_133_332 ();
 sg13g2_fill_1 FILLER_0_133_343 ();
 sg13g2_fill_2 FILLER_0_133_394 ();
 sg13g2_fill_1 FILLER_0_133_396 ();
 sg13g2_fill_2 FILLER_0_133_405 ();
 sg13g2_fill_4 FILLER_0_133_433 ();
 sg13g2_fill_1 FILLER_0_133_437 ();
 sg13g2_fill_4 FILLER_0_133_442 ();
 sg13g2_fill_4 FILLER_0_133_477 ();
 sg13g2_fill_2 FILLER_0_133_481 ();
 sg13g2_fill_1 FILLER_0_133_502 ();
 sg13g2_fill_1 FILLER_0_133_552 ();
 sg13g2_fill_4 FILLER_0_133_567 ();
 sg13g2_fill_2 FILLER_0_133_571 ();
 sg13g2_fill_2 FILLER_0_133_596 ();
 sg13g2_fill_1 FILLER_0_133_598 ();
 sg13g2_fill_1 FILLER_0_133_607 ();
 sg13g2_fill_1 FILLER_0_133_663 ();
 sg13g2_fill_8 FILLER_0_133_691 ();
 sg13g2_fill_2 FILLER_0_133_699 ();
 sg13g2_fill_1 FILLER_0_133_701 ();
 sg13g2_fill_8 FILLER_0_133_711 ();
 sg13g2_fill_8 FILLER_0_133_719 ();
 sg13g2_fill_1 FILLER_0_133_731 ();
 sg13g2_fill_2 FILLER_0_133_737 ();
 sg13g2_fill_1 FILLER_0_133_796 ();
 sg13g2_fill_2 FILLER_0_133_831 ();
 sg13g2_fill_1 FILLER_0_133_833 ();
 sg13g2_fill_4 FILLER_0_133_879 ();
 sg13g2_fill_2 FILLER_0_133_883 ();
 sg13g2_fill_1 FILLER_0_133_911 ();
 sg13g2_fill_2 FILLER_0_133_938 ();
 sg13g2_fill_8 FILLER_0_133_970 ();
 sg13g2_fill_1 FILLER_0_133_978 ();
 sg13g2_fill_8 FILLER_0_133_1005 ();
 sg13g2_fill_8 FILLER_0_133_1013 ();
 sg13g2_fill_4 FILLER_0_133_1026 ();
 sg13g2_fill_2 FILLER_0_133_1030 ();
 sg13g2_fill_8 FILLER_0_133_1042 ();
 sg13g2_fill_4 FILLER_0_133_1050 ();
 sg13g2_fill_4 FILLER_0_133_1068 ();
 sg13g2_fill_2 FILLER_0_133_1098 ();
 sg13g2_fill_8 FILLER_0_133_1104 ();
 sg13g2_fill_8 FILLER_0_133_1112 ();
 sg13g2_fill_8 FILLER_0_133_1120 ();
 sg13g2_fill_8 FILLER_0_133_1128 ();
 sg13g2_fill_8 FILLER_0_133_1136 ();
 sg13g2_fill_8 FILLER_0_133_1144 ();
 sg13g2_fill_8 FILLER_0_133_1152 ();
 sg13g2_fill_8 FILLER_0_133_1160 ();
 sg13g2_fill_8 FILLER_0_133_1168 ();
 sg13g2_fill_8 FILLER_0_133_1176 ();
 sg13g2_fill_8 FILLER_0_133_1184 ();
 sg13g2_fill_8 FILLER_0_133_1192 ();
 sg13g2_fill_8 FILLER_0_133_1200 ();
 sg13g2_fill_8 FILLER_0_133_1208 ();
 sg13g2_fill_8 FILLER_0_133_1216 ();
 sg13g2_fill_4 FILLER_0_133_1224 ();
 sg13g2_fill_8 FILLER_0_134_0 ();
 sg13g2_fill_8 FILLER_0_134_8 ();
 sg13g2_fill_8 FILLER_0_134_16 ();
 sg13g2_fill_8 FILLER_0_134_24 ();
 sg13g2_fill_8 FILLER_0_134_32 ();
 sg13g2_fill_8 FILLER_0_134_40 ();
 sg13g2_fill_8 FILLER_0_134_48 ();
 sg13g2_fill_4 FILLER_0_134_56 ();
 sg13g2_fill_2 FILLER_0_134_100 ();
 sg13g2_fill_2 FILLER_0_134_111 ();
 sg13g2_fill_1 FILLER_0_134_113 ();
 sg13g2_fill_1 FILLER_0_134_136 ();
 sg13g2_fill_1 FILLER_0_134_146 ();
 sg13g2_fill_4 FILLER_0_134_151 ();
 sg13g2_fill_8 FILLER_0_134_160 ();
 sg13g2_fill_8 FILLER_0_134_168 ();
 sg13g2_fill_8 FILLER_0_134_176 ();
 sg13g2_fill_8 FILLER_0_134_184 ();
 sg13g2_fill_8 FILLER_0_134_192 ();
 sg13g2_fill_8 FILLER_0_134_200 ();
 sg13g2_fill_8 FILLER_0_134_208 ();
 sg13g2_fill_8 FILLER_0_134_216 ();
 sg13g2_fill_8 FILLER_0_134_224 ();
 sg13g2_fill_8 FILLER_0_134_232 ();
 sg13g2_fill_4 FILLER_0_134_240 ();
 sg13g2_fill_8 FILLER_0_134_283 ();
 sg13g2_decap_8 FILLER_0_134_291 ();
 sg13g2_fill_8 FILLER_0_134_302 ();
 sg13g2_fill_8 FILLER_0_134_310 ();
 sg13g2_decap_8 FILLER_0_134_318 ();
 sg13g2_fill_4 FILLER_0_134_329 ();
 sg13g2_fill_2 FILLER_0_134_333 ();
 sg13g2_fill_8 FILLER_0_134_339 ();
 sg13g2_fill_1 FILLER_0_134_347 ();
 sg13g2_fill_2 FILLER_0_134_360 ();
 sg13g2_fill_4 FILLER_0_134_388 ();
 sg13g2_fill_2 FILLER_0_134_392 ();
 sg13g2_fill_8 FILLER_0_134_404 ();
 sg13g2_fill_1 FILLER_0_134_412 ();
 sg13g2_fill_1 FILLER_0_134_417 ();
 sg13g2_fill_1 FILLER_0_134_428 ();
 sg13g2_fill_8 FILLER_0_134_433 ();
 sg13g2_fill_8 FILLER_0_134_451 ();
 sg13g2_fill_1 FILLER_0_134_459 ();
 sg13g2_fill_8 FILLER_0_134_464 ();
 sg13g2_fill_2 FILLER_0_134_472 ();
 sg13g2_fill_1 FILLER_0_134_474 ();
 sg13g2_fill_1 FILLER_0_134_501 ();
 sg13g2_fill_2 FILLER_0_134_533 ();
 sg13g2_fill_1 FILLER_0_134_535 ();
 sg13g2_fill_1 FILLER_0_134_540 ();
 sg13g2_fill_1 FILLER_0_134_567 ();
 sg13g2_fill_2 FILLER_0_134_594 ();
 sg13g2_fill_1 FILLER_0_134_596 ();
 sg13g2_fill_1 FILLER_0_134_633 ();
 sg13g2_decap_8 FILLER_0_134_668 ();
 sg13g2_fill_1 FILLER_0_134_679 ();
 sg13g2_decap_8 FILLER_0_134_684 ();
 sg13g2_fill_8 FILLER_0_134_721 ();
 sg13g2_fill_4 FILLER_0_134_729 ();
 sg13g2_fill_1 FILLER_0_134_733 ();
 sg13g2_fill_8 FILLER_0_134_780 ();
 sg13g2_fill_8 FILLER_0_134_788 ();
 sg13g2_fill_2 FILLER_0_134_796 ();
 sg13g2_fill_1 FILLER_0_134_798 ();
 sg13g2_fill_8 FILLER_0_134_822 ();
 sg13g2_fill_8 FILLER_0_134_830 ();
 sg13g2_fill_4 FILLER_0_134_838 ();
 sg13g2_fill_8 FILLER_0_134_895 ();
 sg13g2_fill_8 FILLER_0_134_903 ();
 sg13g2_fill_4 FILLER_0_134_911 ();
 sg13g2_fill_1 FILLER_0_134_915 ();
 sg13g2_fill_2 FILLER_0_134_942 ();
 sg13g2_fill_1 FILLER_0_134_944 ();
 sg13g2_fill_8 FILLER_0_134_976 ();
 sg13g2_fill_2 FILLER_0_134_984 ();
 sg13g2_fill_4 FILLER_0_134_1038 ();
 sg13g2_fill_1 FILLER_0_134_1042 ();
 sg13g2_fill_8 FILLER_0_134_1103 ();
 sg13g2_fill_8 FILLER_0_134_1111 ();
 sg13g2_fill_8 FILLER_0_134_1119 ();
 sg13g2_fill_8 FILLER_0_134_1127 ();
 sg13g2_fill_8 FILLER_0_134_1135 ();
 sg13g2_fill_8 FILLER_0_134_1143 ();
 sg13g2_fill_8 FILLER_0_134_1151 ();
 sg13g2_fill_8 FILLER_0_134_1159 ();
 sg13g2_fill_8 FILLER_0_134_1167 ();
 sg13g2_fill_8 FILLER_0_134_1175 ();
 sg13g2_fill_8 FILLER_0_134_1183 ();
 sg13g2_fill_8 FILLER_0_134_1191 ();
 sg13g2_fill_8 FILLER_0_134_1199 ();
 sg13g2_fill_8 FILLER_0_134_1207 ();
 sg13g2_fill_8 FILLER_0_134_1215 ();
 sg13g2_fill_4 FILLER_0_134_1223 ();
 sg13g2_fill_1 FILLER_0_134_1227 ();
 sg13g2_fill_8 FILLER_0_135_0 ();
 sg13g2_fill_8 FILLER_0_135_8 ();
 sg13g2_fill_8 FILLER_0_135_16 ();
 sg13g2_fill_8 FILLER_0_135_24 ();
 sg13g2_fill_8 FILLER_0_135_32 ();
 sg13g2_fill_8 FILLER_0_135_40 ();
 sg13g2_fill_8 FILLER_0_135_48 ();
 sg13g2_fill_8 FILLER_0_135_56 ();
 sg13g2_fill_2 FILLER_0_135_64 ();
 sg13g2_fill_1 FILLER_0_135_66 ();
 sg13g2_fill_4 FILLER_0_135_71 ();
 sg13g2_fill_1 FILLER_0_135_75 ();
 sg13g2_fill_1 FILLER_0_135_86 ();
 sg13g2_fill_2 FILLER_0_135_96 ();
 sg13g2_fill_1 FILLER_0_135_98 ();
 sg13g2_fill_8 FILLER_0_135_116 ();
 sg13g2_fill_2 FILLER_0_135_124 ();
 sg13g2_fill_8 FILLER_0_135_157 ();
 sg13g2_fill_8 FILLER_0_135_165 ();
 sg13g2_fill_8 FILLER_0_135_173 ();
 sg13g2_fill_8 FILLER_0_135_181 ();
 sg13g2_fill_8 FILLER_0_135_189 ();
 sg13g2_fill_8 FILLER_0_135_197 ();
 sg13g2_fill_8 FILLER_0_135_205 ();
 sg13g2_fill_8 FILLER_0_135_213 ();
 sg13g2_fill_8 FILLER_0_135_221 ();
 sg13g2_decap_8 FILLER_0_135_229 ();
 sg13g2_fill_2 FILLER_0_135_272 ();
 sg13g2_fill_2 FILLER_0_135_289 ();
 sg13g2_fill_1 FILLER_0_135_359 ();
 sg13g2_fill_2 FILLER_0_135_369 ();
 sg13g2_fill_1 FILLER_0_135_371 ();
 sg13g2_fill_4 FILLER_0_135_386 ();
 sg13g2_fill_2 FILLER_0_135_390 ();
 sg13g2_fill_8 FILLER_0_135_396 ();
 sg13g2_fill_8 FILLER_0_135_404 ();
 sg13g2_fill_1 FILLER_0_135_412 ();
 sg13g2_fill_1 FILLER_0_135_418 ();
 sg13g2_fill_1 FILLER_0_135_480 ();
 sg13g2_fill_2 FILLER_0_135_485 ();
 sg13g2_fill_2 FILLER_0_135_492 ();
 sg13g2_fill_2 FILLER_0_135_504 ();
 sg13g2_fill_1 FILLER_0_135_506 ();
 sg13g2_fill_8 FILLER_0_135_537 ();
 sg13g2_fill_4 FILLER_0_135_545 ();
 sg13g2_fill_1 FILLER_0_135_549 ();
 sg13g2_fill_8 FILLER_0_135_554 ();
 sg13g2_fill_8 FILLER_0_135_562 ();
 sg13g2_fill_2 FILLER_0_135_575 ();
 sg13g2_fill_2 FILLER_0_135_581 ();
 sg13g2_fill_1 FILLER_0_135_595 ();
 sg13g2_fill_1 FILLER_0_135_606 ();
 sg13g2_fill_1 FILLER_0_135_633 ();
 sg13g2_fill_1 FILLER_0_135_639 ();
 sg13g2_fill_2 FILLER_0_135_697 ();
 sg13g2_fill_8 FILLER_0_135_704 ();
 sg13g2_fill_8 FILLER_0_135_712 ();
 sg13g2_fill_8 FILLER_0_135_720 ();
 sg13g2_fill_4 FILLER_0_135_728 ();
 sg13g2_fill_2 FILLER_0_135_740 ();
 sg13g2_fill_2 FILLER_0_135_758 ();
 sg13g2_fill_1 FILLER_0_135_760 ();
 sg13g2_fill_2 FILLER_0_135_776 ();
 sg13g2_fill_8 FILLER_0_135_782 ();
 sg13g2_fill_4 FILLER_0_135_790 ();
 sg13g2_fill_2 FILLER_0_135_794 ();
 sg13g2_fill_2 FILLER_0_135_817 ();
 sg13g2_fill_1 FILLER_0_135_819 ();
 sg13g2_fill_2 FILLER_0_135_846 ();
 sg13g2_fill_1 FILLER_0_135_848 ();
 sg13g2_fill_8 FILLER_0_135_894 ();
 sg13g2_fill_2 FILLER_0_135_902 ();
 sg13g2_fill_1 FILLER_0_135_904 ();
 sg13g2_fill_8 FILLER_0_135_913 ();
 sg13g2_fill_1 FILLER_0_135_921 ();
 sg13g2_decap_8 FILLER_0_135_926 ();
 sg13g2_fill_4 FILLER_0_135_943 ();
 sg13g2_fill_2 FILLER_0_135_947 ();
 sg13g2_fill_2 FILLER_0_135_953 ();
 sg13g2_fill_1 FILLER_0_135_955 ();
 sg13g2_fill_8 FILLER_0_135_1088 ();
 sg13g2_fill_8 FILLER_0_135_1096 ();
 sg13g2_fill_8 FILLER_0_135_1104 ();
 sg13g2_fill_8 FILLER_0_135_1112 ();
 sg13g2_fill_8 FILLER_0_135_1120 ();
 sg13g2_fill_8 FILLER_0_135_1128 ();
 sg13g2_fill_8 FILLER_0_135_1136 ();
 sg13g2_fill_8 FILLER_0_135_1144 ();
 sg13g2_fill_8 FILLER_0_135_1152 ();
 sg13g2_fill_8 FILLER_0_135_1160 ();
 sg13g2_fill_8 FILLER_0_135_1168 ();
 sg13g2_fill_8 FILLER_0_135_1176 ();
 sg13g2_fill_8 FILLER_0_135_1184 ();
 sg13g2_fill_8 FILLER_0_135_1192 ();
 sg13g2_fill_8 FILLER_0_135_1200 ();
 sg13g2_fill_8 FILLER_0_135_1208 ();
 sg13g2_fill_8 FILLER_0_135_1216 ();
 sg13g2_fill_4 FILLER_0_135_1224 ();
 sg13g2_fill_8 FILLER_0_136_0 ();
 sg13g2_fill_8 FILLER_0_136_8 ();
 sg13g2_fill_8 FILLER_0_136_16 ();
 sg13g2_fill_8 FILLER_0_136_24 ();
 sg13g2_fill_8 FILLER_0_136_32 ();
 sg13g2_fill_8 FILLER_0_136_40 ();
 sg13g2_fill_8 FILLER_0_136_48 ();
 sg13g2_fill_1 FILLER_0_136_56 ();
 sg13g2_fill_2 FILLER_0_136_83 ();
 sg13g2_fill_2 FILLER_0_136_95 ();
 sg13g2_fill_1 FILLER_0_136_123 ();
 sg13g2_decap_8 FILLER_0_136_132 ();
 sg13g2_fill_8 FILLER_0_136_169 ();
 sg13g2_fill_8 FILLER_0_136_177 ();
 sg13g2_fill_8 FILLER_0_136_185 ();
 sg13g2_fill_8 FILLER_0_136_193 ();
 sg13g2_fill_8 FILLER_0_136_201 ();
 sg13g2_fill_8 FILLER_0_136_209 ();
 sg13g2_fill_8 FILLER_0_136_217 ();
 sg13g2_fill_8 FILLER_0_136_225 ();
 sg13g2_decap_8 FILLER_0_136_233 ();
 sg13g2_fill_1 FILLER_0_136_253 ();
 sg13g2_fill_1 FILLER_0_136_264 ();
 sg13g2_fill_2 FILLER_0_136_291 ();
 sg13g2_fill_1 FILLER_0_136_329 ();
 sg13g2_fill_8 FILLER_0_136_345 ();
 sg13g2_fill_8 FILLER_0_136_353 ();
 sg13g2_decap_8 FILLER_0_136_361 ();
 sg13g2_fill_8 FILLER_0_136_395 ();
 sg13g2_fill_4 FILLER_0_136_433 ();
 sg13g2_fill_1 FILLER_0_136_437 ();
 sg13g2_decap_8 FILLER_0_136_468 ();
 sg13g2_fill_8 FILLER_0_136_506 ();
 sg13g2_fill_4 FILLER_0_136_514 ();
 sg13g2_fill_2 FILLER_0_136_518 ();
 sg13g2_fill_4 FILLER_0_136_535 ();
 sg13g2_fill_1 FILLER_0_136_539 ();
 sg13g2_fill_8 FILLER_0_136_570 ();
 sg13g2_fill_8 FILLER_0_136_578 ();
 sg13g2_fill_8 FILLER_0_136_586 ();
 sg13g2_fill_8 FILLER_0_136_594 ();
 sg13g2_fill_8 FILLER_0_136_602 ();
 sg13g2_fill_1 FILLER_0_136_610 ();
 sg13g2_fill_2 FILLER_0_136_625 ();
 sg13g2_fill_1 FILLER_0_136_627 ();
 sg13g2_fill_1 FILLER_0_136_647 ();
 sg13g2_fill_2 FILLER_0_136_652 ();
 sg13g2_fill_2 FILLER_0_136_685 ();
 sg13g2_fill_2 FILLER_0_136_697 ();
 sg13g2_fill_4 FILLER_0_136_724 ();
 sg13g2_fill_1 FILLER_0_136_728 ();
 sg13g2_fill_8 FILLER_0_136_755 ();
 sg13g2_fill_4 FILLER_0_136_763 ();
 sg13g2_fill_1 FILLER_0_136_793 ();
 sg13g2_fill_1 FILLER_0_136_830 ();
 sg13g2_fill_2 FILLER_0_136_835 ();
 sg13g2_fill_1 FILLER_0_136_837 ();
 sg13g2_fill_2 FILLER_0_136_869 ();
 sg13g2_fill_1 FILLER_0_136_871 ();
 sg13g2_fill_1 FILLER_0_136_886 ();
 sg13g2_fill_4 FILLER_0_136_891 ();
 sg13g2_fill_2 FILLER_0_136_895 ();
 sg13g2_fill_4 FILLER_0_136_907 ();
 sg13g2_fill_2 FILLER_0_136_911 ();
 sg13g2_fill_8 FILLER_0_136_922 ();
 sg13g2_fill_8 FILLER_0_136_930 ();
 sg13g2_fill_8 FILLER_0_136_938 ();
 sg13g2_fill_8 FILLER_0_136_946 ();
 sg13g2_fill_8 FILLER_0_136_954 ();
 sg13g2_fill_8 FILLER_0_136_962 ();
 sg13g2_fill_2 FILLER_0_136_970 ();
 sg13g2_fill_8 FILLER_0_136_976 ();
 sg13g2_fill_8 FILLER_0_136_984 ();
 sg13g2_fill_8 FILLER_0_136_992 ();
 sg13g2_fill_2 FILLER_0_136_1000 ();
 sg13g2_fill_2 FILLER_0_136_1006 ();
 sg13g2_fill_4 FILLER_0_136_1012 ();
 sg13g2_fill_2 FILLER_0_136_1016 ();
 sg13g2_fill_2 FILLER_0_136_1056 ();
 sg13g2_fill_8 FILLER_0_136_1071 ();
 sg13g2_fill_8 FILLER_0_136_1079 ();
 sg13g2_fill_8 FILLER_0_136_1087 ();
 sg13g2_fill_8 FILLER_0_136_1095 ();
 sg13g2_fill_8 FILLER_0_136_1103 ();
 sg13g2_fill_8 FILLER_0_136_1111 ();
 sg13g2_fill_8 FILLER_0_136_1119 ();
 sg13g2_fill_8 FILLER_0_136_1127 ();
 sg13g2_fill_8 FILLER_0_136_1135 ();
 sg13g2_fill_8 FILLER_0_136_1143 ();
 sg13g2_fill_8 FILLER_0_136_1151 ();
 sg13g2_fill_8 FILLER_0_136_1159 ();
 sg13g2_fill_8 FILLER_0_136_1167 ();
 sg13g2_fill_8 FILLER_0_136_1175 ();
 sg13g2_fill_8 FILLER_0_136_1183 ();
 sg13g2_fill_8 FILLER_0_136_1191 ();
 sg13g2_fill_8 FILLER_0_136_1199 ();
 sg13g2_fill_8 FILLER_0_136_1207 ();
 sg13g2_fill_8 FILLER_0_136_1215 ();
 sg13g2_fill_4 FILLER_0_136_1223 ();
 sg13g2_fill_1 FILLER_0_136_1227 ();
 sg13g2_fill_8 FILLER_0_137_0 ();
 sg13g2_fill_8 FILLER_0_137_8 ();
 sg13g2_fill_8 FILLER_0_137_16 ();
 sg13g2_fill_8 FILLER_0_137_24 ();
 sg13g2_fill_4 FILLER_0_137_32 ();
 sg13g2_fill_1 FILLER_0_137_36 ();
 sg13g2_fill_4 FILLER_0_137_41 ();
 sg13g2_fill_1 FILLER_0_137_45 ();
 sg13g2_fill_1 FILLER_0_137_160 ();
 sg13g2_fill_8 FILLER_0_137_166 ();
 sg13g2_fill_8 FILLER_0_137_174 ();
 sg13g2_fill_8 FILLER_0_137_182 ();
 sg13g2_fill_8 FILLER_0_137_190 ();
 sg13g2_fill_8 FILLER_0_137_198 ();
 sg13g2_fill_8 FILLER_0_137_206 ();
 sg13g2_fill_8 FILLER_0_137_214 ();
 sg13g2_fill_8 FILLER_0_137_222 ();
 sg13g2_fill_8 FILLER_0_137_230 ();
 sg13g2_fill_8 FILLER_0_137_238 ();
 sg13g2_fill_4 FILLER_0_137_246 ();
 sg13g2_fill_2 FILLER_0_137_250 ();
 sg13g2_fill_4 FILLER_0_137_293 ();
 sg13g2_fill_4 FILLER_0_137_311 ();
 sg13g2_fill_2 FILLER_0_137_315 ();
 sg13g2_fill_2 FILLER_0_137_327 ();
 sg13g2_fill_1 FILLER_0_137_329 ();
 sg13g2_fill_4 FILLER_0_137_382 ();
 sg13g2_fill_4 FILLER_0_137_435 ();
 sg13g2_fill_2 FILLER_0_137_439 ();
 sg13g2_fill_4 FILLER_0_137_456 ();
 sg13g2_fill_8 FILLER_0_137_468 ();
 sg13g2_fill_8 FILLER_0_137_476 ();
 sg13g2_fill_4 FILLER_0_137_488 ();
 sg13g2_fill_4 FILLER_0_137_511 ();
 sg13g2_fill_1 FILLER_0_137_515 ();
 sg13g2_fill_8 FILLER_0_137_546 ();
 sg13g2_fill_1 FILLER_0_137_554 ();
 sg13g2_fill_1 FILLER_0_137_560 ();
 sg13g2_fill_1 FILLER_0_137_571 ();
 sg13g2_fill_8 FILLER_0_137_576 ();
 sg13g2_fill_8 FILLER_0_137_584 ();
 sg13g2_decap_8 FILLER_0_137_592 ();
 sg13g2_fill_8 FILLER_0_137_625 ();
 sg13g2_fill_8 FILLER_0_137_633 ();
 sg13g2_fill_8 FILLER_0_137_641 ();
 sg13g2_fill_8 FILLER_0_137_649 ();
 sg13g2_fill_8 FILLER_0_137_657 ();
 sg13g2_fill_1 FILLER_0_137_665 ();
 sg13g2_fill_8 FILLER_0_137_670 ();
 sg13g2_fill_1 FILLER_0_137_678 ();
 sg13g2_fill_8 FILLER_0_137_689 ();
 sg13g2_fill_8 FILLER_0_137_697 ();
 sg13g2_fill_2 FILLER_0_137_705 ();
 sg13g2_fill_1 FILLER_0_137_707 ();
 sg13g2_fill_4 FILLER_0_137_713 ();
 sg13g2_fill_1 FILLER_0_137_717 ();
 sg13g2_fill_1 FILLER_0_137_733 ();
 sg13g2_fill_1 FILLER_0_137_769 ();
 sg13g2_fill_2 FILLER_0_137_775 ();
 sg13g2_fill_1 FILLER_0_137_777 ();
 sg13g2_fill_8 FILLER_0_137_782 ();
 sg13g2_decap_8 FILLER_0_137_790 ();
 sg13g2_fill_1 FILLER_0_137_801 ();
 sg13g2_fill_1 FILLER_0_137_806 ();
 sg13g2_fill_2 FILLER_0_137_833 ();
 sg13g2_fill_2 FILLER_0_137_840 ();
 sg13g2_fill_1 FILLER_0_137_842 ();
 sg13g2_fill_2 FILLER_0_137_847 ();
 sg13g2_fill_2 FILLER_0_137_859 ();
 sg13g2_fill_1 FILLER_0_137_861 ();
 sg13g2_fill_2 FILLER_0_137_866 ();
 sg13g2_fill_1 FILLER_0_137_880 ();
 sg13g2_fill_8 FILLER_0_137_937 ();
 sg13g2_fill_8 FILLER_0_137_945 ();
 sg13g2_fill_8 FILLER_0_137_953 ();
 sg13g2_fill_8 FILLER_0_137_961 ();
 sg13g2_fill_8 FILLER_0_137_969 ();
 sg13g2_fill_8 FILLER_0_137_977 ();
 sg13g2_fill_8 FILLER_0_137_985 ();
 sg13g2_fill_8 FILLER_0_137_993 ();
 sg13g2_fill_2 FILLER_0_137_1001 ();
 sg13g2_fill_8 FILLER_0_137_1011 ();
 sg13g2_fill_8 FILLER_0_137_1019 ();
 sg13g2_fill_1 FILLER_0_137_1027 ();
 sg13g2_fill_8 FILLER_0_137_1036 ();
 sg13g2_fill_4 FILLER_0_137_1044 ();
 sg13g2_fill_1 FILLER_0_137_1048 ();
 sg13g2_fill_8 FILLER_0_137_1057 ();
 sg13g2_fill_8 FILLER_0_137_1065 ();
 sg13g2_fill_8 FILLER_0_137_1073 ();
 sg13g2_fill_8 FILLER_0_137_1081 ();
 sg13g2_fill_8 FILLER_0_137_1089 ();
 sg13g2_fill_8 FILLER_0_137_1097 ();
 sg13g2_fill_8 FILLER_0_137_1105 ();
 sg13g2_fill_8 FILLER_0_137_1113 ();
 sg13g2_fill_8 FILLER_0_137_1121 ();
 sg13g2_fill_8 FILLER_0_137_1129 ();
 sg13g2_fill_8 FILLER_0_137_1137 ();
 sg13g2_fill_8 FILLER_0_137_1145 ();
 sg13g2_fill_8 FILLER_0_137_1153 ();
 sg13g2_fill_8 FILLER_0_137_1161 ();
 sg13g2_fill_8 FILLER_0_137_1169 ();
 sg13g2_fill_8 FILLER_0_137_1177 ();
 sg13g2_fill_8 FILLER_0_137_1185 ();
 sg13g2_fill_8 FILLER_0_137_1193 ();
 sg13g2_fill_8 FILLER_0_137_1201 ();
 sg13g2_fill_8 FILLER_0_137_1209 ();
 sg13g2_fill_8 FILLER_0_137_1217 ();
 sg13g2_fill_2 FILLER_0_137_1225 ();
 sg13g2_fill_1 FILLER_0_137_1227 ();
 sg13g2_fill_8 FILLER_0_138_0 ();
 sg13g2_fill_8 FILLER_0_138_8 ();
 sg13g2_fill_8 FILLER_0_138_16 ();
 sg13g2_fill_4 FILLER_0_138_24 ();
 sg13g2_fill_2 FILLER_0_138_28 ();
 sg13g2_fill_4 FILLER_0_138_90 ();
 sg13g2_fill_4 FILLER_0_138_133 ();
 sg13g2_fill_1 FILLER_0_138_145 ();
 sg13g2_fill_2 FILLER_0_138_151 ();
 sg13g2_fill_8 FILLER_0_138_192 ();
 sg13g2_fill_8 FILLER_0_138_200 ();
 sg13g2_fill_8 FILLER_0_138_208 ();
 sg13g2_fill_8 FILLER_0_138_216 ();
 sg13g2_fill_8 FILLER_0_138_224 ();
 sg13g2_fill_8 FILLER_0_138_232 ();
 sg13g2_fill_8 FILLER_0_138_240 ();
 sg13g2_fill_8 FILLER_0_138_248 ();
 sg13g2_fill_4 FILLER_0_138_256 ();
 sg13g2_fill_4 FILLER_0_138_264 ();
 sg13g2_fill_8 FILLER_0_138_272 ();
 sg13g2_fill_8 FILLER_0_138_280 ();
 sg13g2_fill_4 FILLER_0_138_288 ();
 sg13g2_fill_2 FILLER_0_138_292 ();
 sg13g2_fill_8 FILLER_0_138_299 ();
 sg13g2_fill_8 FILLER_0_138_307 ();
 sg13g2_fill_8 FILLER_0_138_315 ();
 sg13g2_fill_4 FILLER_0_138_346 ();
 sg13g2_fill_1 FILLER_0_138_350 ();
 sg13g2_fill_1 FILLER_0_138_413 ();
 sg13g2_fill_4 FILLER_0_138_429 ();
 sg13g2_fill_2 FILLER_0_138_433 ();
 sg13g2_fill_1 FILLER_0_138_445 ();
 sg13g2_fill_8 FILLER_0_138_465 ();
 sg13g2_fill_8 FILLER_0_138_473 ();
 sg13g2_fill_4 FILLER_0_138_481 ();
 sg13g2_fill_2 FILLER_0_138_485 ();
 sg13g2_fill_2 FILLER_0_138_496 ();
 sg13g2_fill_1 FILLER_0_138_595 ();
 sg13g2_fill_1 FILLER_0_138_600 ();
 sg13g2_fill_2 FILLER_0_138_606 ();
 sg13g2_fill_2 FILLER_0_138_634 ();
 sg13g2_fill_2 FILLER_0_138_641 ();
 sg13g2_fill_1 FILLER_0_138_643 ();
 sg13g2_fill_8 FILLER_0_138_648 ();
 sg13g2_fill_8 FILLER_0_138_656 ();
 sg13g2_fill_4 FILLER_0_138_664 ();
 sg13g2_fill_2 FILLER_0_138_668 ();
 sg13g2_fill_4 FILLER_0_138_674 ();
 sg13g2_fill_2 FILLER_0_138_678 ();
 sg13g2_fill_8 FILLER_0_138_695 ();
 sg13g2_fill_1 FILLER_0_138_773 ();
 sg13g2_fill_1 FILLER_0_138_804 ();
 sg13g2_fill_8 FILLER_0_138_820 ();
 sg13g2_fill_8 FILLER_0_138_828 ();
 sg13g2_fill_1 FILLER_0_138_878 ();
 sg13g2_fill_1 FILLER_0_138_905 ();
 sg13g2_fill_2 FILLER_0_138_916 ();
 sg13g2_fill_1 FILLER_0_138_918 ();
 sg13g2_fill_4 FILLER_0_138_945 ();
 sg13g2_fill_8 FILLER_0_138_953 ();
 sg13g2_fill_8 FILLER_0_138_961 ();
 sg13g2_fill_8 FILLER_0_138_969 ();
 sg13g2_fill_8 FILLER_0_138_977 ();
 sg13g2_fill_8 FILLER_0_138_985 ();
 sg13g2_fill_8 FILLER_0_138_993 ();
 sg13g2_fill_8 FILLER_0_138_1001 ();
 sg13g2_fill_8 FILLER_0_138_1009 ();
 sg13g2_fill_8 FILLER_0_138_1017 ();
 sg13g2_fill_8 FILLER_0_138_1025 ();
 sg13g2_fill_8 FILLER_0_138_1033 ();
 sg13g2_fill_8 FILLER_0_138_1041 ();
 sg13g2_fill_8 FILLER_0_138_1049 ();
 sg13g2_fill_8 FILLER_0_138_1057 ();
 sg13g2_fill_8 FILLER_0_138_1065 ();
 sg13g2_fill_8 FILLER_0_138_1073 ();
 sg13g2_fill_8 FILLER_0_138_1081 ();
 sg13g2_fill_8 FILLER_0_138_1089 ();
 sg13g2_fill_8 FILLER_0_138_1097 ();
 sg13g2_fill_8 FILLER_0_138_1105 ();
 sg13g2_fill_8 FILLER_0_138_1113 ();
 sg13g2_fill_8 FILLER_0_138_1121 ();
 sg13g2_fill_8 FILLER_0_138_1129 ();
 sg13g2_fill_8 FILLER_0_138_1137 ();
 sg13g2_fill_8 FILLER_0_138_1145 ();
 sg13g2_fill_8 FILLER_0_138_1153 ();
 sg13g2_fill_8 FILLER_0_138_1161 ();
 sg13g2_fill_8 FILLER_0_138_1169 ();
 sg13g2_fill_8 FILLER_0_138_1177 ();
 sg13g2_fill_8 FILLER_0_138_1185 ();
 sg13g2_fill_8 FILLER_0_138_1193 ();
 sg13g2_fill_8 FILLER_0_138_1201 ();
 sg13g2_fill_8 FILLER_0_138_1209 ();
 sg13g2_fill_8 FILLER_0_138_1217 ();
 sg13g2_fill_2 FILLER_0_138_1225 ();
 sg13g2_fill_1 FILLER_0_138_1227 ();
 sg13g2_fill_8 FILLER_0_139_0 ();
 sg13g2_fill_8 FILLER_0_139_8 ();
 sg13g2_fill_8 FILLER_0_139_16 ();
 sg13g2_fill_8 FILLER_0_139_24 ();
 sg13g2_fill_8 FILLER_0_139_32 ();
 sg13g2_fill_8 FILLER_0_139_40 ();
 sg13g2_fill_4 FILLER_0_139_48 ();
 sg13g2_fill_8 FILLER_0_139_57 ();
 sg13g2_fill_2 FILLER_0_139_65 ();
 sg13g2_fill_4 FILLER_0_139_76 ();
 sg13g2_fill_1 FILLER_0_139_80 ();
 sg13g2_fill_2 FILLER_0_139_107 ();
 sg13g2_fill_4 FILLER_0_139_113 ();
 sg13g2_fill_1 FILLER_0_139_117 ();
 sg13g2_fill_2 FILLER_0_139_122 ();
 sg13g2_fill_2 FILLER_0_139_155 ();
 sg13g2_fill_8 FILLER_0_139_188 ();
 sg13g2_fill_8 FILLER_0_139_196 ();
 sg13g2_fill_8 FILLER_0_139_204 ();
 sg13g2_fill_8 FILLER_0_139_212 ();
 sg13g2_fill_8 FILLER_0_139_220 ();
 sg13g2_fill_8 FILLER_0_139_228 ();
 sg13g2_fill_8 FILLER_0_139_236 ();
 sg13g2_fill_8 FILLER_0_139_244 ();
 sg13g2_fill_8 FILLER_0_139_252 ();
 sg13g2_fill_8 FILLER_0_139_260 ();
 sg13g2_fill_8 FILLER_0_139_268 ();
 sg13g2_fill_4 FILLER_0_139_276 ();
 sg13g2_fill_2 FILLER_0_139_340 ();
 sg13g2_fill_8 FILLER_0_139_346 ();
 sg13g2_fill_2 FILLER_0_139_354 ();
 sg13g2_fill_1 FILLER_0_139_398 ();
 sg13g2_fill_4 FILLER_0_139_444 ();
 sg13g2_fill_1 FILLER_0_139_448 ();
 sg13g2_fill_1 FILLER_0_139_475 ();
 sg13g2_fill_2 FILLER_0_139_552 ();
 sg13g2_fill_1 FILLER_0_139_564 ();
 sg13g2_fill_2 FILLER_0_139_575 ();
 sg13g2_fill_2 FILLER_0_139_587 ();
 sg13g2_fill_2 FILLER_0_139_615 ();
 sg13g2_fill_1 FILLER_0_139_617 ();
 sg13g2_fill_2 FILLER_0_139_622 ();
 sg13g2_fill_2 FILLER_0_139_660 ();
 sg13g2_fill_1 FILLER_0_139_662 ();
 sg13g2_fill_8 FILLER_0_139_693 ();
 sg13g2_fill_8 FILLER_0_139_731 ();
 sg13g2_fill_1 FILLER_0_139_739 ();
 sg13g2_fill_1 FILLER_0_139_748 ();
 sg13g2_fill_2 FILLER_0_139_754 ();
 sg13g2_fill_2 FILLER_0_139_766 ();
 sg13g2_fill_2 FILLER_0_139_772 ();
 sg13g2_fill_8 FILLER_0_139_779 ();
 sg13g2_fill_8 FILLER_0_139_787 ();
 sg13g2_fill_4 FILLER_0_139_795 ();
 sg13g2_fill_4 FILLER_0_139_804 ();
 sg13g2_fill_2 FILLER_0_139_901 ();
 sg13g2_fill_2 FILLER_0_139_918 ();
 sg13g2_decap_8 FILLER_0_139_935 ();
 sg13g2_fill_8 FILLER_0_139_968 ();
 sg13g2_fill_8 FILLER_0_139_976 ();
 sg13g2_fill_8 FILLER_0_139_984 ();
 sg13g2_fill_8 FILLER_0_139_992 ();
 sg13g2_fill_8 FILLER_0_139_1000 ();
 sg13g2_fill_8 FILLER_0_139_1008 ();
 sg13g2_fill_8 FILLER_0_139_1016 ();
 sg13g2_fill_8 FILLER_0_139_1024 ();
 sg13g2_fill_8 FILLER_0_139_1032 ();
 sg13g2_fill_8 FILLER_0_139_1040 ();
 sg13g2_fill_8 FILLER_0_139_1048 ();
 sg13g2_fill_8 FILLER_0_139_1056 ();
 sg13g2_fill_8 FILLER_0_139_1064 ();
 sg13g2_fill_8 FILLER_0_139_1072 ();
 sg13g2_fill_8 FILLER_0_139_1080 ();
 sg13g2_fill_8 FILLER_0_139_1088 ();
 sg13g2_fill_8 FILLER_0_139_1096 ();
 sg13g2_fill_8 FILLER_0_139_1104 ();
 sg13g2_fill_8 FILLER_0_139_1112 ();
 sg13g2_fill_8 FILLER_0_139_1120 ();
 sg13g2_fill_8 FILLER_0_139_1128 ();
 sg13g2_fill_8 FILLER_0_139_1136 ();
 sg13g2_fill_8 FILLER_0_139_1144 ();
 sg13g2_fill_8 FILLER_0_139_1152 ();
 sg13g2_fill_8 FILLER_0_139_1160 ();
 sg13g2_fill_8 FILLER_0_139_1168 ();
 sg13g2_fill_8 FILLER_0_139_1176 ();
 sg13g2_fill_8 FILLER_0_139_1184 ();
 sg13g2_fill_8 FILLER_0_139_1192 ();
 sg13g2_fill_8 FILLER_0_139_1200 ();
 sg13g2_fill_8 FILLER_0_139_1208 ();
 sg13g2_fill_8 FILLER_0_139_1216 ();
 sg13g2_fill_4 FILLER_0_139_1224 ();
 sg13g2_fill_8 FILLER_0_140_0 ();
 sg13g2_fill_8 FILLER_0_140_8 ();
 sg13g2_fill_8 FILLER_0_140_16 ();
 sg13g2_fill_8 FILLER_0_140_24 ();
 sg13g2_fill_8 FILLER_0_140_32 ();
 sg13g2_fill_8 FILLER_0_140_40 ();
 sg13g2_fill_8 FILLER_0_140_78 ();
 sg13g2_fill_8 FILLER_0_140_90 ();
 sg13g2_fill_4 FILLER_0_140_98 ();
 sg13g2_fill_8 FILLER_0_140_107 ();
 sg13g2_decap_8 FILLER_0_140_115 ();
 sg13g2_fill_8 FILLER_0_140_152 ();
 sg13g2_fill_4 FILLER_0_140_160 ();
 sg13g2_fill_1 FILLER_0_140_168 ();
 sg13g2_fill_8 FILLER_0_140_173 ();
 sg13g2_fill_8 FILLER_0_140_181 ();
 sg13g2_fill_8 FILLER_0_140_189 ();
 sg13g2_fill_8 FILLER_0_140_197 ();
 sg13g2_fill_8 FILLER_0_140_205 ();
 sg13g2_fill_8 FILLER_0_140_213 ();
 sg13g2_fill_8 FILLER_0_140_221 ();
 sg13g2_fill_8 FILLER_0_140_229 ();
 sg13g2_fill_8 FILLER_0_140_237 ();
 sg13g2_fill_8 FILLER_0_140_245 ();
 sg13g2_fill_8 FILLER_0_140_253 ();
 sg13g2_fill_2 FILLER_0_140_261 ();
 sg13g2_fill_1 FILLER_0_140_319 ();
 sg13g2_fill_8 FILLER_0_140_351 ();
 sg13g2_fill_8 FILLER_0_140_359 ();
 sg13g2_fill_4 FILLER_0_140_367 ();
 sg13g2_fill_1 FILLER_0_140_371 ();
 sg13g2_fill_8 FILLER_0_140_376 ();
 sg13g2_fill_8 FILLER_0_140_384 ();
 sg13g2_fill_8 FILLER_0_140_392 ();
 sg13g2_fill_8 FILLER_0_140_400 ();
 sg13g2_fill_2 FILLER_0_140_408 ();
 sg13g2_fill_1 FILLER_0_140_410 ();
 sg13g2_fill_8 FILLER_0_140_467 ();
 sg13g2_decap_8 FILLER_0_140_475 ();
 sg13g2_fill_4 FILLER_0_140_486 ();
 sg13g2_fill_2 FILLER_0_140_498 ();
 sg13g2_fill_8 FILLER_0_140_514 ();
 sg13g2_fill_1 FILLER_0_140_522 ();
 sg13g2_fill_2 FILLER_0_140_527 ();
 sg13g2_fill_2 FILLER_0_140_534 ();
 sg13g2_fill_1 FILLER_0_140_536 ();
 sg13g2_fill_2 FILLER_0_140_547 ();
 sg13g2_fill_2 FILLER_0_140_558 ();
 sg13g2_fill_1 FILLER_0_140_604 ();
 sg13g2_fill_2 FILLER_0_140_609 ();
 sg13g2_fill_2 FILLER_0_140_616 ();
 sg13g2_fill_2 FILLER_0_140_628 ();
 sg13g2_fill_2 FILLER_0_140_661 ();
 sg13g2_fill_1 FILLER_0_140_704 ();
 sg13g2_fill_1 FILLER_0_140_709 ();
 sg13g2_fill_8 FILLER_0_140_736 ();
 sg13g2_fill_4 FILLER_0_140_744 ();
 sg13g2_fill_2 FILLER_0_140_753 ();
 sg13g2_fill_2 FILLER_0_140_765 ();
 sg13g2_fill_1 FILLER_0_140_767 ();
 sg13g2_fill_2 FILLER_0_140_794 ();
 sg13g2_fill_1 FILLER_0_140_796 ();
 sg13g2_fill_2 FILLER_0_140_807 ();
 sg13g2_fill_1 FILLER_0_140_819 ();
 sg13g2_fill_8 FILLER_0_140_824 ();
 sg13g2_fill_8 FILLER_0_140_832 ();
 sg13g2_fill_2 FILLER_0_140_840 ();
 sg13g2_fill_1 FILLER_0_140_847 ();
 sg13g2_fill_1 FILLER_0_140_862 ();
 sg13g2_fill_1 FILLER_0_140_873 ();
 sg13g2_fill_2 FILLER_0_140_884 ();
 sg13g2_fill_8 FILLER_0_140_896 ();
 sg13g2_fill_8 FILLER_0_140_904 ();
 sg13g2_fill_4 FILLER_0_140_912 ();
 sg13g2_fill_4 FILLER_0_140_926 ();
 sg13g2_fill_2 FILLER_0_140_930 ();
 sg13g2_fill_8 FILLER_0_140_936 ();
 sg13g2_fill_8 FILLER_0_140_944 ();
 sg13g2_fill_8 FILLER_0_140_952 ();
 sg13g2_fill_8 FILLER_0_140_960 ();
 sg13g2_fill_8 FILLER_0_140_968 ();
 sg13g2_fill_8 FILLER_0_140_976 ();
 sg13g2_fill_8 FILLER_0_140_984 ();
 sg13g2_fill_8 FILLER_0_140_992 ();
 sg13g2_fill_8 FILLER_0_140_1000 ();
 sg13g2_fill_8 FILLER_0_140_1008 ();
 sg13g2_fill_8 FILLER_0_140_1016 ();
 sg13g2_fill_8 FILLER_0_140_1024 ();
 sg13g2_fill_8 FILLER_0_140_1032 ();
 sg13g2_fill_8 FILLER_0_140_1040 ();
 sg13g2_fill_8 FILLER_0_140_1048 ();
 sg13g2_fill_8 FILLER_0_140_1056 ();
 sg13g2_fill_8 FILLER_0_140_1064 ();
 sg13g2_fill_8 FILLER_0_140_1072 ();
 sg13g2_fill_8 FILLER_0_140_1080 ();
 sg13g2_fill_8 FILLER_0_140_1088 ();
 sg13g2_fill_8 FILLER_0_140_1096 ();
 sg13g2_fill_8 FILLER_0_140_1104 ();
 sg13g2_fill_8 FILLER_0_140_1112 ();
 sg13g2_fill_8 FILLER_0_140_1120 ();
 sg13g2_fill_8 FILLER_0_140_1128 ();
 sg13g2_fill_8 FILLER_0_140_1136 ();
 sg13g2_fill_8 FILLER_0_140_1144 ();
 sg13g2_fill_8 FILLER_0_140_1152 ();
 sg13g2_fill_8 FILLER_0_140_1160 ();
 sg13g2_fill_8 FILLER_0_140_1168 ();
 sg13g2_fill_8 FILLER_0_140_1176 ();
 sg13g2_fill_8 FILLER_0_140_1184 ();
 sg13g2_fill_8 FILLER_0_140_1192 ();
 sg13g2_fill_8 FILLER_0_140_1200 ();
 sg13g2_fill_8 FILLER_0_140_1208 ();
 sg13g2_fill_8 FILLER_0_140_1216 ();
 sg13g2_fill_4 FILLER_0_140_1224 ();
 sg13g2_fill_8 FILLER_0_141_0 ();
 sg13g2_fill_8 FILLER_0_141_8 ();
 sg13g2_fill_8 FILLER_0_141_16 ();
 sg13g2_fill_8 FILLER_0_141_24 ();
 sg13g2_fill_4 FILLER_0_141_32 ();
 sg13g2_fill_2 FILLER_0_141_36 ();
 sg13g2_fill_2 FILLER_0_141_81 ();
 sg13g2_fill_1 FILLER_0_141_83 ();
 sg13g2_fill_8 FILLER_0_141_115 ();
 sg13g2_fill_2 FILLER_0_141_123 ();
 sg13g2_fill_2 FILLER_0_141_130 ();
 sg13g2_fill_1 FILLER_0_141_132 ();
 sg13g2_fill_8 FILLER_0_141_141 ();
 sg13g2_fill_8 FILLER_0_141_149 ();
 sg13g2_fill_8 FILLER_0_141_157 ();
 sg13g2_fill_8 FILLER_0_141_165 ();
 sg13g2_fill_8 FILLER_0_141_173 ();
 sg13g2_fill_8 FILLER_0_141_181 ();
 sg13g2_fill_8 FILLER_0_141_189 ();
 sg13g2_fill_8 FILLER_0_141_197 ();
 sg13g2_fill_8 FILLER_0_141_205 ();
 sg13g2_fill_8 FILLER_0_141_213 ();
 sg13g2_fill_8 FILLER_0_141_221 ();
 sg13g2_fill_8 FILLER_0_141_229 ();
 sg13g2_fill_8 FILLER_0_141_237 ();
 sg13g2_fill_8 FILLER_0_141_245 ();
 sg13g2_fill_8 FILLER_0_141_253 ();
 sg13g2_fill_4 FILLER_0_141_261 ();
 sg13g2_fill_2 FILLER_0_141_265 ();
 sg13g2_decap_8 FILLER_0_141_293 ();
 sg13g2_fill_1 FILLER_0_141_304 ();
 sg13g2_fill_1 FILLER_0_141_310 ();
 sg13g2_fill_1 FILLER_0_141_321 ();
 sg13g2_fill_1 FILLER_0_141_326 ();
 sg13g2_fill_2 FILLER_0_141_337 ();
 sg13g2_fill_2 FILLER_0_141_365 ();
 sg13g2_fill_1 FILLER_0_141_367 ();
 sg13g2_fill_8 FILLER_0_141_394 ();
 sg13g2_fill_8 FILLER_0_141_402 ();
 sg13g2_fill_8 FILLER_0_141_410 ();
 sg13g2_fill_8 FILLER_0_141_435 ();
 sg13g2_fill_4 FILLER_0_141_443 ();
 sg13g2_fill_1 FILLER_0_141_447 ();
 sg13g2_fill_8 FILLER_0_141_452 ();
 sg13g2_fill_8 FILLER_0_141_460 ();
 sg13g2_fill_4 FILLER_0_141_468 ();
 sg13g2_fill_2 FILLER_0_141_498 ();
 sg13g2_fill_1 FILLER_0_141_500 ();
 sg13g2_fill_1 FILLER_0_141_514 ();
 sg13g2_fill_2 FILLER_0_141_519 ();
 sg13g2_fill_1 FILLER_0_141_521 ();
 sg13g2_fill_2 FILLER_0_141_526 ();
 sg13g2_fill_1 FILLER_0_141_528 ();
 sg13g2_fill_2 FILLER_0_141_558 ();
 sg13g2_fill_1 FILLER_0_141_572 ();
 sg13g2_fill_4 FILLER_0_141_577 ();
 sg13g2_fill_2 FILLER_0_141_581 ();
 sg13g2_fill_2 FILLER_0_141_593 ();
 sg13g2_fill_1 FILLER_0_141_595 ();
 sg13g2_fill_8 FILLER_0_141_600 ();
 sg13g2_fill_2 FILLER_0_141_608 ();
 sg13g2_fill_8 FILLER_0_141_615 ();
 sg13g2_fill_1 FILLER_0_141_623 ();
 sg13g2_fill_8 FILLER_0_141_666 ();
 sg13g2_fill_4 FILLER_0_141_674 ();
 sg13g2_fill_1 FILLER_0_141_687 ();
 sg13g2_fill_1 FILLER_0_141_713 ();
 sg13g2_fill_1 FILLER_0_141_724 ();
 sg13g2_fill_8 FILLER_0_141_729 ();
 sg13g2_fill_2 FILLER_0_141_737 ();
 sg13g2_fill_2 FILLER_0_141_765 ();
 sg13g2_fill_8 FILLER_0_141_873 ();
 sg13g2_fill_1 FILLER_0_141_881 ();
 sg13g2_fill_4 FILLER_0_141_894 ();
 sg13g2_fill_1 FILLER_0_141_898 ();
 sg13g2_fill_8 FILLER_0_141_904 ();
 sg13g2_fill_4 FILLER_0_141_912 ();
 sg13g2_fill_8 FILLER_0_141_955 ();
 sg13g2_fill_8 FILLER_0_141_963 ();
 sg13g2_fill_8 FILLER_0_141_971 ();
 sg13g2_fill_8 FILLER_0_141_979 ();
 sg13g2_fill_8 FILLER_0_141_987 ();
 sg13g2_fill_8 FILLER_0_141_995 ();
 sg13g2_fill_8 FILLER_0_141_1003 ();
 sg13g2_fill_8 FILLER_0_141_1011 ();
 sg13g2_fill_8 FILLER_0_141_1019 ();
 sg13g2_fill_8 FILLER_0_141_1027 ();
 sg13g2_fill_8 FILLER_0_141_1035 ();
 sg13g2_fill_8 FILLER_0_141_1043 ();
 sg13g2_fill_8 FILLER_0_141_1051 ();
 sg13g2_fill_8 FILLER_0_141_1059 ();
 sg13g2_fill_8 FILLER_0_141_1067 ();
 sg13g2_fill_8 FILLER_0_141_1075 ();
 sg13g2_fill_8 FILLER_0_141_1083 ();
 sg13g2_fill_8 FILLER_0_141_1091 ();
 sg13g2_fill_8 FILLER_0_141_1099 ();
 sg13g2_fill_8 FILLER_0_141_1107 ();
 sg13g2_fill_8 FILLER_0_141_1115 ();
 sg13g2_fill_8 FILLER_0_141_1123 ();
 sg13g2_fill_8 FILLER_0_141_1131 ();
 sg13g2_fill_8 FILLER_0_141_1139 ();
 sg13g2_fill_8 FILLER_0_141_1147 ();
 sg13g2_fill_8 FILLER_0_141_1155 ();
 sg13g2_fill_8 FILLER_0_141_1163 ();
 sg13g2_fill_8 FILLER_0_141_1171 ();
 sg13g2_fill_8 FILLER_0_141_1179 ();
 sg13g2_fill_8 FILLER_0_141_1187 ();
 sg13g2_fill_8 FILLER_0_141_1195 ();
 sg13g2_fill_8 FILLER_0_141_1203 ();
 sg13g2_fill_8 FILLER_0_141_1211 ();
 sg13g2_fill_8 FILLER_0_141_1219 ();
 sg13g2_fill_1 FILLER_0_141_1227 ();
 sg13g2_fill_8 FILLER_0_142_0 ();
 sg13g2_fill_8 FILLER_0_142_8 ();
 sg13g2_fill_8 FILLER_0_142_16 ();
 sg13g2_fill_8 FILLER_0_142_24 ();
 sg13g2_fill_8 FILLER_0_142_32 ();
 sg13g2_decap_8 FILLER_0_142_71 ();
 sg13g2_fill_4 FILLER_0_142_124 ();
 sg13g2_fill_1 FILLER_0_142_128 ();
 sg13g2_fill_8 FILLER_0_142_155 ();
 sg13g2_fill_8 FILLER_0_142_163 ();
 sg13g2_fill_8 FILLER_0_142_171 ();
 sg13g2_fill_8 FILLER_0_142_179 ();
 sg13g2_fill_8 FILLER_0_142_187 ();
 sg13g2_fill_8 FILLER_0_142_195 ();
 sg13g2_fill_8 FILLER_0_142_203 ();
 sg13g2_fill_8 FILLER_0_142_211 ();
 sg13g2_fill_8 FILLER_0_142_219 ();
 sg13g2_fill_8 FILLER_0_142_227 ();
 sg13g2_fill_8 FILLER_0_142_235 ();
 sg13g2_fill_8 FILLER_0_142_243 ();
 sg13g2_fill_8 FILLER_0_142_251 ();
 sg13g2_fill_8 FILLER_0_142_259 ();
 sg13g2_decap_8 FILLER_0_142_267 ();
 sg13g2_fill_8 FILLER_0_142_293 ();
 sg13g2_fill_8 FILLER_0_142_301 ();
 sg13g2_fill_4 FILLER_0_142_309 ();
 sg13g2_fill_1 FILLER_0_142_313 ();
 sg13g2_fill_4 FILLER_0_142_318 ();
 sg13g2_fill_2 FILLER_0_142_330 ();
 sg13g2_fill_4 FILLER_0_142_336 ();
 sg13g2_fill_1 FILLER_0_142_345 ();
 sg13g2_fill_1 FILLER_0_142_350 ();
 sg13g2_fill_4 FILLER_0_142_361 ();
 sg13g2_fill_2 FILLER_0_142_370 ();
 sg13g2_fill_8 FILLER_0_142_434 ();
 sg13g2_decap_8 FILLER_0_142_442 ();
 sg13g2_fill_4 FILLER_0_142_453 ();
 sg13g2_fill_1 FILLER_0_142_457 ();
 sg13g2_decap_8 FILLER_0_142_472 ();
 sg13g2_fill_4 FILLER_0_142_483 ();
 sg13g2_fill_1 FILLER_0_142_497 ();
 sg13g2_fill_2 FILLER_0_142_524 ();
 sg13g2_fill_1 FILLER_0_142_536 ();
 sg13g2_fill_1 FILLER_0_142_542 ();
 sg13g2_fill_8 FILLER_0_142_569 ();
 sg13g2_fill_2 FILLER_0_142_586 ();
 sg13g2_fill_2 FILLER_0_142_592 ();
 sg13g2_fill_1 FILLER_0_142_594 ();
 sg13g2_fill_4 FILLER_0_142_626 ();
 sg13g2_fill_8 FILLER_0_142_661 ();
 sg13g2_decap_8 FILLER_0_142_669 ();
 sg13g2_fill_2 FILLER_0_142_702 ();
 sg13g2_fill_1 FILLER_0_142_709 ();
 sg13g2_fill_2 FILLER_0_142_718 ();
 sg13g2_fill_8 FILLER_0_142_728 ();
 sg13g2_decap_8 FILLER_0_142_736 ();
 sg13g2_fill_4 FILLER_0_142_752 ();
 sg13g2_fill_1 FILLER_0_142_783 ();
 sg13g2_fill_1 FILLER_0_142_794 ();
 sg13g2_fill_1 FILLER_0_142_803 ();
 sg13g2_fill_1 FILLER_0_142_809 ();
 sg13g2_fill_8 FILLER_0_142_827 ();
 sg13g2_fill_8 FILLER_0_142_835 ();
 sg13g2_fill_8 FILLER_0_142_847 ();
 sg13g2_fill_4 FILLER_0_142_855 ();
 sg13g2_fill_2 FILLER_0_142_859 ();
 sg13g2_fill_4 FILLER_0_142_865 ();
 sg13g2_fill_4 FILLER_0_142_873 ();
 sg13g2_fill_8 FILLER_0_142_949 ();
 sg13g2_fill_8 FILLER_0_142_957 ();
 sg13g2_fill_8 FILLER_0_142_965 ();
 sg13g2_fill_8 FILLER_0_142_973 ();
 sg13g2_fill_8 FILLER_0_142_981 ();
 sg13g2_fill_8 FILLER_0_142_989 ();
 sg13g2_fill_8 FILLER_0_142_997 ();
 sg13g2_fill_8 FILLER_0_142_1005 ();
 sg13g2_fill_8 FILLER_0_142_1013 ();
 sg13g2_fill_8 FILLER_0_142_1021 ();
 sg13g2_fill_8 FILLER_0_142_1029 ();
 sg13g2_fill_8 FILLER_0_142_1037 ();
 sg13g2_fill_8 FILLER_0_142_1045 ();
 sg13g2_fill_8 FILLER_0_142_1053 ();
 sg13g2_fill_8 FILLER_0_142_1061 ();
 sg13g2_fill_8 FILLER_0_142_1069 ();
 sg13g2_fill_8 FILLER_0_142_1077 ();
 sg13g2_fill_8 FILLER_0_142_1085 ();
 sg13g2_fill_8 FILLER_0_142_1093 ();
 sg13g2_fill_8 FILLER_0_142_1101 ();
 sg13g2_fill_8 FILLER_0_142_1109 ();
 sg13g2_fill_8 FILLER_0_142_1117 ();
 sg13g2_fill_8 FILLER_0_142_1125 ();
 sg13g2_fill_8 FILLER_0_142_1133 ();
 sg13g2_fill_8 FILLER_0_142_1141 ();
 sg13g2_fill_8 FILLER_0_142_1149 ();
 sg13g2_fill_8 FILLER_0_142_1157 ();
 sg13g2_fill_8 FILLER_0_142_1165 ();
 sg13g2_fill_8 FILLER_0_142_1173 ();
 sg13g2_fill_8 FILLER_0_142_1181 ();
 sg13g2_fill_8 FILLER_0_142_1189 ();
 sg13g2_fill_8 FILLER_0_142_1197 ();
 sg13g2_fill_8 FILLER_0_142_1205 ();
 sg13g2_fill_8 FILLER_0_142_1213 ();
 sg13g2_decap_8 FILLER_0_142_1221 ();
 sg13g2_fill_8 FILLER_0_143_0 ();
 sg13g2_fill_8 FILLER_0_143_8 ();
 sg13g2_fill_8 FILLER_0_143_16 ();
 sg13g2_fill_8 FILLER_0_143_24 ();
 sg13g2_fill_8 FILLER_0_143_32 ();
 sg13g2_fill_8 FILLER_0_143_40 ();
 sg13g2_fill_1 FILLER_0_143_48 ();
 sg13g2_fill_8 FILLER_0_143_53 ();
 sg13g2_fill_8 FILLER_0_143_61 ();
 sg13g2_fill_8 FILLER_0_143_69 ();
 sg13g2_fill_4 FILLER_0_143_77 ();
 sg13g2_fill_2 FILLER_0_143_81 ();
 sg13g2_fill_8 FILLER_0_143_113 ();
 sg13g2_fill_8 FILLER_0_143_121 ();
 sg13g2_fill_4 FILLER_0_143_129 ();
 sg13g2_fill_2 FILLER_0_143_133 ();
 sg13g2_fill_8 FILLER_0_143_139 ();
 sg13g2_fill_8 FILLER_0_143_147 ();
 sg13g2_fill_8 FILLER_0_143_155 ();
 sg13g2_fill_8 FILLER_0_143_163 ();
 sg13g2_fill_8 FILLER_0_143_171 ();
 sg13g2_fill_8 FILLER_0_143_179 ();
 sg13g2_fill_8 FILLER_0_143_187 ();
 sg13g2_fill_8 FILLER_0_143_195 ();
 sg13g2_fill_8 FILLER_0_143_203 ();
 sg13g2_fill_8 FILLER_0_143_211 ();
 sg13g2_fill_8 FILLER_0_143_219 ();
 sg13g2_fill_8 FILLER_0_143_227 ();
 sg13g2_fill_8 FILLER_0_143_235 ();
 sg13g2_fill_8 FILLER_0_143_243 ();
 sg13g2_fill_8 FILLER_0_143_251 ();
 sg13g2_fill_8 FILLER_0_143_259 ();
 sg13g2_fill_2 FILLER_0_143_267 ();
 sg13g2_fill_8 FILLER_0_143_277 ();
 sg13g2_fill_8 FILLER_0_143_285 ();
 sg13g2_fill_8 FILLER_0_143_293 ();
 sg13g2_fill_8 FILLER_0_143_301 ();
 sg13g2_fill_4 FILLER_0_143_309 ();
 sg13g2_fill_2 FILLER_0_143_313 ();
 sg13g2_fill_4 FILLER_0_143_323 ();
 sg13g2_fill_1 FILLER_0_143_327 ();
 sg13g2_fill_2 FILLER_0_143_333 ();
 sg13g2_fill_1 FILLER_0_143_335 ();
 sg13g2_fill_8 FILLER_0_143_341 ();
 sg13g2_fill_2 FILLER_0_143_349 ();
 sg13g2_fill_1 FILLER_0_143_422 ();
 sg13g2_fill_1 FILLER_0_143_480 ();
 sg13g2_fill_1 FILLER_0_143_507 ();
 sg13g2_fill_2 FILLER_0_143_534 ();
 sg13g2_fill_1 FILLER_0_143_541 ();
 sg13g2_fill_2 FILLER_0_143_568 ();
 sg13g2_fill_1 FILLER_0_143_596 ();
 sg13g2_fill_2 FILLER_0_143_601 ();
 sg13g2_fill_2 FILLER_0_143_644 ();
 sg13g2_fill_8 FILLER_0_143_650 ();
 sg13g2_fill_8 FILLER_0_143_658 ();
 sg13g2_fill_8 FILLER_0_143_666 ();
 sg13g2_fill_4 FILLER_0_143_674 ();
 sg13g2_fill_1 FILLER_0_143_678 ();
 sg13g2_fill_4 FILLER_0_143_684 ();
 sg13g2_fill_2 FILLER_0_143_692 ();
 sg13g2_fill_1 FILLER_0_143_704 ();
 sg13g2_fill_8 FILLER_0_143_740 ();
 sg13g2_fill_2 FILLER_0_143_748 ();
 sg13g2_fill_8 FILLER_0_143_776 ();
 sg13g2_fill_2 FILLER_0_143_792 ();
 sg13g2_fill_1 FILLER_0_143_794 ();
 sg13g2_fill_8 FILLER_0_143_821 ();
 sg13g2_fill_8 FILLER_0_143_829 ();
 sg13g2_fill_8 FILLER_0_143_837 ();
 sg13g2_fill_8 FILLER_0_143_845 ();
 sg13g2_fill_1 FILLER_0_143_858 ();
 sg13g2_fill_1 FILLER_0_143_869 ();
 sg13g2_fill_1 FILLER_0_143_922 ();
 sg13g2_fill_8 FILLER_0_143_954 ();
 sg13g2_fill_8 FILLER_0_143_962 ();
 sg13g2_fill_8 FILLER_0_143_970 ();
 sg13g2_fill_8 FILLER_0_143_978 ();
 sg13g2_fill_8 FILLER_0_143_986 ();
 sg13g2_fill_8 FILLER_0_143_994 ();
 sg13g2_fill_8 FILLER_0_143_1002 ();
 sg13g2_fill_8 FILLER_0_143_1010 ();
 sg13g2_fill_8 FILLER_0_143_1018 ();
 sg13g2_fill_8 FILLER_0_143_1026 ();
 sg13g2_fill_8 FILLER_0_143_1034 ();
 sg13g2_fill_8 FILLER_0_143_1042 ();
 sg13g2_fill_8 FILLER_0_143_1050 ();
 sg13g2_fill_8 FILLER_0_143_1058 ();
 sg13g2_fill_8 FILLER_0_143_1066 ();
 sg13g2_fill_8 FILLER_0_143_1074 ();
 sg13g2_fill_8 FILLER_0_143_1082 ();
 sg13g2_fill_8 FILLER_0_143_1090 ();
 sg13g2_fill_8 FILLER_0_143_1098 ();
 sg13g2_fill_8 FILLER_0_143_1106 ();
 sg13g2_fill_8 FILLER_0_143_1114 ();
 sg13g2_fill_8 FILLER_0_143_1122 ();
 sg13g2_fill_8 FILLER_0_143_1130 ();
 sg13g2_fill_8 FILLER_0_143_1138 ();
 sg13g2_fill_8 FILLER_0_143_1146 ();
 sg13g2_fill_8 FILLER_0_143_1154 ();
 sg13g2_fill_8 FILLER_0_143_1162 ();
 sg13g2_fill_8 FILLER_0_143_1170 ();
 sg13g2_fill_8 FILLER_0_143_1178 ();
 sg13g2_fill_8 FILLER_0_143_1186 ();
 sg13g2_fill_8 FILLER_0_143_1194 ();
 sg13g2_fill_8 FILLER_0_143_1202 ();
 sg13g2_fill_8 FILLER_0_143_1210 ();
 sg13g2_fill_8 FILLER_0_143_1218 ();
 sg13g2_fill_2 FILLER_0_143_1226 ();
 sg13g2_fill_8 FILLER_0_144_0 ();
 sg13g2_fill_8 FILLER_0_144_8 ();
 sg13g2_fill_8 FILLER_0_144_16 ();
 sg13g2_fill_8 FILLER_0_144_24 ();
 sg13g2_fill_8 FILLER_0_144_32 ();
 sg13g2_fill_8 FILLER_0_144_40 ();
 sg13g2_fill_8 FILLER_0_144_48 ();
 sg13g2_fill_8 FILLER_0_144_56 ();
 sg13g2_fill_8 FILLER_0_144_64 ();
 sg13g2_fill_8 FILLER_0_144_72 ();
 sg13g2_fill_8 FILLER_0_144_80 ();
 sg13g2_fill_1 FILLER_0_144_88 ();
 sg13g2_fill_2 FILLER_0_144_93 ();
 sg13g2_fill_1 FILLER_0_144_95 ();
 sg13g2_fill_8 FILLER_0_144_100 ();
 sg13g2_fill_8 FILLER_0_144_108 ();
 sg13g2_fill_8 FILLER_0_144_116 ();
 sg13g2_fill_8 FILLER_0_144_124 ();
 sg13g2_fill_8 FILLER_0_144_132 ();
 sg13g2_fill_8 FILLER_0_144_140 ();
 sg13g2_fill_8 FILLER_0_144_148 ();
 sg13g2_fill_8 FILLER_0_144_156 ();
 sg13g2_fill_8 FILLER_0_144_164 ();
 sg13g2_fill_8 FILLER_0_144_172 ();
 sg13g2_fill_8 FILLER_0_144_180 ();
 sg13g2_fill_8 FILLER_0_144_188 ();
 sg13g2_fill_8 FILLER_0_144_196 ();
 sg13g2_fill_8 FILLER_0_144_204 ();
 sg13g2_fill_8 FILLER_0_144_212 ();
 sg13g2_fill_8 FILLER_0_144_220 ();
 sg13g2_fill_8 FILLER_0_144_228 ();
 sg13g2_fill_8 FILLER_0_144_236 ();
 sg13g2_fill_8 FILLER_0_144_244 ();
 sg13g2_fill_8 FILLER_0_144_252 ();
 sg13g2_fill_8 FILLER_0_144_260 ();
 sg13g2_fill_4 FILLER_0_144_268 ();
 sg13g2_fill_1 FILLER_0_144_297 ();
 sg13g2_fill_2 FILLER_0_144_303 ();
 sg13g2_fill_1 FILLER_0_144_305 ();
 sg13g2_fill_2 FILLER_0_144_332 ();
 sg13g2_fill_4 FILLER_0_144_360 ();
 sg13g2_fill_4 FILLER_0_144_369 ();
 sg13g2_fill_2 FILLER_0_144_377 ();
 sg13g2_fill_4 FILLER_0_144_383 ();
 sg13g2_fill_2 FILLER_0_144_397 ();
 sg13g2_fill_4 FILLER_0_144_404 ();
 sg13g2_fill_1 FILLER_0_144_412 ();
 sg13g2_fill_1 FILLER_0_144_423 ();
 sg13g2_fill_1 FILLER_0_144_429 ();
 sg13g2_fill_1 FILLER_0_144_434 ();
 sg13g2_fill_1 FILLER_0_144_440 ();
 sg13g2_fill_1 FILLER_0_144_467 ();
 sg13g2_fill_4 FILLER_0_144_480 ();
 sg13g2_fill_2 FILLER_0_144_484 ();
 sg13g2_fill_2 FILLER_0_144_510 ();
 sg13g2_fill_1 FILLER_0_144_512 ();
 sg13g2_fill_2 FILLER_0_144_528 ();
 sg13g2_fill_4 FILLER_0_144_543 ();
 sg13g2_decap_8 FILLER_0_144_551 ();
 sg13g2_fill_8 FILLER_0_144_562 ();
 sg13g2_fill_8 FILLER_0_144_570 ();
 sg13g2_fill_8 FILLER_0_144_578 ();
 sg13g2_decap_8 FILLER_0_144_586 ();
 sg13g2_fill_4 FILLER_0_144_601 ();
 sg13g2_fill_1 FILLER_0_144_605 ();
 sg13g2_fill_2 FILLER_0_144_629 ();
 sg13g2_fill_4 FILLER_0_144_657 ();
 sg13g2_fill_1 FILLER_0_144_661 ();
 sg13g2_fill_4 FILLER_0_144_670 ();
 sg13g2_fill_2 FILLER_0_144_674 ();
 sg13g2_fill_4 FILLER_0_144_753 ();
 sg13g2_fill_2 FILLER_0_144_757 ();
 sg13g2_fill_8 FILLER_0_144_763 ();
 sg13g2_fill_8 FILLER_0_144_771 ();
 sg13g2_fill_4 FILLER_0_144_779 ();
 sg13g2_fill_8 FILLER_0_144_791 ();
 sg13g2_fill_8 FILLER_0_144_799 ();
 sg13g2_fill_2 FILLER_0_144_807 ();
 sg13g2_fill_4 FILLER_0_144_835 ();
 sg13g2_fill_2 FILLER_0_144_839 ();
 sg13g2_fill_2 FILLER_0_144_846 ();
 sg13g2_fill_2 FILLER_0_144_874 ();
 sg13g2_fill_1 FILLER_0_144_876 ();
 sg13g2_fill_4 FILLER_0_144_881 ();
 sg13g2_fill_1 FILLER_0_144_895 ();
 sg13g2_fill_1 FILLER_0_144_911 ();
 sg13g2_fill_1 FILLER_0_144_937 ();
 sg13g2_fill_8 FILLER_0_144_946 ();
 sg13g2_fill_8 FILLER_0_144_954 ();
 sg13g2_fill_8 FILLER_0_144_962 ();
 sg13g2_fill_8 FILLER_0_144_970 ();
 sg13g2_fill_8 FILLER_0_144_978 ();
 sg13g2_fill_8 FILLER_0_144_986 ();
 sg13g2_fill_8 FILLER_0_144_994 ();
 sg13g2_fill_8 FILLER_0_144_1002 ();
 sg13g2_fill_8 FILLER_0_144_1010 ();
 sg13g2_fill_8 FILLER_0_144_1018 ();
 sg13g2_fill_8 FILLER_0_144_1026 ();
 sg13g2_fill_8 FILLER_0_144_1034 ();
 sg13g2_fill_8 FILLER_0_144_1042 ();
 sg13g2_fill_8 FILLER_0_144_1050 ();
 sg13g2_fill_8 FILLER_0_144_1058 ();
 sg13g2_fill_8 FILLER_0_144_1066 ();
 sg13g2_fill_8 FILLER_0_144_1074 ();
 sg13g2_fill_8 FILLER_0_144_1082 ();
 sg13g2_fill_8 FILLER_0_144_1090 ();
 sg13g2_fill_8 FILLER_0_144_1098 ();
 sg13g2_fill_8 FILLER_0_144_1106 ();
 sg13g2_fill_8 FILLER_0_144_1114 ();
 sg13g2_fill_8 FILLER_0_144_1122 ();
 sg13g2_fill_8 FILLER_0_144_1130 ();
 sg13g2_fill_8 FILLER_0_144_1138 ();
 sg13g2_fill_8 FILLER_0_144_1146 ();
 sg13g2_fill_8 FILLER_0_144_1154 ();
 sg13g2_fill_8 FILLER_0_144_1162 ();
 sg13g2_fill_8 FILLER_0_144_1170 ();
 sg13g2_fill_8 FILLER_0_144_1178 ();
 sg13g2_fill_8 FILLER_0_144_1186 ();
 sg13g2_fill_8 FILLER_0_144_1194 ();
 sg13g2_fill_8 FILLER_0_144_1202 ();
 sg13g2_fill_8 FILLER_0_144_1210 ();
 sg13g2_fill_8 FILLER_0_144_1218 ();
 sg13g2_fill_2 FILLER_0_144_1226 ();
 sg13g2_fill_8 FILLER_0_145_0 ();
 sg13g2_fill_8 FILLER_0_145_8 ();
 sg13g2_fill_8 FILLER_0_145_16 ();
 sg13g2_fill_8 FILLER_0_145_24 ();
 sg13g2_fill_8 FILLER_0_145_32 ();
 sg13g2_fill_8 FILLER_0_145_40 ();
 sg13g2_fill_8 FILLER_0_145_48 ();
 sg13g2_fill_8 FILLER_0_145_56 ();
 sg13g2_fill_8 FILLER_0_145_64 ();
 sg13g2_fill_8 FILLER_0_145_72 ();
 sg13g2_fill_8 FILLER_0_145_80 ();
 sg13g2_fill_8 FILLER_0_145_88 ();
 sg13g2_fill_8 FILLER_0_145_96 ();
 sg13g2_fill_8 FILLER_0_145_104 ();
 sg13g2_fill_8 FILLER_0_145_112 ();
 sg13g2_fill_8 FILLER_0_145_120 ();
 sg13g2_fill_8 FILLER_0_145_128 ();
 sg13g2_fill_8 FILLER_0_145_136 ();
 sg13g2_fill_8 FILLER_0_145_144 ();
 sg13g2_fill_8 FILLER_0_145_152 ();
 sg13g2_fill_8 FILLER_0_145_160 ();
 sg13g2_fill_8 FILLER_0_145_168 ();
 sg13g2_fill_8 FILLER_0_145_176 ();
 sg13g2_fill_8 FILLER_0_145_184 ();
 sg13g2_fill_8 FILLER_0_145_192 ();
 sg13g2_fill_8 FILLER_0_145_200 ();
 sg13g2_fill_8 FILLER_0_145_208 ();
 sg13g2_fill_8 FILLER_0_145_216 ();
 sg13g2_fill_8 FILLER_0_145_224 ();
 sg13g2_fill_8 FILLER_0_145_232 ();
 sg13g2_fill_8 FILLER_0_145_240 ();
 sg13g2_fill_4 FILLER_0_145_248 ();
 sg13g2_fill_2 FILLER_0_145_252 ();
 sg13g2_fill_4 FILLER_0_145_336 ();
 sg13g2_fill_8 FILLER_0_145_344 ();
 sg13g2_fill_4 FILLER_0_145_352 ();
 sg13g2_fill_8 FILLER_0_145_366 ();
 sg13g2_fill_4 FILLER_0_145_374 ();
 sg13g2_fill_8 FILLER_0_145_393 ();
 sg13g2_fill_8 FILLER_0_145_401 ();
 sg13g2_fill_8 FILLER_0_145_409 ();
 sg13g2_fill_8 FILLER_0_145_417 ();
 sg13g2_fill_2 FILLER_0_145_425 ();
 sg13g2_fill_1 FILLER_0_145_427 ();
 sg13g2_fill_2 FILLER_0_145_454 ();
 sg13g2_fill_1 FILLER_0_145_456 ();
 sg13g2_fill_8 FILLER_0_145_476 ();
 sg13g2_fill_8 FILLER_0_145_484 ();
 sg13g2_fill_8 FILLER_0_145_492 ();
 sg13g2_fill_8 FILLER_0_145_500 ();
 sg13g2_fill_8 FILLER_0_145_508 ();
 sg13g2_fill_8 FILLER_0_145_516 ();
 sg13g2_decap_8 FILLER_0_145_524 ();
 sg13g2_fill_2 FILLER_0_145_561 ();
 sg13g2_fill_1 FILLER_0_145_577 ();
 sg13g2_fill_1 FILLER_0_145_582 ();
 sg13g2_fill_2 FILLER_0_145_602 ();
 sg13g2_fill_8 FILLER_0_145_608 ();
 sg13g2_fill_8 FILLER_0_145_616 ();
 sg13g2_fill_2 FILLER_0_145_624 ();
 sg13g2_fill_1 FILLER_0_145_626 ();
 sg13g2_fill_2 FILLER_0_145_663 ();
 sg13g2_fill_2 FILLER_0_145_705 ();
 sg13g2_fill_1 FILLER_0_145_711 ();
 sg13g2_fill_2 FILLER_0_145_720 ();
 sg13g2_fill_1 FILLER_0_145_722 ();
 sg13g2_fill_2 FILLER_0_145_727 ();
 sg13g2_fill_1 FILLER_0_145_729 ();
 sg13g2_fill_8 FILLER_0_145_744 ();
 sg13g2_fill_4 FILLER_0_145_752 ();
 sg13g2_fill_1 FILLER_0_145_756 ();
 sg13g2_fill_1 FILLER_0_145_779 ();
 sg13g2_fill_1 FILLER_0_145_806 ();
 sg13g2_fill_1 FILLER_0_145_811 ();
 sg13g2_fill_1 FILLER_0_145_826 ();
 sg13g2_fill_2 FILLER_0_145_857 ();
 sg13g2_fill_2 FILLER_0_145_874 ();
 sg13g2_fill_1 FILLER_0_145_876 ();
 sg13g2_fill_4 FILLER_0_145_896 ();
 sg13g2_fill_1 FILLER_0_145_905 ();
 sg13g2_fill_8 FILLER_0_145_918 ();
 sg13g2_fill_8 FILLER_0_145_926 ();
 sg13g2_fill_8 FILLER_0_145_934 ();
 sg13g2_fill_8 FILLER_0_145_942 ();
 sg13g2_fill_8 FILLER_0_145_950 ();
 sg13g2_fill_8 FILLER_0_145_958 ();
 sg13g2_fill_8 FILLER_0_145_966 ();
 sg13g2_fill_8 FILLER_0_145_974 ();
 sg13g2_fill_8 FILLER_0_145_982 ();
 sg13g2_fill_8 FILLER_0_145_990 ();
 sg13g2_fill_8 FILLER_0_145_998 ();
 sg13g2_fill_8 FILLER_0_145_1006 ();
 sg13g2_fill_8 FILLER_0_145_1014 ();
 sg13g2_fill_8 FILLER_0_145_1022 ();
 sg13g2_fill_8 FILLER_0_145_1030 ();
 sg13g2_fill_8 FILLER_0_145_1038 ();
 sg13g2_fill_8 FILLER_0_145_1046 ();
 sg13g2_fill_8 FILLER_0_145_1054 ();
 sg13g2_fill_8 FILLER_0_145_1062 ();
 sg13g2_fill_8 FILLER_0_145_1070 ();
 sg13g2_fill_8 FILLER_0_145_1078 ();
 sg13g2_fill_8 FILLER_0_145_1086 ();
 sg13g2_fill_8 FILLER_0_145_1094 ();
 sg13g2_fill_8 FILLER_0_145_1102 ();
 sg13g2_fill_8 FILLER_0_145_1110 ();
 sg13g2_fill_8 FILLER_0_145_1118 ();
 sg13g2_fill_8 FILLER_0_145_1126 ();
 sg13g2_fill_8 FILLER_0_145_1134 ();
 sg13g2_fill_8 FILLER_0_145_1142 ();
 sg13g2_fill_8 FILLER_0_145_1150 ();
 sg13g2_fill_8 FILLER_0_145_1158 ();
 sg13g2_fill_8 FILLER_0_145_1166 ();
 sg13g2_fill_8 FILLER_0_145_1174 ();
 sg13g2_fill_8 FILLER_0_145_1182 ();
 sg13g2_fill_8 FILLER_0_145_1190 ();
 sg13g2_fill_8 FILLER_0_145_1198 ();
 sg13g2_fill_8 FILLER_0_145_1206 ();
 sg13g2_fill_8 FILLER_0_145_1214 ();
 sg13g2_fill_4 FILLER_0_145_1222 ();
 sg13g2_fill_2 FILLER_0_145_1226 ();
 sg13g2_fill_8 FILLER_0_146_0 ();
 sg13g2_fill_8 FILLER_0_146_8 ();
 sg13g2_fill_8 FILLER_0_146_16 ();
 sg13g2_fill_8 FILLER_0_146_24 ();
 sg13g2_fill_8 FILLER_0_146_32 ();
 sg13g2_fill_8 FILLER_0_146_40 ();
 sg13g2_fill_8 FILLER_0_146_48 ();
 sg13g2_fill_8 FILLER_0_146_56 ();
 sg13g2_fill_8 FILLER_0_146_64 ();
 sg13g2_fill_8 FILLER_0_146_72 ();
 sg13g2_fill_8 FILLER_0_146_80 ();
 sg13g2_fill_8 FILLER_0_146_88 ();
 sg13g2_fill_8 FILLER_0_146_96 ();
 sg13g2_fill_8 FILLER_0_146_104 ();
 sg13g2_fill_8 FILLER_0_146_112 ();
 sg13g2_fill_8 FILLER_0_146_120 ();
 sg13g2_fill_8 FILLER_0_146_128 ();
 sg13g2_fill_8 FILLER_0_146_136 ();
 sg13g2_fill_8 FILLER_0_146_144 ();
 sg13g2_fill_8 FILLER_0_146_152 ();
 sg13g2_fill_8 FILLER_0_146_160 ();
 sg13g2_fill_8 FILLER_0_146_168 ();
 sg13g2_fill_8 FILLER_0_146_176 ();
 sg13g2_fill_8 FILLER_0_146_184 ();
 sg13g2_fill_8 FILLER_0_146_192 ();
 sg13g2_fill_8 FILLER_0_146_200 ();
 sg13g2_fill_8 FILLER_0_146_208 ();
 sg13g2_fill_8 FILLER_0_146_216 ();
 sg13g2_fill_8 FILLER_0_146_224 ();
 sg13g2_fill_8 FILLER_0_146_232 ();
 sg13g2_fill_8 FILLER_0_146_240 ();
 sg13g2_fill_8 FILLER_0_146_248 ();
 sg13g2_fill_4 FILLER_0_146_256 ();
 sg13g2_fill_2 FILLER_0_146_260 ();
 sg13g2_fill_2 FILLER_0_146_266 ();
 sg13g2_fill_1 FILLER_0_146_268 ();
 sg13g2_fill_1 FILLER_0_146_305 ();
 sg13g2_fill_2 FILLER_0_146_331 ();
 sg13g2_fill_1 FILLER_0_146_333 ();
 sg13g2_fill_2 FILLER_0_146_360 ();
 sg13g2_fill_2 FILLER_0_146_372 ();
 sg13g2_fill_1 FILLER_0_146_374 ();
 sg13g2_fill_1 FILLER_0_146_385 ();
 sg13g2_fill_2 FILLER_0_146_412 ();
 sg13g2_fill_1 FILLER_0_146_414 ();
 sg13g2_fill_2 FILLER_0_146_420 ();
 sg13g2_fill_1 FILLER_0_146_422 ();
 sg13g2_fill_1 FILLER_0_146_454 ();
 sg13g2_fill_2 FILLER_0_146_481 ();
 sg13g2_fill_1 FILLER_0_146_483 ();
 sg13g2_fill_4 FILLER_0_146_510 ();
 sg13g2_fill_2 FILLER_0_146_580 ();
 sg13g2_fill_1 FILLER_0_146_586 ();
 sg13g2_decap_8 FILLER_0_146_613 ();
 sg13g2_fill_2 FILLER_0_146_635 ();
 sg13g2_fill_1 FILLER_0_146_637 ();
 sg13g2_fill_4 FILLER_0_146_642 ();
 sg13g2_fill_8 FILLER_0_146_650 ();
 sg13g2_fill_4 FILLER_0_146_658 ();
 sg13g2_fill_2 FILLER_0_146_693 ();
 sg13g2_fill_2 FILLER_0_146_705 ();
 sg13g2_fill_1 FILLER_0_146_707 ();
 sg13g2_fill_2 FILLER_0_146_734 ();
 sg13g2_fill_1 FILLER_0_146_736 ();
 sg13g2_fill_2 FILLER_0_146_747 ();
 sg13g2_fill_1 FILLER_0_146_749 ();
 sg13g2_fill_1 FILLER_0_146_812 ();
 sg13g2_fill_1 FILLER_0_146_839 ();
 sg13g2_fill_1 FILLER_0_146_844 ();
 sg13g2_fill_1 FILLER_0_146_850 ();
 sg13g2_fill_2 FILLER_0_146_885 ();
 sg13g2_fill_1 FILLER_0_146_887 ();
 sg13g2_fill_2 FILLER_0_146_914 ();
 sg13g2_fill_8 FILLER_0_146_931 ();
 sg13g2_fill_8 FILLER_0_146_939 ();
 sg13g2_fill_8 FILLER_0_146_947 ();
 sg13g2_fill_8 FILLER_0_146_955 ();
 sg13g2_fill_8 FILLER_0_146_963 ();
 sg13g2_fill_8 FILLER_0_146_971 ();
 sg13g2_fill_8 FILLER_0_146_979 ();
 sg13g2_fill_8 FILLER_0_146_987 ();
 sg13g2_fill_8 FILLER_0_146_995 ();
 sg13g2_fill_8 FILLER_0_146_1003 ();
 sg13g2_fill_8 FILLER_0_146_1011 ();
 sg13g2_fill_8 FILLER_0_146_1019 ();
 sg13g2_fill_8 FILLER_0_146_1027 ();
 sg13g2_fill_8 FILLER_0_146_1035 ();
 sg13g2_fill_8 FILLER_0_146_1043 ();
 sg13g2_fill_8 FILLER_0_146_1051 ();
 sg13g2_fill_8 FILLER_0_146_1059 ();
 sg13g2_fill_8 FILLER_0_146_1067 ();
 sg13g2_fill_8 FILLER_0_146_1075 ();
 sg13g2_fill_8 FILLER_0_146_1083 ();
 sg13g2_fill_8 FILLER_0_146_1091 ();
 sg13g2_fill_8 FILLER_0_146_1099 ();
 sg13g2_fill_8 FILLER_0_146_1107 ();
 sg13g2_fill_8 FILLER_0_146_1115 ();
 sg13g2_fill_8 FILLER_0_146_1123 ();
 sg13g2_fill_8 FILLER_0_146_1131 ();
 sg13g2_fill_8 FILLER_0_146_1139 ();
 sg13g2_fill_8 FILLER_0_146_1147 ();
 sg13g2_fill_8 FILLER_0_146_1155 ();
 sg13g2_fill_8 FILLER_0_146_1163 ();
 sg13g2_fill_8 FILLER_0_146_1171 ();
 sg13g2_fill_8 FILLER_0_146_1179 ();
 sg13g2_fill_8 FILLER_0_146_1187 ();
 sg13g2_fill_8 FILLER_0_146_1195 ();
 sg13g2_fill_8 FILLER_0_146_1203 ();
 sg13g2_fill_8 FILLER_0_146_1211 ();
 sg13g2_fill_8 FILLER_0_146_1219 ();
 sg13g2_fill_1 FILLER_0_146_1227 ();
 sg13g2_fill_8 FILLER_0_147_0 ();
 sg13g2_fill_8 FILLER_0_147_8 ();
 sg13g2_fill_8 FILLER_0_147_16 ();
 sg13g2_fill_8 FILLER_0_147_24 ();
 sg13g2_fill_8 FILLER_0_147_32 ();
 sg13g2_fill_8 FILLER_0_147_40 ();
 sg13g2_fill_8 FILLER_0_147_48 ();
 sg13g2_fill_8 FILLER_0_147_56 ();
 sg13g2_fill_8 FILLER_0_147_64 ();
 sg13g2_fill_8 FILLER_0_147_72 ();
 sg13g2_fill_8 FILLER_0_147_80 ();
 sg13g2_fill_8 FILLER_0_147_88 ();
 sg13g2_fill_8 FILLER_0_147_96 ();
 sg13g2_fill_8 FILLER_0_147_104 ();
 sg13g2_fill_8 FILLER_0_147_112 ();
 sg13g2_fill_8 FILLER_0_147_120 ();
 sg13g2_fill_8 FILLER_0_147_128 ();
 sg13g2_fill_8 FILLER_0_147_136 ();
 sg13g2_fill_8 FILLER_0_147_144 ();
 sg13g2_fill_8 FILLER_0_147_152 ();
 sg13g2_fill_8 FILLER_0_147_160 ();
 sg13g2_fill_8 FILLER_0_147_168 ();
 sg13g2_fill_8 FILLER_0_147_176 ();
 sg13g2_fill_8 FILLER_0_147_184 ();
 sg13g2_fill_8 FILLER_0_147_192 ();
 sg13g2_fill_8 FILLER_0_147_200 ();
 sg13g2_fill_8 FILLER_0_147_208 ();
 sg13g2_fill_8 FILLER_0_147_216 ();
 sg13g2_fill_8 FILLER_0_147_224 ();
 sg13g2_fill_8 FILLER_0_147_232 ();
 sg13g2_fill_8 FILLER_0_147_240 ();
 sg13g2_fill_8 FILLER_0_147_248 ();
 sg13g2_fill_2 FILLER_0_147_256 ();
 sg13g2_fill_1 FILLER_0_147_258 ();
 sg13g2_fill_8 FILLER_0_147_263 ();
 sg13g2_fill_4 FILLER_0_147_271 ();
 sg13g2_fill_8 FILLER_0_147_280 ();
 sg13g2_fill_2 FILLER_0_147_288 ();
 sg13g2_fill_1 FILLER_0_147_290 ();
 sg13g2_fill_8 FILLER_0_147_295 ();
 sg13g2_fill_8 FILLER_0_147_303 ();
 sg13g2_fill_4 FILLER_0_147_311 ();
 sg13g2_fill_2 FILLER_0_147_315 ();
 sg13g2_fill_8 FILLER_0_147_321 ();
 sg13g2_fill_2 FILLER_0_147_329 ();
 sg13g2_fill_1 FILLER_0_147_331 ();
 sg13g2_fill_1 FILLER_0_147_377 ();
 sg13g2_fill_1 FILLER_0_147_462 ();
 sg13g2_fill_1 FILLER_0_147_473 ();
 sg13g2_fill_1 FILLER_0_147_478 ();
 sg13g2_fill_1 FILLER_0_147_489 ();
 sg13g2_fill_1 FILLER_0_147_495 ();
 sg13g2_fill_2 FILLER_0_147_548 ();
 sg13g2_fill_1 FILLER_0_147_550 ();
 sg13g2_fill_1 FILLER_0_147_555 ();
 sg13g2_fill_1 FILLER_0_147_561 ();
 sg13g2_fill_2 FILLER_0_147_588 ();
 sg13g2_fill_1 FILLER_0_147_616 ();
 sg13g2_fill_4 FILLER_0_147_625 ();
 sg13g2_fill_8 FILLER_0_147_660 ();
 sg13g2_fill_4 FILLER_0_147_668 ();
 sg13g2_fill_1 FILLER_0_147_676 ();
 sg13g2_fill_8 FILLER_0_147_681 ();
 sg13g2_fill_4 FILLER_0_147_689 ();
 sg13g2_fill_2 FILLER_0_147_693 ();
 sg13g2_fill_2 FILLER_0_147_705 ();
 sg13g2_fill_1 FILLER_0_147_707 ();
 sg13g2_fill_1 FILLER_0_147_712 ();
 sg13g2_fill_1 FILLER_0_147_718 ();
 sg13g2_fill_1 FILLER_0_147_729 ();
 sg13g2_fill_1 FILLER_0_147_756 ();
 sg13g2_fill_2 FILLER_0_147_762 ();
 sg13g2_fill_1 FILLER_0_147_772 ();
 sg13g2_fill_2 FILLER_0_147_777 ();
 sg13g2_fill_1 FILLER_0_147_784 ();
 sg13g2_fill_2 FILLER_0_147_790 ();
 sg13g2_fill_1 FILLER_0_147_802 ();
 sg13g2_fill_2 FILLER_0_147_815 ();
 sg13g2_decap_8 FILLER_0_147_830 ();
 sg13g2_fill_4 FILLER_0_147_847 ();
 sg13g2_fill_2 FILLER_0_147_851 ();
 sg13g2_fill_8 FILLER_0_147_861 ();
 sg13g2_fill_1 FILLER_0_147_869 ();
 sg13g2_fill_8 FILLER_0_147_948 ();
 sg13g2_fill_8 FILLER_0_147_956 ();
 sg13g2_fill_8 FILLER_0_147_964 ();
 sg13g2_fill_8 FILLER_0_147_972 ();
 sg13g2_fill_8 FILLER_0_147_980 ();
 sg13g2_fill_8 FILLER_0_147_988 ();
 sg13g2_fill_8 FILLER_0_147_996 ();
 sg13g2_fill_8 FILLER_0_147_1004 ();
 sg13g2_fill_8 FILLER_0_147_1012 ();
 sg13g2_fill_8 FILLER_0_147_1020 ();
 sg13g2_fill_8 FILLER_0_147_1028 ();
 sg13g2_fill_8 FILLER_0_147_1036 ();
 sg13g2_fill_8 FILLER_0_147_1044 ();
 sg13g2_fill_8 FILLER_0_147_1052 ();
 sg13g2_fill_8 FILLER_0_147_1060 ();
 sg13g2_fill_8 FILLER_0_147_1068 ();
 sg13g2_fill_8 FILLER_0_147_1076 ();
 sg13g2_fill_8 FILLER_0_147_1084 ();
 sg13g2_fill_8 FILLER_0_147_1092 ();
 sg13g2_fill_8 FILLER_0_147_1100 ();
 sg13g2_fill_8 FILLER_0_147_1108 ();
 sg13g2_fill_8 FILLER_0_147_1116 ();
 sg13g2_fill_8 FILLER_0_147_1124 ();
 sg13g2_fill_8 FILLER_0_147_1132 ();
 sg13g2_fill_8 FILLER_0_147_1140 ();
 sg13g2_fill_8 FILLER_0_147_1148 ();
 sg13g2_fill_8 FILLER_0_147_1156 ();
 sg13g2_fill_8 FILLER_0_147_1164 ();
 sg13g2_fill_8 FILLER_0_147_1172 ();
 sg13g2_fill_8 FILLER_0_147_1180 ();
 sg13g2_fill_8 FILLER_0_147_1188 ();
 sg13g2_fill_8 FILLER_0_147_1196 ();
 sg13g2_fill_8 FILLER_0_147_1204 ();
 sg13g2_fill_8 FILLER_0_147_1212 ();
 sg13g2_fill_8 FILLER_0_147_1220 ();
 sg13g2_fill_8 FILLER_0_148_0 ();
 sg13g2_fill_8 FILLER_0_148_8 ();
 sg13g2_fill_8 FILLER_0_148_16 ();
 sg13g2_fill_8 FILLER_0_148_24 ();
 sg13g2_fill_8 FILLER_0_148_32 ();
 sg13g2_fill_8 FILLER_0_148_40 ();
 sg13g2_fill_8 FILLER_0_148_48 ();
 sg13g2_fill_8 FILLER_0_148_56 ();
 sg13g2_fill_8 FILLER_0_148_64 ();
 sg13g2_fill_8 FILLER_0_148_72 ();
 sg13g2_fill_8 FILLER_0_148_80 ();
 sg13g2_fill_8 FILLER_0_148_88 ();
 sg13g2_fill_8 FILLER_0_148_96 ();
 sg13g2_fill_8 FILLER_0_148_104 ();
 sg13g2_fill_8 FILLER_0_148_112 ();
 sg13g2_fill_8 FILLER_0_148_120 ();
 sg13g2_fill_8 FILLER_0_148_128 ();
 sg13g2_fill_8 FILLER_0_148_136 ();
 sg13g2_fill_8 FILLER_0_148_144 ();
 sg13g2_fill_8 FILLER_0_148_152 ();
 sg13g2_fill_8 FILLER_0_148_160 ();
 sg13g2_fill_8 FILLER_0_148_168 ();
 sg13g2_fill_8 FILLER_0_148_176 ();
 sg13g2_fill_8 FILLER_0_148_184 ();
 sg13g2_fill_8 FILLER_0_148_192 ();
 sg13g2_fill_8 FILLER_0_148_200 ();
 sg13g2_fill_8 FILLER_0_148_208 ();
 sg13g2_fill_8 FILLER_0_148_216 ();
 sg13g2_fill_8 FILLER_0_148_224 ();
 sg13g2_fill_8 FILLER_0_148_232 ();
 sg13g2_fill_8 FILLER_0_148_240 ();
 sg13g2_fill_8 FILLER_0_148_248 ();
 sg13g2_fill_8 FILLER_0_148_256 ();
 sg13g2_fill_8 FILLER_0_148_264 ();
 sg13g2_fill_8 FILLER_0_148_272 ();
 sg13g2_fill_8 FILLER_0_148_280 ();
 sg13g2_fill_8 FILLER_0_148_288 ();
 sg13g2_fill_8 FILLER_0_148_296 ();
 sg13g2_fill_8 FILLER_0_148_304 ();
 sg13g2_fill_8 FILLER_0_148_312 ();
 sg13g2_fill_8 FILLER_0_148_320 ();
 sg13g2_fill_8 FILLER_0_148_328 ();
 sg13g2_fill_4 FILLER_0_148_336 ();
 sg13g2_fill_4 FILLER_0_148_345 ();
 sg13g2_fill_2 FILLER_0_148_353 ();
 sg13g2_fill_1 FILLER_0_148_355 ();
 sg13g2_fill_2 FILLER_0_148_405 ();
 sg13g2_fill_1 FILLER_0_148_407 ();
 sg13g2_fill_4 FILLER_0_148_444 ();
 sg13g2_fill_8 FILLER_0_148_474 ();
 sg13g2_fill_2 FILLER_0_148_482 ();
 sg13g2_fill_1 FILLER_0_148_484 ();
 sg13g2_fill_1 FILLER_0_148_495 ();
 sg13g2_fill_2 FILLER_0_148_501 ();
 sg13g2_fill_4 FILLER_0_148_507 ();
 sg13g2_fill_4 FILLER_0_148_516 ();
 sg13g2_fill_2 FILLER_0_148_556 ();
 sg13g2_fill_2 FILLER_0_148_584 ();
 sg13g2_fill_2 FILLER_0_148_596 ();
 sg13g2_fill_4 FILLER_0_148_602 ();
 sg13g2_fill_2 FILLER_0_148_632 ();
 sg13g2_fill_8 FILLER_0_148_648 ();
 sg13g2_fill_8 FILLER_0_148_656 ();
 sg13g2_fill_8 FILLER_0_148_664 ();
 sg13g2_fill_2 FILLER_0_148_672 ();
 sg13g2_fill_2 FILLER_0_148_705 ();
 sg13g2_fill_1 FILLER_0_148_707 ();
 sg13g2_fill_1 FILLER_0_148_739 ();
 sg13g2_fill_8 FILLER_0_148_744 ();
 sg13g2_fill_4 FILLER_0_148_752 ();
 sg13g2_fill_2 FILLER_0_148_756 ();
 sg13g2_fill_4 FILLER_0_148_763 ();
 sg13g2_fill_1 FILLER_0_148_767 ();
 sg13g2_fill_4 FILLER_0_148_778 ();
 sg13g2_fill_1 FILLER_0_148_782 ();
 sg13g2_fill_2 FILLER_0_148_792 ();
 sg13g2_fill_1 FILLER_0_148_794 ();
 sg13g2_fill_4 FILLER_0_148_805 ();
 sg13g2_fill_2 FILLER_0_148_809 ();
 sg13g2_fill_4 FILLER_0_148_826 ();
 sg13g2_fill_1 FILLER_0_148_830 ();
 sg13g2_fill_8 FILLER_0_148_835 ();
 sg13g2_fill_8 FILLER_0_148_843 ();
 sg13g2_fill_4 FILLER_0_148_851 ();
 sg13g2_fill_2 FILLER_0_148_855 ();
 sg13g2_fill_8 FILLER_0_148_869 ();
 sg13g2_fill_1 FILLER_0_148_877 ();
 sg13g2_fill_8 FILLER_0_148_947 ();
 sg13g2_fill_8 FILLER_0_148_955 ();
 sg13g2_fill_8 FILLER_0_148_963 ();
 sg13g2_fill_8 FILLER_0_148_971 ();
 sg13g2_fill_8 FILLER_0_148_979 ();
 sg13g2_fill_8 FILLER_0_148_987 ();
 sg13g2_fill_8 FILLER_0_148_995 ();
 sg13g2_fill_8 FILLER_0_148_1003 ();
 sg13g2_fill_8 FILLER_0_148_1011 ();
 sg13g2_fill_8 FILLER_0_148_1019 ();
 sg13g2_fill_8 FILLER_0_148_1027 ();
 sg13g2_fill_8 FILLER_0_148_1035 ();
 sg13g2_fill_8 FILLER_0_148_1043 ();
 sg13g2_fill_8 FILLER_0_148_1051 ();
 sg13g2_fill_8 FILLER_0_148_1059 ();
 sg13g2_fill_8 FILLER_0_148_1067 ();
 sg13g2_fill_8 FILLER_0_148_1075 ();
 sg13g2_fill_8 FILLER_0_148_1083 ();
 sg13g2_fill_8 FILLER_0_148_1091 ();
 sg13g2_fill_8 FILLER_0_148_1099 ();
 sg13g2_fill_8 FILLER_0_148_1107 ();
 sg13g2_fill_8 FILLER_0_148_1115 ();
 sg13g2_fill_8 FILLER_0_148_1123 ();
 sg13g2_fill_8 FILLER_0_148_1131 ();
 sg13g2_fill_8 FILLER_0_148_1139 ();
 sg13g2_fill_8 FILLER_0_148_1147 ();
 sg13g2_fill_8 FILLER_0_148_1155 ();
 sg13g2_fill_8 FILLER_0_148_1163 ();
 sg13g2_fill_8 FILLER_0_148_1171 ();
 sg13g2_fill_8 FILLER_0_148_1179 ();
 sg13g2_fill_8 FILLER_0_148_1187 ();
 sg13g2_fill_8 FILLER_0_148_1195 ();
 sg13g2_fill_8 FILLER_0_148_1203 ();
 sg13g2_fill_8 FILLER_0_148_1211 ();
 sg13g2_fill_8 FILLER_0_148_1219 ();
 sg13g2_fill_1 FILLER_0_148_1227 ();
 sg13g2_fill_8 FILLER_0_149_0 ();
 sg13g2_fill_8 FILLER_0_149_8 ();
 sg13g2_fill_8 FILLER_0_149_16 ();
 sg13g2_fill_8 FILLER_0_149_24 ();
 sg13g2_fill_8 FILLER_0_149_32 ();
 sg13g2_fill_8 FILLER_0_149_40 ();
 sg13g2_fill_8 FILLER_0_149_48 ();
 sg13g2_fill_8 FILLER_0_149_56 ();
 sg13g2_fill_8 FILLER_0_149_64 ();
 sg13g2_fill_8 FILLER_0_149_72 ();
 sg13g2_fill_8 FILLER_0_149_80 ();
 sg13g2_fill_8 FILLER_0_149_88 ();
 sg13g2_fill_8 FILLER_0_149_96 ();
 sg13g2_fill_8 FILLER_0_149_104 ();
 sg13g2_fill_8 FILLER_0_149_112 ();
 sg13g2_fill_8 FILLER_0_149_120 ();
 sg13g2_fill_8 FILLER_0_149_128 ();
 sg13g2_fill_8 FILLER_0_149_136 ();
 sg13g2_fill_8 FILLER_0_149_144 ();
 sg13g2_fill_8 FILLER_0_149_152 ();
 sg13g2_fill_8 FILLER_0_149_160 ();
 sg13g2_fill_8 FILLER_0_149_168 ();
 sg13g2_fill_8 FILLER_0_149_176 ();
 sg13g2_fill_8 FILLER_0_149_184 ();
 sg13g2_fill_8 FILLER_0_149_192 ();
 sg13g2_fill_8 FILLER_0_149_200 ();
 sg13g2_fill_8 FILLER_0_149_208 ();
 sg13g2_fill_8 FILLER_0_149_216 ();
 sg13g2_fill_8 FILLER_0_149_224 ();
 sg13g2_fill_8 FILLER_0_149_232 ();
 sg13g2_fill_8 FILLER_0_149_240 ();
 sg13g2_fill_8 FILLER_0_149_248 ();
 sg13g2_fill_8 FILLER_0_149_256 ();
 sg13g2_fill_8 FILLER_0_149_264 ();
 sg13g2_fill_8 FILLER_0_149_272 ();
 sg13g2_fill_8 FILLER_0_149_280 ();
 sg13g2_fill_8 FILLER_0_149_288 ();
 sg13g2_fill_8 FILLER_0_149_296 ();
 sg13g2_fill_8 FILLER_0_149_304 ();
 sg13g2_fill_8 FILLER_0_149_312 ();
 sg13g2_fill_8 FILLER_0_149_320 ();
 sg13g2_fill_8 FILLER_0_149_328 ();
 sg13g2_fill_8 FILLER_0_149_336 ();
 sg13g2_fill_8 FILLER_0_149_344 ();
 sg13g2_fill_8 FILLER_0_149_352 ();
 sg13g2_fill_8 FILLER_0_149_360 ();
 sg13g2_fill_8 FILLER_0_149_368 ();
 sg13g2_fill_2 FILLER_0_149_376 ();
 sg13g2_fill_1 FILLER_0_149_378 ();
 sg13g2_fill_8 FILLER_0_149_383 ();
 sg13g2_fill_1 FILLER_0_149_391 ();
 sg13g2_fill_1 FILLER_0_149_396 ();
 sg13g2_fill_8 FILLER_0_149_401 ();
 sg13g2_fill_2 FILLER_0_149_409 ();
 sg13g2_fill_1 FILLER_0_149_411 ();
 sg13g2_fill_4 FILLER_0_149_425 ();
 sg13g2_fill_2 FILLER_0_149_429 ();
 sg13g2_fill_8 FILLER_0_149_441 ();
 sg13g2_fill_1 FILLER_0_149_449 ();
 sg13g2_fill_1 FILLER_0_149_459 ();
 sg13g2_fill_8 FILLER_0_149_478 ();
 sg13g2_decap_8 FILLER_0_149_486 ();
 sg13g2_fill_2 FILLER_0_149_501 ();
 sg13g2_fill_1 FILLER_0_149_503 ();
 sg13g2_fill_8 FILLER_0_149_514 ();
 sg13g2_fill_4 FILLER_0_149_522 ();
 sg13g2_fill_1 FILLER_0_149_526 ();
 sg13g2_decap_8 FILLER_0_149_535 ();
 sg13g2_fill_8 FILLER_0_149_546 ();
 sg13g2_fill_4 FILLER_0_149_554 ();
 sg13g2_fill_2 FILLER_0_149_573 ();
 sg13g2_fill_1 FILLER_0_149_575 ();
 sg13g2_fill_2 FILLER_0_149_585 ();
 sg13g2_fill_1 FILLER_0_149_587 ();
 sg13g2_fill_4 FILLER_0_149_608 ();
 sg13g2_fill_1 FILLER_0_149_612 ();
 sg13g2_fill_8 FILLER_0_149_617 ();
 sg13g2_fill_2 FILLER_0_149_625 ();
 sg13g2_fill_4 FILLER_0_149_662 ();
 sg13g2_fill_2 FILLER_0_149_666 ();
 sg13g2_fill_1 FILLER_0_149_694 ();
 sg13g2_fill_1 FILLER_0_149_705 ();
 sg13g2_fill_1 FILLER_0_149_715 ();
 sg13g2_fill_2 FILLER_0_149_735 ();
 sg13g2_fill_1 FILLER_0_149_737 ();
 sg13g2_fill_4 FILLER_0_149_746 ();
 sg13g2_fill_1 FILLER_0_149_750 ();
 sg13g2_decap_8 FILLER_0_149_777 ();
 sg13g2_fill_8 FILLER_0_149_837 ();
 sg13g2_fill_4 FILLER_0_149_845 ();
 sg13g2_fill_1 FILLER_0_149_849 ();
 sg13g2_fill_8 FILLER_0_149_876 ();
 sg13g2_fill_8 FILLER_0_149_884 ();
 sg13g2_fill_2 FILLER_0_149_892 ();
 sg13g2_fill_4 FILLER_0_149_898 ();
 sg13g2_fill_8 FILLER_0_149_906 ();
 sg13g2_fill_2 FILLER_0_149_914 ();
 sg13g2_fill_1 FILLER_0_149_916 ();
 sg13g2_fill_4 FILLER_0_149_922 ();
 sg13g2_fill_2 FILLER_0_149_926 ();
 sg13g2_fill_8 FILLER_0_149_936 ();
 sg13g2_fill_8 FILLER_0_149_944 ();
 sg13g2_fill_8 FILLER_0_149_952 ();
 sg13g2_fill_8 FILLER_0_149_960 ();
 sg13g2_fill_8 FILLER_0_149_968 ();
 sg13g2_fill_8 FILLER_0_149_976 ();
 sg13g2_fill_8 FILLER_0_149_984 ();
 sg13g2_fill_8 FILLER_0_149_992 ();
 sg13g2_fill_8 FILLER_0_149_1000 ();
 sg13g2_fill_8 FILLER_0_149_1008 ();
 sg13g2_fill_8 FILLER_0_149_1016 ();
 sg13g2_fill_8 FILLER_0_149_1024 ();
 sg13g2_fill_8 FILLER_0_149_1032 ();
 sg13g2_fill_8 FILLER_0_149_1040 ();
 sg13g2_fill_8 FILLER_0_149_1048 ();
 sg13g2_fill_8 FILLER_0_149_1056 ();
 sg13g2_fill_8 FILLER_0_149_1064 ();
 sg13g2_fill_8 FILLER_0_149_1072 ();
 sg13g2_fill_8 FILLER_0_149_1080 ();
 sg13g2_fill_8 FILLER_0_149_1088 ();
 sg13g2_fill_8 FILLER_0_149_1096 ();
 sg13g2_fill_8 FILLER_0_149_1104 ();
 sg13g2_fill_8 FILLER_0_149_1112 ();
 sg13g2_fill_8 FILLER_0_149_1120 ();
 sg13g2_fill_8 FILLER_0_149_1128 ();
 sg13g2_fill_8 FILLER_0_149_1136 ();
 sg13g2_fill_8 FILLER_0_149_1144 ();
 sg13g2_fill_8 FILLER_0_149_1152 ();
 sg13g2_fill_8 FILLER_0_149_1160 ();
 sg13g2_fill_8 FILLER_0_149_1168 ();
 sg13g2_fill_8 FILLER_0_149_1176 ();
 sg13g2_fill_8 FILLER_0_149_1184 ();
 sg13g2_fill_8 FILLER_0_149_1192 ();
 sg13g2_fill_8 FILLER_0_149_1200 ();
 sg13g2_fill_8 FILLER_0_149_1208 ();
 sg13g2_fill_8 FILLER_0_149_1216 ();
 sg13g2_fill_4 FILLER_0_149_1224 ();
 sg13g2_fill_8 FILLER_0_150_0 ();
 sg13g2_fill_8 FILLER_0_150_8 ();
 sg13g2_fill_8 FILLER_0_150_16 ();
 sg13g2_fill_8 FILLER_0_150_24 ();
 sg13g2_fill_8 FILLER_0_150_32 ();
 sg13g2_fill_8 FILLER_0_150_40 ();
 sg13g2_fill_8 FILLER_0_150_48 ();
 sg13g2_fill_8 FILLER_0_150_56 ();
 sg13g2_fill_8 FILLER_0_150_64 ();
 sg13g2_fill_8 FILLER_0_150_72 ();
 sg13g2_fill_8 FILLER_0_150_80 ();
 sg13g2_fill_8 FILLER_0_150_88 ();
 sg13g2_fill_8 FILLER_0_150_96 ();
 sg13g2_fill_8 FILLER_0_150_104 ();
 sg13g2_fill_8 FILLER_0_150_112 ();
 sg13g2_fill_8 FILLER_0_150_120 ();
 sg13g2_fill_8 FILLER_0_150_128 ();
 sg13g2_fill_8 FILLER_0_150_136 ();
 sg13g2_fill_8 FILLER_0_150_144 ();
 sg13g2_fill_8 FILLER_0_150_152 ();
 sg13g2_fill_8 FILLER_0_150_160 ();
 sg13g2_fill_8 FILLER_0_150_168 ();
 sg13g2_fill_8 FILLER_0_150_176 ();
 sg13g2_fill_8 FILLER_0_150_184 ();
 sg13g2_fill_8 FILLER_0_150_192 ();
 sg13g2_fill_8 FILLER_0_150_200 ();
 sg13g2_fill_8 FILLER_0_150_208 ();
 sg13g2_fill_8 FILLER_0_150_216 ();
 sg13g2_fill_8 FILLER_0_150_224 ();
 sg13g2_fill_8 FILLER_0_150_232 ();
 sg13g2_fill_8 FILLER_0_150_240 ();
 sg13g2_fill_8 FILLER_0_150_248 ();
 sg13g2_fill_8 FILLER_0_150_256 ();
 sg13g2_fill_8 FILLER_0_150_264 ();
 sg13g2_fill_8 FILLER_0_150_272 ();
 sg13g2_fill_8 FILLER_0_150_280 ();
 sg13g2_fill_8 FILLER_0_150_288 ();
 sg13g2_fill_8 FILLER_0_150_296 ();
 sg13g2_fill_8 FILLER_0_150_304 ();
 sg13g2_fill_8 FILLER_0_150_312 ();
 sg13g2_fill_8 FILLER_0_150_320 ();
 sg13g2_fill_8 FILLER_0_150_328 ();
 sg13g2_fill_8 FILLER_0_150_336 ();
 sg13g2_fill_8 FILLER_0_150_344 ();
 sg13g2_fill_8 FILLER_0_150_352 ();
 sg13g2_fill_8 FILLER_0_150_360 ();
 sg13g2_fill_8 FILLER_0_150_368 ();
 sg13g2_fill_8 FILLER_0_150_376 ();
 sg13g2_fill_8 FILLER_0_150_384 ();
 sg13g2_fill_8 FILLER_0_150_392 ();
 sg13g2_fill_8 FILLER_0_150_400 ();
 sg13g2_fill_8 FILLER_0_150_408 ();
 sg13g2_fill_8 FILLER_0_150_416 ();
 sg13g2_fill_8 FILLER_0_150_424 ();
 sg13g2_fill_2 FILLER_0_150_442 ();
 sg13g2_fill_8 FILLER_0_150_474 ();
 sg13g2_fill_4 FILLER_0_150_482 ();
 sg13g2_fill_1 FILLER_0_150_486 ();
 sg13g2_fill_4 FILLER_0_150_513 ();
 sg13g2_decap_8 FILLER_0_150_521 ();
 sg13g2_fill_4 FILLER_0_150_537 ();
 sg13g2_fill_2 FILLER_0_150_541 ();
 sg13g2_fill_2 FILLER_0_150_553 ();
 sg13g2_fill_1 FILLER_0_150_555 ();
 sg13g2_fill_2 FILLER_0_150_576 ();
 sg13g2_fill_8 FILLER_0_150_586 ();
 sg13g2_fill_2 FILLER_0_150_594 ();
 sg13g2_fill_1 FILLER_0_150_596 ();
 sg13g2_fill_2 FILLER_0_150_601 ();
 sg13g2_fill_4 FILLER_0_150_608 ();
 sg13g2_fill_2 FILLER_0_150_612 ();
 sg13g2_fill_4 FILLER_0_150_627 ();
 sg13g2_fill_1 FILLER_0_150_631 ();
 sg13g2_fill_8 FILLER_0_150_647 ();
 sg13g2_fill_8 FILLER_0_150_655 ();
 sg13g2_fill_4 FILLER_0_150_663 ();
 sg13g2_fill_2 FILLER_0_150_667 ();
 sg13g2_fill_8 FILLER_0_150_681 ();
 sg13g2_fill_8 FILLER_0_150_689 ();
 sg13g2_fill_2 FILLER_0_150_697 ();
 sg13g2_fill_1 FILLER_0_150_699 ();
 sg13g2_fill_8 FILLER_0_150_710 ();
 sg13g2_fill_1 FILLER_0_150_718 ();
 sg13g2_fill_8 FILLER_0_150_729 ();
 sg13g2_fill_4 FILLER_0_150_737 ();
 sg13g2_fill_1 FILLER_0_150_741 ();
 sg13g2_fill_2 FILLER_0_150_812 ();
 sg13g2_fill_2 FILLER_0_150_844 ();
 sg13g2_fill_8 FILLER_0_150_892 ();
 sg13g2_fill_8 FILLER_0_150_900 ();
 sg13g2_decap_8 FILLER_0_150_908 ();
 sg13g2_fill_8 FILLER_0_150_933 ();
 sg13g2_fill_8 FILLER_0_150_941 ();
 sg13g2_fill_8 FILLER_0_150_949 ();
 sg13g2_fill_8 FILLER_0_150_957 ();
 sg13g2_fill_8 FILLER_0_150_965 ();
 sg13g2_fill_8 FILLER_0_150_973 ();
 sg13g2_fill_8 FILLER_0_150_981 ();
 sg13g2_fill_8 FILLER_0_150_989 ();
 sg13g2_fill_8 FILLER_0_150_997 ();
 sg13g2_fill_8 FILLER_0_150_1005 ();
 sg13g2_fill_8 FILLER_0_150_1013 ();
 sg13g2_fill_8 FILLER_0_150_1021 ();
 sg13g2_fill_8 FILLER_0_150_1029 ();
 sg13g2_fill_8 FILLER_0_150_1037 ();
 sg13g2_fill_8 FILLER_0_150_1045 ();
 sg13g2_fill_8 FILLER_0_150_1053 ();
 sg13g2_fill_8 FILLER_0_150_1061 ();
 sg13g2_fill_8 FILLER_0_150_1069 ();
 sg13g2_fill_8 FILLER_0_150_1077 ();
 sg13g2_fill_8 FILLER_0_150_1085 ();
 sg13g2_fill_8 FILLER_0_150_1093 ();
 sg13g2_fill_8 FILLER_0_150_1101 ();
 sg13g2_fill_8 FILLER_0_150_1109 ();
 sg13g2_fill_8 FILLER_0_150_1117 ();
 sg13g2_fill_8 FILLER_0_150_1125 ();
 sg13g2_fill_8 FILLER_0_150_1133 ();
 sg13g2_fill_8 FILLER_0_150_1141 ();
 sg13g2_fill_8 FILLER_0_150_1149 ();
 sg13g2_fill_8 FILLER_0_150_1157 ();
 sg13g2_fill_8 FILLER_0_150_1165 ();
 sg13g2_fill_8 FILLER_0_150_1173 ();
 sg13g2_fill_8 FILLER_0_150_1181 ();
 sg13g2_fill_8 FILLER_0_150_1189 ();
 sg13g2_fill_8 FILLER_0_150_1197 ();
 sg13g2_fill_8 FILLER_0_150_1205 ();
 sg13g2_fill_8 FILLER_0_150_1213 ();
 sg13g2_decap_8 FILLER_0_150_1221 ();
 sg13g2_fill_8 FILLER_0_151_0 ();
 sg13g2_fill_8 FILLER_0_151_8 ();
 sg13g2_fill_8 FILLER_0_151_16 ();
 sg13g2_fill_8 FILLER_0_151_24 ();
 sg13g2_fill_8 FILLER_0_151_32 ();
 sg13g2_fill_8 FILLER_0_151_40 ();
 sg13g2_fill_8 FILLER_0_151_48 ();
 sg13g2_fill_8 FILLER_0_151_56 ();
 sg13g2_fill_8 FILLER_0_151_64 ();
 sg13g2_fill_8 FILLER_0_151_72 ();
 sg13g2_fill_8 FILLER_0_151_80 ();
 sg13g2_fill_8 FILLER_0_151_88 ();
 sg13g2_fill_8 FILLER_0_151_96 ();
 sg13g2_fill_8 FILLER_0_151_104 ();
 sg13g2_fill_8 FILLER_0_151_112 ();
 sg13g2_fill_8 FILLER_0_151_120 ();
 sg13g2_fill_8 FILLER_0_151_128 ();
 sg13g2_fill_8 FILLER_0_151_136 ();
 sg13g2_fill_8 FILLER_0_151_144 ();
 sg13g2_fill_8 FILLER_0_151_152 ();
 sg13g2_fill_8 FILLER_0_151_160 ();
 sg13g2_fill_8 FILLER_0_151_168 ();
 sg13g2_fill_8 FILLER_0_151_176 ();
 sg13g2_fill_8 FILLER_0_151_184 ();
 sg13g2_fill_8 FILLER_0_151_192 ();
 sg13g2_fill_8 FILLER_0_151_200 ();
 sg13g2_fill_8 FILLER_0_151_208 ();
 sg13g2_fill_8 FILLER_0_151_216 ();
 sg13g2_fill_8 FILLER_0_151_224 ();
 sg13g2_fill_8 FILLER_0_151_232 ();
 sg13g2_fill_8 FILLER_0_151_240 ();
 sg13g2_fill_8 FILLER_0_151_248 ();
 sg13g2_fill_8 FILLER_0_151_256 ();
 sg13g2_fill_8 FILLER_0_151_264 ();
 sg13g2_fill_8 FILLER_0_151_272 ();
 sg13g2_fill_8 FILLER_0_151_280 ();
 sg13g2_fill_8 FILLER_0_151_288 ();
 sg13g2_fill_8 FILLER_0_151_296 ();
 sg13g2_fill_8 FILLER_0_151_304 ();
 sg13g2_fill_8 FILLER_0_151_312 ();
 sg13g2_fill_8 FILLER_0_151_320 ();
 sg13g2_fill_8 FILLER_0_151_328 ();
 sg13g2_fill_8 FILLER_0_151_336 ();
 sg13g2_fill_8 FILLER_0_151_344 ();
 sg13g2_fill_8 FILLER_0_151_352 ();
 sg13g2_fill_8 FILLER_0_151_360 ();
 sg13g2_fill_8 FILLER_0_151_368 ();
 sg13g2_fill_8 FILLER_0_151_376 ();
 sg13g2_fill_8 FILLER_0_151_384 ();
 sg13g2_fill_8 FILLER_0_151_392 ();
 sg13g2_fill_8 FILLER_0_151_400 ();
 sg13g2_fill_1 FILLER_0_151_408 ();
 sg13g2_fill_1 FILLER_0_151_435 ();
 sg13g2_fill_2 FILLER_0_151_441 ();
 sg13g2_fill_2 FILLER_0_151_453 ();
 sg13g2_fill_2 FILLER_0_151_460 ();
 sg13g2_fill_4 FILLER_0_151_472 ();
 sg13g2_fill_2 FILLER_0_151_476 ();
 sg13g2_fill_4 FILLER_0_151_518 ();
 sg13g2_fill_1 FILLER_0_151_526 ();
 sg13g2_fill_4 FILLER_0_151_553 ();
 sg13g2_fill_2 FILLER_0_151_562 ();
 sg13g2_fill_1 FILLER_0_151_564 ();
 sg13g2_fill_1 FILLER_0_151_617 ();
 sg13g2_fill_2 FILLER_0_151_633 ();
 sg13g2_fill_1 FILLER_0_151_635 ();
 sg13g2_fill_8 FILLER_0_151_662 ();
 sg13g2_decap_8 FILLER_0_151_670 ();
 sg13g2_fill_4 FILLER_0_151_703 ();
 sg13g2_fill_4 FILLER_0_151_712 ();
 sg13g2_fill_2 FILLER_0_151_716 ();
 sg13g2_fill_2 FILLER_0_151_758 ();
 sg13g2_fill_1 FILLER_0_151_760 ();
 sg13g2_fill_2 FILLER_0_151_789 ();
 sg13g2_fill_1 FILLER_0_151_791 ();
 sg13g2_fill_4 FILLER_0_151_802 ();
 sg13g2_fill_2 FILLER_0_151_837 ();
 sg13g2_fill_4 FILLER_0_151_849 ();
 sg13g2_fill_4 FILLER_0_151_903 ();
 sg13g2_fill_1 FILLER_0_151_907 ();
 sg13g2_fill_1 FILLER_0_151_934 ();
 sg13g2_fill_8 FILLER_0_151_939 ();
 sg13g2_fill_8 FILLER_0_151_947 ();
 sg13g2_fill_8 FILLER_0_151_955 ();
 sg13g2_fill_8 FILLER_0_151_963 ();
 sg13g2_fill_8 FILLER_0_151_971 ();
 sg13g2_fill_8 FILLER_0_151_979 ();
 sg13g2_fill_8 FILLER_0_151_987 ();
 sg13g2_fill_8 FILLER_0_151_995 ();
 sg13g2_fill_8 FILLER_0_151_1003 ();
 sg13g2_fill_8 FILLER_0_151_1011 ();
 sg13g2_fill_8 FILLER_0_151_1019 ();
 sg13g2_fill_8 FILLER_0_151_1027 ();
 sg13g2_fill_8 FILLER_0_151_1035 ();
 sg13g2_fill_8 FILLER_0_151_1043 ();
 sg13g2_fill_8 FILLER_0_151_1051 ();
 sg13g2_fill_8 FILLER_0_151_1059 ();
 sg13g2_fill_8 FILLER_0_151_1067 ();
 sg13g2_fill_8 FILLER_0_151_1075 ();
 sg13g2_fill_8 FILLER_0_151_1083 ();
 sg13g2_fill_8 FILLER_0_151_1091 ();
 sg13g2_fill_8 FILLER_0_151_1099 ();
 sg13g2_fill_8 FILLER_0_151_1107 ();
 sg13g2_fill_8 FILLER_0_151_1115 ();
 sg13g2_fill_8 FILLER_0_151_1123 ();
 sg13g2_fill_8 FILLER_0_151_1131 ();
 sg13g2_fill_8 FILLER_0_151_1139 ();
 sg13g2_fill_8 FILLER_0_151_1147 ();
 sg13g2_fill_8 FILLER_0_151_1155 ();
 sg13g2_fill_8 FILLER_0_151_1163 ();
 sg13g2_fill_8 FILLER_0_151_1171 ();
 sg13g2_fill_8 FILLER_0_151_1179 ();
 sg13g2_fill_8 FILLER_0_151_1187 ();
 sg13g2_fill_8 FILLER_0_151_1195 ();
 sg13g2_fill_8 FILLER_0_151_1203 ();
 sg13g2_fill_8 FILLER_0_151_1211 ();
 sg13g2_fill_8 FILLER_0_151_1219 ();
 sg13g2_fill_1 FILLER_0_151_1227 ();
 sg13g2_fill_8 FILLER_0_152_0 ();
 sg13g2_fill_8 FILLER_0_152_8 ();
 sg13g2_fill_8 FILLER_0_152_16 ();
 sg13g2_fill_8 FILLER_0_152_24 ();
 sg13g2_fill_8 FILLER_0_152_32 ();
 sg13g2_fill_8 FILLER_0_152_40 ();
 sg13g2_fill_8 FILLER_0_152_48 ();
 sg13g2_fill_8 FILLER_0_152_56 ();
 sg13g2_fill_8 FILLER_0_152_64 ();
 sg13g2_fill_8 FILLER_0_152_72 ();
 sg13g2_fill_8 FILLER_0_152_80 ();
 sg13g2_fill_8 FILLER_0_152_88 ();
 sg13g2_fill_8 FILLER_0_152_96 ();
 sg13g2_fill_8 FILLER_0_152_104 ();
 sg13g2_fill_8 FILLER_0_152_112 ();
 sg13g2_fill_8 FILLER_0_152_120 ();
 sg13g2_fill_8 FILLER_0_152_128 ();
 sg13g2_fill_8 FILLER_0_152_136 ();
 sg13g2_fill_8 FILLER_0_152_144 ();
 sg13g2_fill_8 FILLER_0_152_152 ();
 sg13g2_fill_8 FILLER_0_152_160 ();
 sg13g2_fill_8 FILLER_0_152_168 ();
 sg13g2_fill_8 FILLER_0_152_176 ();
 sg13g2_fill_8 FILLER_0_152_184 ();
 sg13g2_fill_8 FILLER_0_152_192 ();
 sg13g2_fill_8 FILLER_0_152_200 ();
 sg13g2_fill_8 FILLER_0_152_208 ();
 sg13g2_fill_8 FILLER_0_152_216 ();
 sg13g2_fill_8 FILLER_0_152_224 ();
 sg13g2_fill_8 FILLER_0_152_232 ();
 sg13g2_fill_8 FILLER_0_152_240 ();
 sg13g2_fill_8 FILLER_0_152_248 ();
 sg13g2_fill_8 FILLER_0_152_256 ();
 sg13g2_fill_8 FILLER_0_152_264 ();
 sg13g2_fill_8 FILLER_0_152_272 ();
 sg13g2_fill_8 FILLER_0_152_280 ();
 sg13g2_fill_8 FILLER_0_152_288 ();
 sg13g2_fill_8 FILLER_0_152_296 ();
 sg13g2_fill_8 FILLER_0_152_304 ();
 sg13g2_fill_8 FILLER_0_152_312 ();
 sg13g2_fill_8 FILLER_0_152_320 ();
 sg13g2_fill_8 FILLER_0_152_328 ();
 sg13g2_fill_8 FILLER_0_152_336 ();
 sg13g2_fill_8 FILLER_0_152_344 ();
 sg13g2_fill_8 FILLER_0_152_352 ();
 sg13g2_fill_8 FILLER_0_152_360 ();
 sg13g2_fill_8 FILLER_0_152_368 ();
 sg13g2_fill_8 FILLER_0_152_376 ();
 sg13g2_fill_8 FILLER_0_152_384 ();
 sg13g2_fill_8 FILLER_0_152_392 ();
 sg13g2_fill_8 FILLER_0_152_400 ();
 sg13g2_fill_1 FILLER_0_152_438 ();
 sg13g2_fill_1 FILLER_0_152_444 ();
 sg13g2_fill_1 FILLER_0_152_450 ();
 sg13g2_decap_8 FILLER_0_152_477 ();
 sg13g2_fill_1 FILLER_0_152_560 ();
 sg13g2_fill_2 FILLER_0_152_566 ();
 sg13g2_fill_8 FILLER_0_152_572 ();
 sg13g2_fill_1 FILLER_0_152_580 ();
 sg13g2_fill_1 FILLER_0_152_648 ();
 sg13g2_fill_8 FILLER_0_152_653 ();
 sg13g2_fill_8 FILLER_0_152_661 ();
 sg13g2_fill_4 FILLER_0_152_669 ();
 sg13g2_fill_8 FILLER_0_152_738 ();
 sg13g2_fill_4 FILLER_0_152_746 ();
 sg13g2_fill_2 FILLER_0_152_750 ();
 sg13g2_fill_1 FILLER_0_152_778 ();
 sg13g2_fill_2 FILLER_0_152_789 ();
 sg13g2_fill_1 FILLER_0_152_817 ();
 sg13g2_fill_2 FILLER_0_152_823 ();
 sg13g2_decap_8 FILLER_0_152_861 ();
 sg13g2_fill_1 FILLER_0_152_886 ();
 sg13g2_fill_2 FILLER_0_152_913 ();
 sg13g2_decap_8 FILLER_0_152_930 ();
 sg13g2_fill_8 FILLER_0_152_941 ();
 sg13g2_fill_8 FILLER_0_152_949 ();
 sg13g2_fill_8 FILLER_0_152_957 ();
 sg13g2_fill_8 FILLER_0_152_965 ();
 sg13g2_fill_8 FILLER_0_152_973 ();
 sg13g2_fill_8 FILLER_0_152_981 ();
 sg13g2_fill_8 FILLER_0_152_989 ();
 sg13g2_fill_8 FILLER_0_152_997 ();
 sg13g2_fill_8 FILLER_0_152_1005 ();
 sg13g2_fill_8 FILLER_0_152_1013 ();
 sg13g2_fill_8 FILLER_0_152_1021 ();
 sg13g2_fill_8 FILLER_0_152_1029 ();
 sg13g2_fill_8 FILLER_0_152_1037 ();
 sg13g2_fill_8 FILLER_0_152_1045 ();
 sg13g2_fill_8 FILLER_0_152_1053 ();
 sg13g2_fill_8 FILLER_0_152_1061 ();
 sg13g2_fill_8 FILLER_0_152_1069 ();
 sg13g2_fill_8 FILLER_0_152_1077 ();
 sg13g2_fill_8 FILLER_0_152_1085 ();
 sg13g2_fill_8 FILLER_0_152_1093 ();
 sg13g2_fill_8 FILLER_0_152_1101 ();
 sg13g2_fill_8 FILLER_0_152_1109 ();
 sg13g2_fill_8 FILLER_0_152_1117 ();
 sg13g2_fill_8 FILLER_0_152_1125 ();
 sg13g2_fill_8 FILLER_0_152_1133 ();
 sg13g2_fill_8 FILLER_0_152_1141 ();
 sg13g2_fill_8 FILLER_0_152_1149 ();
 sg13g2_fill_8 FILLER_0_152_1157 ();
 sg13g2_fill_8 FILLER_0_152_1165 ();
 sg13g2_fill_8 FILLER_0_152_1173 ();
 sg13g2_fill_8 FILLER_0_152_1181 ();
 sg13g2_fill_8 FILLER_0_152_1189 ();
 sg13g2_fill_8 FILLER_0_152_1197 ();
 sg13g2_fill_8 FILLER_0_152_1205 ();
 sg13g2_fill_8 FILLER_0_152_1213 ();
 sg13g2_decap_8 FILLER_0_152_1221 ();
 sg13g2_fill_8 FILLER_0_153_0 ();
 sg13g2_fill_8 FILLER_0_153_8 ();
 sg13g2_fill_8 FILLER_0_153_16 ();
 sg13g2_fill_8 FILLER_0_153_24 ();
 sg13g2_fill_8 FILLER_0_153_32 ();
 sg13g2_fill_8 FILLER_0_153_40 ();
 sg13g2_fill_8 FILLER_0_153_48 ();
 sg13g2_fill_8 FILLER_0_153_56 ();
 sg13g2_fill_8 FILLER_0_153_64 ();
 sg13g2_fill_8 FILLER_0_153_72 ();
 sg13g2_fill_8 FILLER_0_153_80 ();
 sg13g2_fill_8 FILLER_0_153_88 ();
 sg13g2_fill_8 FILLER_0_153_96 ();
 sg13g2_fill_8 FILLER_0_153_104 ();
 sg13g2_fill_8 FILLER_0_153_112 ();
 sg13g2_fill_8 FILLER_0_153_120 ();
 sg13g2_fill_8 FILLER_0_153_128 ();
 sg13g2_fill_8 FILLER_0_153_136 ();
 sg13g2_fill_8 FILLER_0_153_144 ();
 sg13g2_fill_8 FILLER_0_153_152 ();
 sg13g2_fill_8 FILLER_0_153_160 ();
 sg13g2_fill_8 FILLER_0_153_168 ();
 sg13g2_fill_8 FILLER_0_153_176 ();
 sg13g2_fill_8 FILLER_0_153_184 ();
 sg13g2_fill_8 FILLER_0_153_192 ();
 sg13g2_fill_8 FILLER_0_153_200 ();
 sg13g2_fill_8 FILLER_0_153_208 ();
 sg13g2_fill_8 FILLER_0_153_216 ();
 sg13g2_fill_8 FILLER_0_153_224 ();
 sg13g2_fill_8 FILLER_0_153_232 ();
 sg13g2_fill_8 FILLER_0_153_240 ();
 sg13g2_fill_8 FILLER_0_153_248 ();
 sg13g2_fill_8 FILLER_0_153_256 ();
 sg13g2_fill_8 FILLER_0_153_264 ();
 sg13g2_fill_8 FILLER_0_153_272 ();
 sg13g2_fill_8 FILLER_0_153_280 ();
 sg13g2_fill_8 FILLER_0_153_288 ();
 sg13g2_fill_8 FILLER_0_153_296 ();
 sg13g2_fill_8 FILLER_0_153_304 ();
 sg13g2_fill_8 FILLER_0_153_312 ();
 sg13g2_fill_8 FILLER_0_153_320 ();
 sg13g2_fill_8 FILLER_0_153_328 ();
 sg13g2_fill_8 FILLER_0_153_336 ();
 sg13g2_fill_8 FILLER_0_153_344 ();
 sg13g2_fill_8 FILLER_0_153_352 ();
 sg13g2_fill_8 FILLER_0_153_360 ();
 sg13g2_fill_8 FILLER_0_153_368 ();
 sg13g2_fill_8 FILLER_0_153_376 ();
 sg13g2_fill_8 FILLER_0_153_384 ();
 sg13g2_fill_8 FILLER_0_153_392 ();
 sg13g2_fill_8 FILLER_0_153_400 ();
 sg13g2_fill_8 FILLER_0_153_408 ();
 sg13g2_fill_4 FILLER_0_153_416 ();
 sg13g2_fill_2 FILLER_0_153_420 ();
 sg13g2_fill_8 FILLER_0_153_436 ();
 sg13g2_fill_4 FILLER_0_153_478 ();
 sg13g2_fill_4 FILLER_0_153_486 ();
 sg13g2_fill_1 FILLER_0_153_490 ();
 sg13g2_fill_2 FILLER_0_153_500 ();
 sg13g2_fill_4 FILLER_0_153_533 ();
 sg13g2_fill_2 FILLER_0_153_537 ();
 sg13g2_fill_8 FILLER_0_153_583 ();
 sg13g2_fill_2 FILLER_0_153_595 ();
 sg13g2_fill_2 FILLER_0_153_617 ();
 sg13g2_fill_8 FILLER_0_153_649 ();
 sg13g2_fill_8 FILLER_0_153_657 ();
 sg13g2_fill_8 FILLER_0_153_665 ();
 sg13g2_fill_8 FILLER_0_153_673 ();
 sg13g2_fill_2 FILLER_0_153_681 ();
 sg13g2_decap_8 FILLER_0_153_687 ();
 sg13g2_fill_1 FILLER_0_153_699 ();
 sg13g2_fill_2 FILLER_0_153_710 ();
 sg13g2_fill_8 FILLER_0_153_726 ();
 sg13g2_fill_8 FILLER_0_153_734 ();
 sg13g2_fill_8 FILLER_0_153_742 ();
 sg13g2_fill_8 FILLER_0_153_750 ();
 sg13g2_fill_2 FILLER_0_153_766 ();
 sg13g2_fill_4 FILLER_0_153_783 ();
 sg13g2_decap_8 FILLER_0_153_792 ();
 sg13g2_decap_8 FILLER_0_153_803 ();
 sg13g2_fill_2 FILLER_0_153_845 ();
 sg13g2_fill_1 FILLER_0_153_847 ();
 sg13g2_fill_8 FILLER_0_153_917 ();
 sg13g2_fill_2 FILLER_0_153_925 ();
 sg13g2_fill_1 FILLER_0_153_927 ();
 sg13g2_fill_8 FILLER_0_153_954 ();
 sg13g2_fill_8 FILLER_0_153_962 ();
 sg13g2_fill_8 FILLER_0_153_970 ();
 sg13g2_fill_8 FILLER_0_153_978 ();
 sg13g2_fill_8 FILLER_0_153_986 ();
 sg13g2_fill_8 FILLER_0_153_994 ();
 sg13g2_fill_8 FILLER_0_153_1002 ();
 sg13g2_fill_8 FILLER_0_153_1010 ();
 sg13g2_fill_8 FILLER_0_153_1018 ();
 sg13g2_fill_8 FILLER_0_153_1026 ();
 sg13g2_fill_8 FILLER_0_153_1034 ();
 sg13g2_fill_8 FILLER_0_153_1042 ();
 sg13g2_fill_8 FILLER_0_153_1050 ();
 sg13g2_fill_8 FILLER_0_153_1058 ();
 sg13g2_fill_8 FILLER_0_153_1066 ();
 sg13g2_fill_8 FILLER_0_153_1074 ();
 sg13g2_fill_8 FILLER_0_153_1082 ();
 sg13g2_fill_8 FILLER_0_153_1090 ();
 sg13g2_fill_8 FILLER_0_153_1098 ();
 sg13g2_fill_8 FILLER_0_153_1106 ();
 sg13g2_fill_8 FILLER_0_153_1114 ();
 sg13g2_fill_8 FILLER_0_153_1122 ();
 sg13g2_fill_8 FILLER_0_153_1130 ();
 sg13g2_fill_8 FILLER_0_153_1138 ();
 sg13g2_fill_8 FILLER_0_153_1146 ();
 sg13g2_fill_8 FILLER_0_153_1154 ();
 sg13g2_fill_8 FILLER_0_153_1162 ();
 sg13g2_fill_8 FILLER_0_153_1170 ();
 sg13g2_fill_8 FILLER_0_153_1178 ();
 sg13g2_fill_8 FILLER_0_153_1186 ();
 sg13g2_fill_8 FILLER_0_153_1194 ();
 sg13g2_fill_8 FILLER_0_153_1202 ();
 sg13g2_fill_8 FILLER_0_153_1210 ();
 sg13g2_fill_8 FILLER_0_153_1218 ();
 sg13g2_fill_2 FILLER_0_153_1226 ();
 sg13g2_fill_8 FILLER_0_154_0 ();
 sg13g2_fill_8 FILLER_0_154_8 ();
 sg13g2_fill_8 FILLER_0_154_16 ();
 sg13g2_fill_8 FILLER_0_154_24 ();
 sg13g2_fill_8 FILLER_0_154_32 ();
 sg13g2_fill_8 FILLER_0_154_40 ();
 sg13g2_fill_8 FILLER_0_154_48 ();
 sg13g2_fill_8 FILLER_0_154_56 ();
 sg13g2_fill_8 FILLER_0_154_64 ();
 sg13g2_fill_8 FILLER_0_154_72 ();
 sg13g2_fill_8 FILLER_0_154_80 ();
 sg13g2_fill_8 FILLER_0_154_88 ();
 sg13g2_fill_8 FILLER_0_154_96 ();
 sg13g2_fill_8 FILLER_0_154_104 ();
 sg13g2_fill_8 FILLER_0_154_112 ();
 sg13g2_fill_8 FILLER_0_154_120 ();
 sg13g2_fill_8 FILLER_0_154_128 ();
 sg13g2_fill_8 FILLER_0_154_136 ();
 sg13g2_fill_8 FILLER_0_154_144 ();
 sg13g2_fill_8 FILLER_0_154_152 ();
 sg13g2_fill_8 FILLER_0_154_160 ();
 sg13g2_fill_8 FILLER_0_154_168 ();
 sg13g2_fill_8 FILLER_0_154_176 ();
 sg13g2_fill_8 FILLER_0_154_184 ();
 sg13g2_fill_8 FILLER_0_154_192 ();
 sg13g2_fill_8 FILLER_0_154_200 ();
 sg13g2_fill_8 FILLER_0_154_208 ();
 sg13g2_fill_8 FILLER_0_154_216 ();
 sg13g2_fill_8 FILLER_0_154_224 ();
 sg13g2_fill_8 FILLER_0_154_232 ();
 sg13g2_fill_8 FILLER_0_154_240 ();
 sg13g2_fill_8 FILLER_0_154_248 ();
 sg13g2_fill_8 FILLER_0_154_256 ();
 sg13g2_fill_8 FILLER_0_154_264 ();
 sg13g2_fill_8 FILLER_0_154_272 ();
 sg13g2_fill_8 FILLER_0_154_280 ();
 sg13g2_fill_8 FILLER_0_154_288 ();
 sg13g2_fill_8 FILLER_0_154_296 ();
 sg13g2_fill_8 FILLER_0_154_304 ();
 sg13g2_fill_8 FILLER_0_154_312 ();
 sg13g2_fill_8 FILLER_0_154_320 ();
 sg13g2_fill_8 FILLER_0_154_328 ();
 sg13g2_fill_8 FILLER_0_154_336 ();
 sg13g2_fill_8 FILLER_0_154_344 ();
 sg13g2_fill_8 FILLER_0_154_352 ();
 sg13g2_fill_8 FILLER_0_154_360 ();
 sg13g2_fill_8 FILLER_0_154_368 ();
 sg13g2_fill_8 FILLER_0_154_376 ();
 sg13g2_fill_8 FILLER_0_154_384 ();
 sg13g2_fill_8 FILLER_0_154_392 ();
 sg13g2_fill_8 FILLER_0_154_400 ();
 sg13g2_fill_8 FILLER_0_154_408 ();
 sg13g2_fill_8 FILLER_0_154_416 ();
 sg13g2_fill_8 FILLER_0_154_424 ();
 sg13g2_fill_8 FILLER_0_154_432 ();
 sg13g2_fill_8 FILLER_0_154_440 ();
 sg13g2_fill_2 FILLER_0_154_448 ();
 sg13g2_fill_4 FILLER_0_154_454 ();
 sg13g2_fill_1 FILLER_0_154_458 ();
 sg13g2_fill_8 FILLER_0_154_463 ();
 sg13g2_fill_2 FILLER_0_154_471 ();
 sg13g2_fill_1 FILLER_0_154_473 ();
 sg13g2_fill_8 FILLER_0_154_500 ();
 sg13g2_fill_8 FILLER_0_154_508 ();
 sg13g2_fill_8 FILLER_0_154_521 ();
 sg13g2_fill_8 FILLER_0_154_529 ();
 sg13g2_fill_4 FILLER_0_154_537 ();
 sg13g2_fill_1 FILLER_0_154_541 ();
 sg13g2_fill_8 FILLER_0_154_568 ();
 sg13g2_fill_8 FILLER_0_154_576 ();
 sg13g2_fill_8 FILLER_0_154_584 ();
 sg13g2_fill_8 FILLER_0_154_592 ();
 sg13g2_fill_8 FILLER_0_154_600 ();
 sg13g2_fill_8 FILLER_0_154_608 ();
 sg13g2_fill_8 FILLER_0_154_616 ();
 sg13g2_fill_4 FILLER_0_154_624 ();
 sg13g2_fill_2 FILLER_0_154_628 ();
 sg13g2_fill_8 FILLER_0_154_634 ();
 sg13g2_fill_8 FILLER_0_154_642 ();
 sg13g2_fill_8 FILLER_0_154_650 ();
 sg13g2_fill_8 FILLER_0_154_658 ();
 sg13g2_fill_8 FILLER_0_154_666 ();
 sg13g2_fill_8 FILLER_0_154_674 ();
 sg13g2_fill_8 FILLER_0_154_682 ();
 sg13g2_fill_8 FILLER_0_154_690 ();
 sg13g2_fill_8 FILLER_0_154_698 ();
 sg13g2_fill_8 FILLER_0_154_706 ();
 sg13g2_fill_8 FILLER_0_154_714 ();
 sg13g2_fill_8 FILLER_0_154_722 ();
 sg13g2_fill_8 FILLER_0_154_730 ();
 sg13g2_fill_8 FILLER_0_154_738 ();
 sg13g2_fill_8 FILLER_0_154_746 ();
 sg13g2_fill_8 FILLER_0_154_780 ();
 sg13g2_fill_8 FILLER_0_154_788 ();
 sg13g2_fill_8 FILLER_0_154_796 ();
 sg13g2_fill_8 FILLER_0_154_804 ();
 sg13g2_fill_4 FILLER_0_154_812 ();
 sg13g2_fill_1 FILLER_0_154_816 ();
 sg13g2_fill_8 FILLER_0_154_821 ();
 sg13g2_fill_8 FILLER_0_154_829 ();
 sg13g2_fill_8 FILLER_0_154_837 ();
 sg13g2_fill_8 FILLER_0_154_845 ();
 sg13g2_fill_4 FILLER_0_154_853 ();
 sg13g2_fill_1 FILLER_0_154_857 ();
 sg13g2_fill_8 FILLER_0_154_862 ();
 sg13g2_fill_8 FILLER_0_154_870 ();
 sg13g2_fill_4 FILLER_0_154_878 ();
 sg13g2_fill_8 FILLER_0_154_887 ();
 sg13g2_fill_8 FILLER_0_154_895 ();
 sg13g2_fill_8 FILLER_0_154_903 ();
 sg13g2_fill_8 FILLER_0_154_911 ();
 sg13g2_fill_8 FILLER_0_154_919 ();
 sg13g2_fill_8 FILLER_0_154_927 ();
 sg13g2_fill_8 FILLER_0_154_935 ();
 sg13g2_fill_8 FILLER_0_154_943 ();
 sg13g2_fill_8 FILLER_0_154_951 ();
 sg13g2_fill_8 FILLER_0_154_959 ();
 sg13g2_fill_8 FILLER_0_154_967 ();
 sg13g2_fill_8 FILLER_0_154_975 ();
 sg13g2_fill_8 FILLER_0_154_983 ();
 sg13g2_fill_8 FILLER_0_154_991 ();
 sg13g2_fill_8 FILLER_0_154_999 ();
 sg13g2_fill_8 FILLER_0_154_1007 ();
 sg13g2_fill_8 FILLER_0_154_1015 ();
 sg13g2_fill_8 FILLER_0_154_1023 ();
 sg13g2_fill_8 FILLER_0_154_1031 ();
 sg13g2_fill_8 FILLER_0_154_1039 ();
 sg13g2_fill_8 FILLER_0_154_1047 ();
 sg13g2_fill_8 FILLER_0_154_1055 ();
 sg13g2_fill_8 FILLER_0_154_1063 ();
 sg13g2_fill_8 FILLER_0_154_1071 ();
 sg13g2_fill_8 FILLER_0_154_1079 ();
 sg13g2_fill_8 FILLER_0_154_1087 ();
 sg13g2_fill_8 FILLER_0_154_1095 ();
 sg13g2_fill_8 FILLER_0_154_1103 ();
 sg13g2_fill_8 FILLER_0_154_1111 ();
 sg13g2_fill_8 FILLER_0_154_1119 ();
 sg13g2_fill_8 FILLER_0_154_1127 ();
 sg13g2_fill_8 FILLER_0_154_1135 ();
 sg13g2_fill_8 FILLER_0_154_1143 ();
 sg13g2_fill_8 FILLER_0_154_1151 ();
 sg13g2_fill_8 FILLER_0_154_1159 ();
 sg13g2_fill_8 FILLER_0_154_1167 ();
 sg13g2_fill_8 FILLER_0_154_1175 ();
 sg13g2_fill_8 FILLER_0_154_1183 ();
 sg13g2_fill_8 FILLER_0_154_1191 ();
 sg13g2_fill_8 FILLER_0_154_1199 ();
 sg13g2_fill_8 FILLER_0_154_1207 ();
 sg13g2_fill_8 FILLER_0_154_1215 ();
 sg13g2_fill_4 FILLER_0_154_1223 ();
 sg13g2_fill_1 FILLER_0_154_1227 ();
endmodule
