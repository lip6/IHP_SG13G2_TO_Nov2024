module martin_top (aux_enable_pad,
    clk_pad,
    lfsr_out_pad,
    rst_pad,
    shreg_in_pad,
    shreg_out_pad,
    wr_enable_pad,
    data_in_pad,
    data_out_pad,
    out_select_pad,
    reg_addr_pad);
 inout aux_enable_pad;
 inout clk_pad;
 inout lfsr_out_pad;
 inout rst_pad;
 inout shreg_in_pad;
 inout shreg_out_pad;
 inout wr_enable_pad;
 inout [7:0] data_in_pad;
 inout [7:0] data_out_pad;
 inout [1:0] out_select_pad;
 inout [2:0] reg_addr_pad;

 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire net606;
 wire net605;
 wire net604;
 wire net603;
 wire _01707_;
 wire net602;
 wire _01709_;
 wire _01710_;
 wire net601;
 wire _01712_;
 wire net600;
 wire net599;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire net598;
 wire _01719_;
 wire net597;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire net596;
 wire _01725_;
 wire _01726_;
 wire net595;
 wire net594;
 wire net593;
 wire _01730_;
 wire net592;
 wire net591;
 wire _01733_;
 wire net590;
 wire net589;
 wire _01736_;
 wire net588;
 wire net587;
 wire net586;
 wire net585;
 wire _01741_;
 wire net584;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire net583;
 wire net582;
 wire net581;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire net580;
 wire net579;
 wire net578;
 wire _01765_;
 wire _01766_;
 wire net577;
 wire net576;
 wire net575;
 wire _01770_;
 wire _01771_;
 wire net574;
 wire _01773_;
 wire net573;
 wire net572;
 wire _01776_;
 wire _01777_;
 wire net571;
 wire net570;
 wire _01780_;
 wire _01781_;
 wire net569;
 wire _01783_;
 wire net568;
 wire net567;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire net566;
 wire _01790_;
 wire _01791_;
 wire net565;
 wire net564;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire net563;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire net562;
 wire _01804_;
 wire net561;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire net560;
 wire net559;
 wire _01814_;
 wire net558;
 wire net557;
 wire net556;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire net555;
 wire _01822_;
 wire net554;
 wire _01824_;
 wire net553;
 wire net552;
 wire net551;
 wire _01828_;
 wire _01829_;
 wire net550;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire net549;
 wire _01835_;
 wire _01836_;
 wire net548;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire net547;
 wire _01842_;
 wire _01843_;
 wire net546;
 wire net545;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire net544;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire net543;
 wire _01861_;
 wire net542;
 wire _01863_;
 wire _01864_;
 wire net541;
 wire net540;
 wire net539;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire net538;
 wire _01873_;
 wire _01874_;
 wire net537;
 wire net536;
 wire _01877_;
 wire _01878_;
 wire net535;
 wire net534;
 wire _01881_;
 wire net533;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire net532;
 wire net531;
 wire net530;
 wire net529;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire net528;
 wire _01901_;
 wire net527;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire net526;
 wire net525;
 wire net524;
 wire net523;
 wire _01918_;
 wire net522;
 wire _01920_;
 wire net521;
 wire _01922_;
 wire _01923_;
 wire net520;
 wire net519;
 wire _01926_;
 wire _01927_;
 wire net518;
 wire net517;
 wire _01930_;
 wire _01931_;
 wire net516;
 wire net515;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire net514;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire net513;
 wire _01945_;
 wire net512;
 wire net511;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire net510;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire net509;
 wire net508;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire net507;
 wire net506;
 wire net505;
 wire net504;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire net503;
 wire _01985_;
 wire _01986_;
 wire net502;
 wire net501;
 wire _01989_;
 wire net500;
 wire _01991_;
 wire _01992_;
 wire net499;
 wire net498;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire net497;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire net496;
 wire _02006_;
 wire net495;
 wire net494;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire net493;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire net492;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire net491;
 wire net490;
 wire net489;
 wire net488;
 wire net487;
 wire net486;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire net485;
 wire _02033_;
 wire net484;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire net483;
 wire net482;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire net481;
 wire net480;
 wire net479;
 wire net478;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire net477;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire net476;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire net475;
 wire net474;
 wire net473;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire net472;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire net471;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire net470;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire net469;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire net468;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire net467;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire net466;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire net465;
 wire _02260_;
 wire _02261_;
 wire net464;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire net463;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire net462;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire net461;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire net460;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire net459;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire net458;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire net457;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire net456;
 wire net455;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire net454;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire net453;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire net452;
 wire _02463_;
 wire net451;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire net450;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire net449;
 wire net448;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire net447;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire net446;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire net445;
 wire _02604_;
 wire net444;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire net443;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire net442;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire net441;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire net440;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire net439;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire net438;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire net437;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire net436;
 wire _02750_;
 wire net435;
 wire _02752_;
 wire net434;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire net433;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire net432;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire net431;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire net430;
 wire _02828_;
 wire _02829_;
 wire net429;
 wire _02831_;
 wire _02832_;
 wire net428;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire net427;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire net426;
 wire _02888_;
 wire _02889_;
 wire net425;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire net424;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire net423;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire net422;
 wire net421;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire net420;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire net419;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire net418;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire net417;
 wire net416;
 wire net415;
 wire net414;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire net413;
 wire net412;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire net411;
 wire net410;
 wire net409;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire net408;
 wire net407;
 wire net406;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire net405;
 wire net404;
 wire _03061_;
 wire net403;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire net402;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire net401;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire net400;
 wire net399;
 wire _03078_;
 wire _03079_;
 wire net398;
 wire net397;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire net396;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire net395;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire net394;
 wire _03117_;
 wire _03118_;
 wire net393;
 wire net392;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire net391;
 wire net390;
 wire _03140_;
 wire net389;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire net388;
 wire net387;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire net386;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire net385;
 wire net384;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire net383;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire net382;
 wire net381;
 wire _03207_;
 wire net380;
 wire net379;
 wire _03210_;
 wire net378;
 wire net377;
 wire net376;
 wire net375;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire net374;
 wire net373;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire net372;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire net371;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire net370;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire net369;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire net368;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire net367;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire net366;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire net365;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire net364;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire net363;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire net362;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire net361;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire net360;
 wire net359;
 wire net358;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire net357;
 wire net356;
 wire net355;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire net354;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire net353;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire net352;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire net351;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire net350;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire net349;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire net348;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire net347;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire net346;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire net345;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire net344;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire net343;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire net342;
 wire net341;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire net340;
 wire net339;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire net338;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire net337;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire net336;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire net335;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire net334;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire net333;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire net332;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire net331;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire net330;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire net329;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire net328;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire net327;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire net326;
 wire net325;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire net324;
 wire net323;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire net322;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire net321;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire net320;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire net319;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire net318;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire net317;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire net316;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire net315;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire net314;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire net313;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire net312;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire net311;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire net310;
 wire net309;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire net308;
 wire net307;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire net306;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire net305;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire net304;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire net303;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire net302;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire net301;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire net300;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire net299;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire net298;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire net297;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire net296;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire net295;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire net294;
 wire net293;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire net292;
 wire net291;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire net290;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire net289;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire net288;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire net287;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire net286;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire net285;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire net284;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire net283;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire net282;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire net281;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire net280;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire net279;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire net278;
 wire net277;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire net276;
 wire net275;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire net274;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire net273;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire net272;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire net271;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire net270;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire net269;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire net268;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire net267;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire net266;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire net265;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire net264;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire net263;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire net262;
 wire net261;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire net260;
 wire net259;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire net258;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire net257;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire net256;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire net255;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire net254;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire net253;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire net252;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire net251;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire net250;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire net249;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire net248;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire net247;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire net246;
 wire net245;
 wire net244;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire net243;
 wire net242;
 wire net241;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire net240;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire net239;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire net238;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire net237;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire net236;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire net235;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire net234;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire net233;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire net232;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire net231;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire net230;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire net229;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire net228;
 wire net227;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire net226;
 wire net225;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire net224;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire net223;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire net222;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire net221;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire net220;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire net219;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire net218;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire net217;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire net216;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire net215;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire net214;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire net213;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire net212;
 wire net211;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire net210;
 wire net209;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire net208;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire net207;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire net206;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire net205;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire net204;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire net203;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire net202;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire net201;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire net200;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire net199;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire net198;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire net197;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire net196;
 wire net195;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire net194;
 wire net193;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire net192;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire net191;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire net190;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire net189;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire net188;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire net187;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire net186;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire net185;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire net184;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire net183;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire net182;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire net181;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire net180;
 wire net179;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire net178;
 wire net177;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire net176;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire net175;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire net174;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire net173;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire net172;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire net171;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire net170;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire net169;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire net168;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire net167;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire net166;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire net165;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire net164;
 wire net163;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire net162;
 wire net161;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire net160;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire net159;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire net158;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire net157;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire net156;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire net155;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire net154;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire net153;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire net152;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire net151;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire net150;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire net149;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire net148;
 wire net147;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire net146;
 wire net145;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire net144;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire net143;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire net142;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire net141;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire net140;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire net139;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire net138;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire net137;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire net136;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire net135;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire net134;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire net133;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire net132;
 wire net131;
 wire net130;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire net129;
 wire net128;
 wire net127;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire net126;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire net125;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire net124;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire net123;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire net122;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire net121;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire net120;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire net119;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire net118;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire net117;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire net116;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire net115;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire net114;
 wire net113;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire net112;
 wire net111;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire net110;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire net109;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire net108;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire net107;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire net106;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire net105;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire net104;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire net103;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire net102;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire net101;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire net100;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire net99;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire net98;
 wire net97;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire net96;
 wire net95;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire net94;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire net93;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire net92;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire net91;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire net90;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire net89;
 wire _04724_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire net88;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire net87;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire net86;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire net85;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire net84;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire net83;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire net82;
 wire net81;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire net80;
 wire net79;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire net78;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire net77;
 wire _04786_;
 wire _04787_;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire net76;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire net75;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire net74;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire net73;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire net72;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire net71;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire net70;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire net69;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire net68;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire net67;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire net66;
 wire net65;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire net64;
 wire net63;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire net62;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire net61;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire net60;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire net59;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire net58;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire net57;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire net56;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire net55;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire net54;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire net53;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire net52;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire net51;
 wire _04932_;
 wire _04933_;
 wire _04934_;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire net50;
 wire net49;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire net48;
 wire net47;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire _04952_;
 wire net46;
 wire _04954_;
 wire _04955_;
 wire _04956_;
 wire net45;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire net44;
 wire _04966_;
 wire _04967_;
 wire _04968_;
 wire net43;
 wire _04970_;
 wire _04971_;
 wire _04972_;
 wire _04973_;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire net42;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire net41;
 wire _04982_;
 wire _04983_;
 wire _04984_;
 wire _04985_;
 wire _04986_;
 wire _04987_;
 wire _04988_;
 wire net40;
 wire _04990_;
 wire _04991_;
 wire _04992_;
 wire net39;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04997_;
 wire _04998_;
 wire _04999_;
 wire _05000_;
 wire net38;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire net37;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire _05012_;
 wire net34;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire net36;
 wire _05018_;
 wire _05019_;
 wire _05020_;
 wire _05021_;
 wire _05022_;
 wire _05023_;
 wire _05024_;
 wire net35;
 wire net33;
 wire _05027_;
 wire _05028_;
 wire _05029_;
 wire net4050;
 wire net31;
 wire _05032_;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire _05036_;
 wire _05037_;
 wire _05038_;
 wire net30;
 wire _05040_;
 wire _05041_;
 wire _05042_;
 wire net29;
 wire _05044_;
 wire _05045_;
 wire _05046_;
 wire _05047_;
 wire _05048_;
 wire _05049_;
 wire _05050_;
 wire net28;
 wire _05052_;
 wire _05053_;
 wire _05054_;
 wire net27;
 wire _05056_;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire _05061_;
 wire _05062_;
 wire net26;
 wire _05064_;
 wire _05065_;
 wire _05066_;
 wire net25;
 wire _05068_;
 wire _05069_;
 wire _05070_;
 wire _05071_;
 wire _05072_;
 wire _05073_;
 wire _05074_;
 wire net24;
 wire _05076_;
 wire _05077_;
 wire _05078_;
 wire net23;
 wire _05080_;
 wire _05081_;
 wire _05082_;
 wire _05083_;
 wire _05084_;
 wire _05085_;
 wire _05086_;
 wire net21;
 wire _05088_;
 wire _05089_;
 wire _05090_;
 wire net4037;
 wire _05092_;
 wire _05093_;
 wire _05094_;
 wire _05095_;
 wire _05096_;
 wire _05097_;
 wire _05098_;
 wire net20;
 wire _05100_;
 wire _05101_;
 wire _05102_;
 wire net19;
 wire _05104_;
 wire _05105_;
 wire _05106_;
 wire _05107_;
 wire _05108_;
 wire _05109_;
 wire _05110_;
 wire net18;
 wire _05112_;
 wire _05113_;
 wire _05114_;
 wire net16;
 wire _05116_;
 wire _05117_;
 wire _05118_;
 wire _05119_;
 wire _05120_;
 wire _05121_;
 wire _05122_;
 wire net15;
 wire _05124_;
 wire _05125_;
 wire _05126_;
 wire net4031;
 wire _05128_;
 wire _05129_;
 wire _05130_;
 wire _05131_;
 wire _05132_;
 wire _05133_;
 wire _05134_;
 wire net14;
 wire _05136_;
 wire _05137_;
 wire _05138_;
 wire net13;
 wire _05140_;
 wire _05141_;
 wire _05142_;
 wire _05143_;
 wire _05144_;
 wire _05145_;
 wire _05146_;
 wire net12;
 wire _05148_;
 wire _05149_;
 wire _05150_;
 wire net11;
 wire _05152_;
 wire _05153_;
 wire _05154_;
 wire _05155_;
 wire _05156_;
 wire _05157_;
 wire _05158_;
 wire net10;
 wire _05160_;
 wire _05161_;
 wire _05162_;
 wire net9;
 wire _05164_;
 wire _05165_;
 wire _05166_;
 wire _05167_;
 wire _05168_;
 wire _05169_;
 wire _05170_;
 wire net7;
 wire _05172_;
 wire _05173_;
 wire _05174_;
 wire _05175_;
 wire _05176_;
 wire _05177_;
 wire _05178_;
 wire _05179_;
 wire _05180_;
 wire _05181_;
 wire net4023;
 wire _05183_;
 wire net6;
 wire _05185_;
 wire net5;
 wire net4;
 wire net3;
 wire _05189_;
 wire _05190_;
 wire _05191_;
 wire _05192_;
 wire _05193_;
 wire _05194_;
 wire _05195_;
 wire _05196_;
 wire _05197_;
 wire _05198_;
 wire _05199_;
 wire _05200_;
 wire _05201_;
 wire _05202_;
 wire net2;
 wire _05204_;
 wire _05205_;
 wire _05206_;
 wire _05207_;
 wire _05208_;
 wire _05209_;
 wire _05210_;
 wire _05211_;
 wire _05212_;
 wire _05213_;
 wire _05214_;
 wire net1;
 wire _05216_;
 wire _05217_;
 wire _05218_;
 wire _05219_;
 wire _05220_;
 wire _05221_;
 wire _05222_;
 wire _05223_;
 wire _05224_;
 wire _05225_;
 wire _05227_;
 wire _05228_;
 wire _05229_;
 wire _05230_;
 wire _05231_;
 wire _05232_;
 wire _05233_;
 wire _05234_;
 wire _05235_;
 wire _05236_;
 wire _05238_;
 wire _05239_;
 wire _05240_;
 wire _05241_;
 wire _05242_;
 wire _05243_;
 wire _05244_;
 wire _05245_;
 wire _05246_;
 wire _05247_;
 wire _05248_;
 wire _05249_;
 wire _05250_;
 wire _05251_;
 wire _05252_;
 wire _05253_;
 wire _05254_;
 wire _05255_;
 wire _05256_;
 wire _05257_;
 wire _05258_;
 wire _05259_;
 wire _05260_;
 wire _05261_;
 wire _05262_;
 wire _05263_;
 wire _05264_;
 wire _05265_;
 wire _05266_;
 wire _05267_;
 wire _05268_;
 wire _05269_;
 wire _05270_;
 wire _05271_;
 wire _05272_;
 wire _05273_;
 wire _05274_;
 wire _05275_;
 wire _05276_;
 wire _05277_;
 wire _05278_;
 wire _05279_;
 wire _05280_;
 wire _05281_;
 wire _05282_;
 wire _05283_;
 wire _05284_;
 wire _05285_;
 wire _05286_;
 wire _05287_;
 wire _05288_;
 wire _05289_;
 wire _05290_;
 wire _05291_;
 wire _05292_;
 wire _05293_;
 wire _05294_;
 wire _05295_;
 wire _05296_;
 wire _05297_;
 wire _05298_;
 wire _05299_;
 wire _05300_;
 wire _05301_;
 wire _05302_;
 wire _05303_;
 wire _05304_;
 wire _05305_;
 wire _05306_;
 wire _05307_;
 wire _05308_;
 wire _05309_;
 wire _05310_;
 wire _05311_;
 wire _05312_;
 wire _05313_;
 wire _05314_;
 wire _05315_;
 wire _05316_;
 wire _05317_;
 wire _05318_;
 wire _05319_;
 wire _05320_;
 wire _05321_;
 wire _05322_;
 wire _05323_;
 wire _05324_;
 wire _05325_;
 wire _05326_;
 wire _05327_;
 wire _05328_;
 wire _05329_;
 wire _05330_;
 wire _05331_;
 wire _05332_;
 wire _05333_;
 wire _05334_;
 wire _05335_;
 wire _05336_;
 wire _05337_;
 wire _05338_;
 wire _05339_;
 wire _05340_;
 wire _05341_;
 wire _05342_;
 wire _05343_;
 wire _05344_;
 wire _05345_;
 wire _05346_;
 wire _05347_;
 wire _05348_;
 wire _05349_;
 wire _05350_;
 wire _05351_;
 wire _05352_;
 wire _05353_;
 wire _05354_;
 wire _05355_;
 wire _05356_;
 wire _05357_;
 wire _05358_;
 wire _05359_;
 wire _05360_;
 wire _05361_;
 wire _05362_;
 wire _05363_;
 wire _05364_;
 wire _05365_;
 wire _05366_;
 wire _05367_;
 wire _05368_;
 wire _05369_;
 wire _05370_;
 wire _05371_;
 wire _05372_;
 wire _05373_;
 wire _05374_;
 wire _05375_;
 wire _05376_;
 wire _05377_;
 wire _05378_;
 wire _05379_;
 wire _05380_;
 wire _05381_;
 wire _05382_;
 wire _05383_;
 wire _05384_;
 wire _05385_;
 wire _05386_;
 wire _05387_;
 wire _05388_;
 wire _05389_;
 wire _05390_;
 wire _05391_;
 wire _05392_;
 wire _05393_;
 wire _05394_;
 wire _05395_;
 wire _05396_;
 wire _05397_;
 wire _05398_;
 wire _05399_;
 wire _05400_;
 wire _05401_;
 wire _05402_;
 wire _05403_;
 wire _05404_;
 wire _05405_;
 wire _05406_;
 wire _05407_;
 wire _05408_;
 wire _05409_;
 wire _05410_;
 wire _05411_;
 wire _05412_;
 wire _05413_;
 wire _05414_;
 wire _05415_;
 wire _05416_;
 wire _05417_;
 wire _05418_;
 wire _05419_;
 wire _05420_;
 wire _05421_;
 wire _05422_;
 wire _05423_;
 wire _05424_;
 wire _05425_;
 wire _05426_;
 wire _05427_;
 wire _05428_;
 wire _05429_;
 wire _05430_;
 wire _05431_;
 wire _05432_;
 wire _05433_;
 wire _05434_;
 wire _05435_;
 wire _05436_;
 wire _05437_;
 wire _05438_;
 wire _05439_;
 wire _05440_;
 wire _05441_;
 wire _05442_;
 wire _05443_;
 wire _05444_;
 wire _05445_;
 wire _05446_;
 wire _05447_;
 wire _05448_;
 wire _05449_;
 wire _05450_;
 wire _05451_;
 wire _05452_;
 wire _05453_;
 wire _05454_;
 wire _05455_;
 wire _05456_;
 wire _05457_;
 wire _05458_;
 wire _05459_;
 wire _05460_;
 wire _05461_;
 wire _05462_;
 wire _05463_;
 wire _05464_;
 wire _05465_;
 wire _05466_;
 wire _05467_;
 wire _05468_;
 wire _05469_;
 wire _05470_;
 wire _05471_;
 wire _05472_;
 wire _05473_;
 wire _05474_;
 wire _05475_;
 wire _05476_;
 wire _05477_;
 wire _05478_;
 wire _05479_;
 wire _05480_;
 wire _05481_;
 wire _05482_;
 wire _05483_;
 wire _05484_;
 wire _05485_;
 wire _05486_;
 wire _05487_;
 wire _05488_;
 wire _05489_;
 wire _05490_;
 wire _05491_;
 wire _05492_;
 wire _05493_;
 wire _05494_;
 wire _05495_;
 wire _05496_;
 wire _05497_;
 wire _05498_;
 wire _05499_;
 wire _05500_;
 wire _05501_;
 wire _05502_;
 wire _05503_;
 wire _05504_;
 wire _05505_;
 wire _05506_;
 wire _05507_;
 wire _05508_;
 wire _05509_;
 wire _05510_;
 wire _05511_;
 wire _05512_;
 wire _05513_;
 wire _05514_;
 wire _05515_;
 wire _05516_;
 wire _05517_;
 wire _05518_;
 wire _05519_;
 wire _05520_;
 wire _05521_;
 wire _05522_;
 wire _05523_;
 wire _05524_;
 wire _05525_;
 wire _05526_;
 wire _05527_;
 wire _05528_;
 wire _05529_;
 wire _05530_;
 wire _05531_;
 wire _05532_;
 wire _05533_;
 wire _05534_;
 wire _05535_;
 wire _05536_;
 wire _05537_;
 wire _05538_;
 wire _05539_;
 wire _05540_;
 wire _05541_;
 wire _05542_;
 wire _05543_;
 wire _05544_;
 wire _05545_;
 wire _05546_;
 wire _05547_;
 wire _05548_;
 wire _05549_;
 wire _05550_;
 wire _05551_;
 wire _05552_;
 wire _05553_;
 wire _05554_;
 wire _05555_;
 wire _05556_;
 wire _05557_;
 wire _05558_;
 wire _05559_;
 wire _05560_;
 wire _05561_;
 wire _05562_;
 wire _05563_;
 wire _05564_;
 wire _05565_;
 wire _05566_;
 wire _05567_;
 wire _05568_;
 wire _05569_;
 wire _05570_;
 wire _05571_;
 wire _05572_;
 wire _05573_;
 wire _05574_;
 wire _05575_;
 wire _05576_;
 wire _05577_;
 wire _05578_;
 wire _05579_;
 wire _05580_;
 wire _05581_;
 wire _05582_;
 wire _05583_;
 wire _05584_;
 wire _05585_;
 wire _05586_;
 wire _05587_;
 wire _05588_;
 wire _05589_;
 wire _05590_;
 wire _05591_;
 wire _05592_;
 wire _05593_;
 wire _05594_;
 wire _05595_;
 wire _05596_;
 wire _05597_;
 wire _05598_;
 wire _05599_;
 wire _05600_;
 wire _05601_;
 wire _05602_;
 wire _05603_;
 wire _05604_;
 wire _05605_;
 wire _05606_;
 wire _05607_;
 wire _05608_;
 wire _05609_;
 wire _05610_;
 wire _05611_;
 wire _05612_;
 wire _05613_;
 wire _05614_;
 wire _05615_;
 wire _05616_;
 wire _05617_;
 wire _05618_;
 wire _05619_;
 wire _05620_;
 wire _05621_;
 wire _05622_;
 wire _05623_;
 wire _05624_;
 wire _05625_;
 wire _05626_;
 wire _05627_;
 wire _05628_;
 wire _05629_;
 wire _05630_;
 wire _05631_;
 wire _05632_;
 wire _05633_;
 wire _05634_;
 wire _05635_;
 wire _05636_;
 wire _05637_;
 wire _05638_;
 wire _05639_;
 wire _05640_;
 wire _05641_;
 wire _05642_;
 wire _05643_;
 wire _05644_;
 wire _05645_;
 wire _05646_;
 wire _05647_;
 wire _05648_;
 wire _05649_;
 wire _05650_;
 wire _05651_;
 wire _05652_;
 wire _05653_;
 wire _05654_;
 wire _05655_;
 wire _05656_;
 wire _05657_;
 wire _05658_;
 wire _05659_;
 wire _05660_;
 wire _05661_;
 wire _05662_;
 wire _05663_;
 wire _05664_;
 wire _05665_;
 wire _05666_;
 wire _05667_;
 wire _05668_;
 wire _05669_;
 wire _05670_;
 wire _05671_;
 wire _05672_;
 wire _05673_;
 wire _05674_;
 wire _05675_;
 wire _05676_;
 wire _05677_;
 wire _05678_;
 wire _05679_;
 wire _05680_;
 wire _05681_;
 wire _05682_;
 wire _05683_;
 wire _05684_;
 wire _05685_;
 wire _05686_;
 wire _05687_;
 wire _05688_;
 wire _05689_;
 wire _05690_;
 wire _05691_;
 wire _05692_;
 wire _05693_;
 wire _05694_;
 wire _05695_;
 wire _05696_;
 wire _05697_;
 wire _05698_;
 wire _05699_;
 wire _05700_;
 wire _05701_;
 wire _05702_;
 wire _05703_;
 wire _05704_;
 wire _05705_;
 wire _05706_;
 wire _05707_;
 wire _05708_;
 wire _05709_;
 wire _05710_;
 wire _05711_;
 wire _05712_;
 wire _05713_;
 wire _05714_;
 wire _05715_;
 wire _05716_;
 wire _05717_;
 wire _05718_;
 wire _05719_;
 wire _05720_;
 wire _05721_;
 wire _05722_;
 wire _05723_;
 wire _05724_;
 wire _05725_;
 wire _05726_;
 wire _05727_;
 wire _05728_;
 wire _05729_;
 wire _05730_;
 wire _05731_;
 wire _05732_;
 wire _05733_;
 wire _05734_;
 wire _05735_;
 wire _05736_;
 wire _05737_;
 wire _05738_;
 wire _05739_;
 wire _05740_;
 wire _05741_;
 wire _05742_;
 wire _05743_;
 wire _05744_;
 wire _05745_;
 wire _05746_;
 wire _05747_;
 wire _05748_;
 wire _05749_;
 wire _05750_;
 wire _05751_;
 wire _05752_;
 wire _05753_;
 wire _05754_;
 wire _05755_;
 wire _05756_;
 wire _05757_;
 wire _05758_;
 wire _05759_;
 wire _05760_;
 wire _05761_;
 wire _05762_;
 wire _05763_;
 wire _05764_;
 wire _05765_;
 wire _05766_;
 wire _05767_;
 wire _05768_;
 wire _05769_;
 wire _05770_;
 wire _05771_;
 wire _05772_;
 wire _05773_;
 wire _05774_;
 wire _05775_;
 wire _05776_;
 wire _05777_;
 wire _05778_;
 wire _05779_;
 wire _05780_;
 wire _05781_;
 wire _05782_;
 wire _05783_;
 wire _05784_;
 wire _05785_;
 wire _05786_;
 wire _05787_;
 wire _05788_;
 wire _05789_;
 wire _05790_;
 wire _05791_;
 wire _05792_;
 wire _05793_;
 wire _05794_;
 wire _05795_;
 wire _05796_;
 wire _05797_;
 wire _05798_;
 wire _05799_;
 wire _05800_;
 wire _05801_;
 wire _05802_;
 wire _05803_;
 wire _05804_;
 wire _05805_;
 wire _05806_;
 wire _05807_;
 wire _05808_;
 wire _05809_;
 wire _05810_;
 wire _05811_;
 wire _05812_;
 wire _05813_;
 wire _05814_;
 wire _05815_;
 wire _05816_;
 wire _05817_;
 wire _05818_;
 wire _05819_;
 wire _05820_;
 wire _05821_;
 wire _05822_;
 wire _05823_;
 wire _05824_;
 wire _05825_;
 wire _05826_;
 wire _05827_;
 wire _05828_;
 wire _05829_;
 wire _05830_;
 wire _05831_;
 wire _05832_;
 wire _05833_;
 wire _05834_;
 wire _05835_;
 wire _05836_;
 wire _05837_;
 wire _05838_;
 wire _05839_;
 wire _05840_;
 wire _05841_;
 wire _05842_;
 wire _05843_;
 wire _05844_;
 wire _05845_;
 wire _05846_;
 wire _05847_;
 wire _05848_;
 wire _05849_;
 wire _05850_;
 wire _05851_;
 wire _05852_;
 wire _05853_;
 wire _05854_;
 wire _05855_;
 wire _05856_;
 wire _05857_;
 wire _05858_;
 wire _05859_;
 wire _05860_;
 wire _05861_;
 wire _05862_;
 wire _05863_;
 wire _05864_;
 wire _05865_;
 wire _05866_;
 wire _05867_;
 wire _05868_;
 wire _05869_;
 wire _05870_;
 wire _05871_;
 wire _05872_;
 wire _05873_;
 wire _05874_;
 wire _05875_;
 wire _05876_;
 wire _05877_;
 wire _05878_;
 wire _05879_;
 wire _05880_;
 wire _05881_;
 wire _05882_;
 wire _05883_;
 wire _05884_;
 wire _05885_;
 wire _05886_;
 wire _05887_;
 wire _05888_;
 wire _05889_;
 wire _05890_;
 wire _05891_;
 wire _05892_;
 wire _05893_;
 wire _05894_;
 wire _05895_;
 wire _05896_;
 wire _05897_;
 wire _05898_;
 wire _05899_;
 wire _05900_;
 wire _05901_;
 wire _05902_;
 wire _05903_;
 wire _05904_;
 wire _05905_;
 wire _05906_;
 wire _05907_;
 wire _05908_;
 wire _05909_;
 wire _05910_;
 wire _05911_;
 wire _05912_;
 wire _05913_;
 wire _05914_;
 wire _05915_;
 wire _05916_;
 wire _05917_;
 wire _05918_;
 wire _05919_;
 wire _05920_;
 wire _05921_;
 wire _05922_;
 wire _05923_;
 wire _05924_;
 wire _05925_;
 wire _05926_;
 wire _05927_;
 wire _05928_;
 wire _05929_;
 wire _05930_;
 wire _05931_;
 wire _05932_;
 wire _05933_;
 wire _05934_;
 wire _05935_;
 wire _05936_;
 wire _05937_;
 wire _05938_;
 wire _05939_;
 wire _05940_;
 wire _05941_;
 wire _05942_;
 wire _05943_;
 wire _05944_;
 wire _05945_;
 wire _05946_;
 wire _05947_;
 wire _05948_;
 wire _05949_;
 wire _05950_;
 wire _05951_;
 wire _05952_;
 wire _05953_;
 wire _05954_;
 wire _05955_;
 wire _05956_;
 wire _05957_;
 wire _05958_;
 wire _05959_;
 wire _05960_;
 wire _05961_;
 wire _05962_;
 wire _05963_;
 wire _05964_;
 wire _05965_;
 wire _05966_;
 wire _05967_;
 wire _05968_;
 wire _05969_;
 wire _05970_;
 wire _05971_;
 wire _05972_;
 wire _05973_;
 wire _05974_;
 wire _05975_;
 wire _05976_;
 wire _05977_;
 wire _05978_;
 wire _05979_;
 wire _05980_;
 wire _05981_;
 wire _05982_;
 wire _05983_;
 wire _05984_;
 wire _05985_;
 wire _05986_;
 wire _05987_;
 wire _05988_;
 wire _05989_;
 wire _05990_;
 wire _05991_;
 wire _05992_;
 wire _05993_;
 wire _05994_;
 wire _05995_;
 wire _05996_;
 wire _05997_;
 wire _05998_;
 wire _05999_;
 wire _06000_;
 wire _06001_;
 wire _06002_;
 wire _06003_;
 wire _06004_;
 wire _06005_;
 wire _06006_;
 wire _06007_;
 wire _06008_;
 wire _06009_;
 wire _06010_;
 wire _06011_;
 wire _06012_;
 wire _06013_;
 wire _06014_;
 wire _06015_;
 wire _06016_;
 wire _06017_;
 wire _06018_;
 wire _06019_;
 wire _06020_;
 wire _06021_;
 wire _06022_;
 wire _06023_;
 wire _06024_;
 wire _06025_;
 wire _06026_;
 wire _06027_;
 wire _06028_;
 wire _06029_;
 wire _06030_;
 wire _06031_;
 wire _06032_;
 wire _06033_;
 wire _06034_;
 wire _06035_;
 wire _06036_;
 wire _06037_;
 wire _06038_;
 wire _06039_;
 wire _06040_;
 wire _06041_;
 wire _06042_;
 wire _06043_;
 wire _06044_;
 wire _06045_;
 wire _06046_;
 wire _06047_;
 wire _06048_;
 wire _06049_;
 wire _06050_;
 wire _06051_;
 wire _06052_;
 wire _06053_;
 wire _06054_;
 wire _06055_;
 wire _06056_;
 wire _06057_;
 wire _06058_;
 wire _06059_;
 wire _06060_;
 wire _06061_;
 wire _06062_;
 wire _06063_;
 wire _06064_;
 wire _06065_;
 wire _06066_;
 wire _06067_;
 wire _06068_;
 wire _06069_;
 wire _06070_;
 wire _06071_;
 wire _06072_;
 wire _06073_;
 wire _06074_;
 wire _06075_;
 wire _06076_;
 wire _06077_;
 wire _06078_;
 wire _06079_;
 wire _06080_;
 wire _06081_;
 wire _06082_;
 wire _06083_;
 wire _06084_;
 wire _06085_;
 wire _06086_;
 wire _06087_;
 wire _06088_;
 wire _06089_;
 wire _06090_;
 wire _06091_;
 wire _06092_;
 wire _06093_;
 wire _06094_;
 wire _06095_;
 wire _06096_;
 wire _06097_;
 wire _06098_;
 wire _06099_;
 wire _06100_;
 wire _06101_;
 wire _06102_;
 wire _06103_;
 wire _06104_;
 wire _06105_;
 wire _06106_;
 wire _06107_;
 wire _06108_;
 wire _06109_;
 wire _06110_;
 wire _06111_;
 wire _06112_;
 wire _06113_;
 wire _06114_;
 wire _06115_;
 wire _06116_;
 wire _06117_;
 wire _06118_;
 wire _06119_;
 wire _06120_;
 wire _06121_;
 wire _06122_;
 wire _06123_;
 wire _06124_;
 wire _06125_;
 wire _06126_;
 wire _06127_;
 wire _06128_;
 wire _06129_;
 wire _06130_;
 wire _06131_;
 wire _06132_;
 wire _06133_;
 wire _06134_;
 wire _06135_;
 wire _06136_;
 wire _06137_;
 wire _06138_;
 wire _06139_;
 wire _06140_;
 wire _06141_;
 wire _06142_;
 wire _06143_;
 wire _06144_;
 wire _06145_;
 wire _06146_;
 wire _06147_;
 wire _06148_;
 wire _06149_;
 wire _06150_;
 wire _06151_;
 wire _06152_;
 wire _06153_;
 wire _06154_;
 wire _06155_;
 wire _06156_;
 wire _06157_;
 wire _06158_;
 wire _06159_;
 wire _06160_;
 wire _06161_;
 wire _06162_;
 wire _06163_;
 wire _06164_;
 wire _06165_;
 wire _06166_;
 wire _06167_;
 wire _06168_;
 wire _06169_;
 wire _06170_;
 wire _06171_;
 wire _06172_;
 wire _06173_;
 wire _06174_;
 wire _06175_;
 wire _06176_;
 wire _06177_;
 wire _06178_;
 wire _06179_;
 wire _06180_;
 wire _06181_;
 wire _06182_;
 wire _06183_;
 wire _06184_;
 wire _06185_;
 wire _06186_;
 wire _06187_;
 wire _06188_;
 wire _06189_;
 wire _06190_;
 wire _06191_;
 wire _06192_;
 wire _06193_;
 wire _06194_;
 wire _06195_;
 wire _06196_;
 wire _06197_;
 wire _06198_;
 wire _06199_;
 wire _06200_;
 wire _06201_;
 wire _06202_;
 wire _06203_;
 wire _06204_;
 wire _06205_;
 wire _06206_;
 wire _06207_;
 wire _06208_;
 wire _06209_;
 wire _06210_;
 wire _06211_;
 wire _06212_;
 wire _06213_;
 wire _06214_;
 wire _06215_;
 wire _06216_;
 wire _06217_;
 wire _06218_;
 wire _06219_;
 wire _06220_;
 wire _06221_;
 wire _06222_;
 wire _06223_;
 wire _06224_;
 wire _06225_;
 wire _06226_;
 wire _06227_;
 wire _06228_;
 wire _06229_;
 wire _06230_;
 wire _06231_;
 wire _06232_;
 wire _06233_;
 wire _06234_;
 wire _06235_;
 wire _06236_;
 wire _06237_;
 wire _06238_;
 wire _06239_;
 wire _06240_;
 wire _06241_;
 wire _06242_;
 wire _06243_;
 wire _06244_;
 wire _06245_;
 wire _06246_;
 wire _06247_;
 wire _06248_;
 wire _06249_;
 wire _06250_;
 wire _06251_;
 wire _06252_;
 wire _06253_;
 wire _06254_;
 wire _06255_;
 wire _06256_;
 wire _06257_;
 wire _06258_;
 wire _06259_;
 wire _06260_;
 wire _06261_;
 wire _06262_;
 wire _06263_;
 wire _06264_;
 wire _06265_;
 wire _06266_;
 wire _06267_;
 wire _06268_;
 wire _06269_;
 wire _06270_;
 wire _06271_;
 wire _06272_;
 wire _06273_;
 wire _06274_;
 wire _06275_;
 wire _06276_;
 wire _06277_;
 wire _06278_;
 wire _06279_;
 wire _06280_;
 wire _06281_;
 wire _06282_;
 wire _06283_;
 wire _06284_;
 wire _06285_;
 wire _06286_;
 wire _06287_;
 wire _06288_;
 wire _06289_;
 wire _06290_;
 wire _06291_;
 wire _06292_;
 wire _06293_;
 wire _06294_;
 wire _06295_;
 wire _06296_;
 wire _06297_;
 wire _06298_;
 wire _06299_;
 wire _06300_;
 wire _06301_;
 wire _06302_;
 wire _06303_;
 wire _06304_;
 wire _06305_;
 wire _06306_;
 wire _06307_;
 wire _06308_;
 wire _06309_;
 wire _06310_;
 wire _06311_;
 wire _06312_;
 wire _06313_;
 wire _06314_;
 wire _06315_;
 wire _06316_;
 wire _06317_;
 wire _06318_;
 wire _06319_;
 wire _06320_;
 wire _06321_;
 wire _06322_;
 wire _06323_;
 wire _06324_;
 wire _06325_;
 wire _06326_;
 wire _06327_;
 wire _06328_;
 wire _06329_;
 wire _06330_;
 wire _06331_;
 wire _06332_;
 wire _06333_;
 wire _06334_;
 wire _06335_;
 wire _06336_;
 wire _06337_;
 wire _06338_;
 wire _06339_;
 wire _06340_;
 wire _06341_;
 wire _06342_;
 wire _06343_;
 wire _06344_;
 wire _06345_;
 wire _06346_;
 wire _06347_;
 wire _06348_;
 wire _06349_;
 wire _06350_;
 wire _06351_;
 wire _06352_;
 wire _06353_;
 wire _06354_;
 wire _06355_;
 wire _06356_;
 wire _06357_;
 wire _06358_;
 wire _06359_;
 wire _06360_;
 wire _06361_;
 wire _06362_;
 wire _06363_;
 wire _06364_;
 wire _06365_;
 wire _06366_;
 wire _06367_;
 wire _06368_;
 wire _06369_;
 wire _06370_;
 wire _06371_;
 wire _06372_;
 wire _06373_;
 wire _06374_;
 wire _06375_;
 wire _06376_;
 wire _06377_;
 wire _06378_;
 wire _06379_;
 wire _06380_;
 wire _06381_;
 wire _06382_;
 wire _06383_;
 wire _06384_;
 wire _06385_;
 wire _06386_;
 wire _06387_;
 wire _06388_;
 wire _06389_;
 wire _06390_;
 wire _06391_;
 wire _06392_;
 wire _06393_;
 wire _06394_;
 wire _06395_;
 wire _06396_;
 wire _06397_;
 wire _06398_;
 wire _06399_;
 wire _06400_;
 wire _06401_;
 wire _06402_;
 wire _06403_;
 wire _06404_;
 wire _06405_;
 wire _06406_;
 wire _06407_;
 wire _06408_;
 wire _06409_;
 wire _06410_;
 wire _06411_;
 wire _06412_;
 wire _06413_;
 wire _06414_;
 wire _06415_;
 wire _06416_;
 wire _06417_;
 wire _06418_;
 wire _06419_;
 wire _06420_;
 wire _06421_;
 wire _06422_;
 wire _06423_;
 wire _06424_;
 wire _06425_;
 wire _06426_;
 wire _06427_;
 wire _06428_;
 wire _06429_;
 wire _06430_;
 wire _06431_;
 wire _06432_;
 wire _06433_;
 wire _06434_;
 wire _06435_;
 wire _06436_;
 wire _06437_;
 wire _06438_;
 wire _06439_;
 wire _06440_;
 wire _06441_;
 wire _06442_;
 wire _06443_;
 wire _06444_;
 wire _06445_;
 wire _06446_;
 wire _06447_;
 wire _06448_;
 wire _06449_;
 wire _06450_;
 wire _06451_;
 wire _06452_;
 wire _06453_;
 wire _06454_;
 wire _06455_;
 wire _06456_;
 wire _06457_;
 wire _06458_;
 wire _06459_;
 wire _06460_;
 wire _06461_;
 wire _06462_;
 wire _06463_;
 wire _06464_;
 wire _06465_;
 wire _06466_;
 wire _06467_;
 wire _06468_;
 wire _06469_;
 wire _06470_;
 wire _06471_;
 wire _06472_;
 wire _06473_;
 wire _06474_;
 wire _06475_;
 wire _06476_;
 wire _06477_;
 wire _06478_;
 wire _06479_;
 wire _06480_;
 wire _06481_;
 wire _06482_;
 wire _06483_;
 wire _06484_;
 wire _06485_;
 wire _06486_;
 wire _06487_;
 wire _06488_;
 wire _06489_;
 wire _06490_;
 wire _06491_;
 wire _06492_;
 wire _06493_;
 wire _06494_;
 wire _06495_;
 wire _06496_;
 wire _06497_;
 wire _06498_;
 wire _06499_;
 wire _06500_;
 wire _06501_;
 wire _06502_;
 wire _06503_;
 wire _06504_;
 wire _06505_;
 wire _06506_;
 wire _06507_;
 wire _06508_;
 wire _06509_;
 wire _06510_;
 wire _06511_;
 wire _06512_;
 wire _06513_;
 wire _06514_;
 wire _06515_;
 wire _06516_;
 wire _06517_;
 wire _06518_;
 wire _06519_;
 wire _06520_;
 wire _06521_;
 wire _06522_;
 wire _06523_;
 wire _06524_;
 wire _06525_;
 wire _06526_;
 wire _06527_;
 wire _06528_;
 wire _06529_;
 wire _06530_;
 wire _06531_;
 wire _06532_;
 wire _06533_;
 wire _06534_;
 wire _06535_;
 wire _06536_;
 wire _06537_;
 wire _06538_;
 wire _06539_;
 wire _06540_;
 wire _06541_;
 wire _06542_;
 wire _06543_;
 wire _06544_;
 wire _06545_;
 wire _06546_;
 wire _06547_;
 wire _06548_;
 wire _06549_;
 wire _06550_;
 wire _06551_;
 wire _06552_;
 wire _06553_;
 wire _06554_;
 wire _06555_;
 wire _06556_;
 wire _06557_;
 wire _06558_;
 wire _06559_;
 wire _06560_;
 wire _06561_;
 wire _06562_;
 wire _06563_;
 wire _06564_;
 wire _06565_;
 wire _06566_;
 wire _06567_;
 wire _06568_;
 wire _06569_;
 wire _06570_;
 wire _06571_;
 wire _06572_;
 wire _06573_;
 wire _06574_;
 wire _06575_;
 wire _06576_;
 wire _06577_;
 wire _06578_;
 wire _06579_;
 wire _06580_;
 wire _06581_;
 wire _06582_;
 wire _06583_;
 wire _06584_;
 wire _06585_;
 wire _06586_;
 wire _06587_;
 wire _06588_;
 wire _06589_;
 wire _06590_;
 wire _06591_;
 wire _06592_;
 wire _06593_;
 wire _06594_;
 wire _06595_;
 wire _06596_;
 wire _06597_;
 wire _06598_;
 wire _06599_;
 wire _06600_;
 wire _06601_;
 wire _06602_;
 wire _06603_;
 wire _06604_;
 wire _06605_;
 wire _06606_;
 wire _06607_;
 wire _06608_;
 wire _06609_;
 wire _06610_;
 wire _06611_;
 wire _06612_;
 wire _06613_;
 wire _06614_;
 wire _06615_;
 wire _06616_;
 wire _06617_;
 wire _06618_;
 wire _06619_;
 wire _06620_;
 wire _06621_;
 wire _06622_;
 wire _06623_;
 wire _06624_;
 wire _06625_;
 wire _06626_;
 wire _06627_;
 wire _06628_;
 wire _06629_;
 wire _06630_;
 wire _06631_;
 wire _06632_;
 wire _06633_;
 wire _06634_;
 wire _06635_;
 wire _06636_;
 wire _06637_;
 wire _06638_;
 wire _06639_;
 wire _06640_;
 wire _06641_;
 wire _06642_;
 wire _06643_;
 wire _06644_;
 wire _06645_;
 wire _06646_;
 wire _06647_;
 wire _06648_;
 wire _06649_;
 wire _06650_;
 wire _06651_;
 wire _06652_;
 wire _06653_;
 wire _06654_;
 wire _06655_;
 wire _06656_;
 wire _06657_;
 wire _06658_;
 wire _06659_;
 wire _06660_;
 wire _06661_;
 wire _06662_;
 wire _06663_;
 wire _06664_;
 wire _06665_;
 wire _06666_;
 wire _06667_;
 wire _06668_;
 wire _06669_;
 wire _06670_;
 wire _06671_;
 wire _06672_;
 wire _06673_;
 wire _06674_;
 wire _06675_;
 wire _06676_;
 wire _06677_;
 wire _06678_;
 wire _06679_;
 wire _06680_;
 wire _06681_;
 wire _06682_;
 wire _06683_;
 wire _06684_;
 wire _06685_;
 wire _06686_;
 wire _06687_;
 wire _06688_;
 wire _06689_;
 wire _06690_;
 wire _06691_;
 wire _06692_;
 wire _06693_;
 wire _06694_;
 wire _06695_;
 wire _06696_;
 wire _06697_;
 wire _06698_;
 wire _06699_;
 wire _06700_;
 wire _06701_;
 wire _06702_;
 wire _06703_;
 wire _06704_;
 wire _06705_;
 wire _06706_;
 wire _06707_;
 wire _06708_;
 wire _06709_;
 wire _06710_;
 wire _06711_;
 wire _06712_;
 wire _06713_;
 wire _06714_;
 wire _06715_;
 wire _06716_;
 wire _06717_;
 wire _06718_;
 wire _06719_;
 wire _06720_;
 wire _06721_;
 wire _06722_;
 wire _06723_;
 wire _06724_;
 wire _06725_;
 wire _06726_;
 wire _06727_;
 wire _06728_;
 wire _06729_;
 wire _06730_;
 wire _06731_;
 wire _06732_;
 wire _06733_;
 wire _06734_;
 wire _06735_;
 wire _06736_;
 wire _06737_;
 wire _06738_;
 wire _06739_;
 wire _06740_;
 wire _06741_;
 wire _06742_;
 wire _06743_;
 wire _06744_;
 wire _06745_;
 wire _06746_;
 wire _06747_;
 wire _06748_;
 wire _06749_;
 wire _06750_;
 wire _06751_;
 wire _06752_;
 wire _06753_;
 wire _06754_;
 wire _06755_;
 wire _06756_;
 wire _06757_;
 wire _06758_;
 wire _06759_;
 wire _06760_;
 wire _06761_;
 wire _06762_;
 wire _06763_;
 wire _06764_;
 wire _06765_;
 wire _06766_;
 wire _06767_;
 wire _06768_;
 wire _06769_;
 wire _06770_;
 wire _06771_;
 wire _06772_;
 wire _06773_;
 wire _06774_;
 wire _06775_;
 wire _06776_;
 wire _06777_;
 wire _06778_;
 wire _06779_;
 wire _06780_;
 wire _06781_;
 wire _06782_;
 wire _06783_;
 wire _06784_;
 wire _06785_;
 wire _06786_;
 wire _06787_;
 wire _06788_;
 wire _06789_;
 wire _06790_;
 wire _06791_;
 wire _06792_;
 wire _06793_;
 wire _06794_;
 wire _06795_;
 wire _06796_;
 wire _06797_;
 wire _06798_;
 wire _06799_;
 wire _06800_;
 wire _06801_;
 wire _06802_;
 wire _06803_;
 wire _06804_;
 wire _06805_;
 wire _06806_;
 wire _06807_;
 wire _06808_;
 wire _06809_;
 wire _06810_;
 wire _06811_;
 wire _06812_;
 wire _06813_;
 wire _06814_;
 wire _06815_;
 wire _06816_;
 wire _06817_;
 wire _06818_;
 wire _06819_;
 wire _06820_;
 wire _06821_;
 wire _06822_;
 wire _06823_;
 wire _06824_;
 wire _06825_;
 wire _06826_;
 wire _06827_;
 wire _06828_;
 wire _06829_;
 wire _06830_;
 wire _06831_;
 wire _06832_;
 wire _06833_;
 wire _06834_;
 wire _06835_;
 wire _06836_;
 wire _06837_;
 wire _06838_;
 wire _06839_;
 wire _06840_;
 wire _06841_;
 wire _06842_;
 wire _06843_;
 wire _06844_;
 wire _06845_;
 wire _06846_;
 wire _06847_;
 wire _06848_;
 wire _06849_;
 wire _06850_;
 wire _06851_;
 wire _06852_;
 wire _06853_;
 wire _06854_;
 wire _06855_;
 wire _06856_;
 wire _06857_;
 wire _06858_;
 wire _06859_;
 wire _06860_;
 wire _06861_;
 wire _06862_;
 wire _06863_;
 wire _06864_;
 wire _06865_;
 wire _06866_;
 wire _06867_;
 wire _06868_;
 wire _06869_;
 wire _06870_;
 wire _06871_;
 wire _06872_;
 wire _06873_;
 wire _06874_;
 wire _06875_;
 wire _06876_;
 wire _06877_;
 wire _06878_;
 wire _06879_;
 wire _06880_;
 wire _06881_;
 wire _06882_;
 wire _06883_;
 wire _06884_;
 wire _06885_;
 wire _06886_;
 wire _06887_;
 wire _06888_;
 wire _06889_;
 wire _06890_;
 wire _06891_;
 wire _06892_;
 wire _06893_;
 wire _06894_;
 wire _06895_;
 wire _06896_;
 wire _06897_;
 wire _06898_;
 wire _06899_;
 wire _06900_;
 wire _06901_;
 wire _06902_;
 wire _06903_;
 wire _06904_;
 wire _06905_;
 wire _06906_;
 wire _06907_;
 wire _06908_;
 wire _06909_;
 wire _06910_;
 wire _06911_;
 wire _06912_;
 wire _06913_;
 wire _06914_;
 wire _06915_;
 wire _06916_;
 wire _06917_;
 wire _06918_;
 wire _06919_;
 wire _06920_;
 wire _06921_;
 wire _06922_;
 wire _06923_;
 wire _06924_;
 wire _06925_;
 wire _06926_;
 wire _06927_;
 wire _06928_;
 wire _06929_;
 wire _06930_;
 wire _06931_;
 wire _06932_;
 wire _06933_;
 wire _06934_;
 wire _06935_;
 wire _06936_;
 wire _06937_;
 wire _06938_;
 wire _06939_;
 wire _06940_;
 wire _06941_;
 wire _06942_;
 wire _06943_;
 wire _06944_;
 wire _06945_;
 wire _06946_;
 wire _06947_;
 wire _06948_;
 wire _06949_;
 wire _06950_;
 wire _06951_;
 wire _06952_;
 wire _06953_;
 wire _06954_;
 wire _06955_;
 wire _06956_;
 wire _06957_;
 wire _06958_;
 wire _06959_;
 wire _06960_;
 wire _06961_;
 wire _06962_;
 wire _06963_;
 wire _06964_;
 wire _06965_;
 wire _06966_;
 wire _06967_;
 wire clknet_leaf_0_clk_p2c;
 wire aux_enable_p2c;
 wire clk_p2c;
 wire data_in_p2c_1;
 wire data_in_p2c_2;
 wire data_in_p2c_3;
 wire data_in_p2c_4;
 wire data_in_p2c_5;
 wire data_in_p2c_6;
 wire data_in_p2c_7;
 wire data_in_p2c_8;
 wire net4049;
 wire net32;
 wire net22;
 wire net17;
 wire net4032;
 wire net8;
 wire net4017;
 wire net4016;
 wire lfsr_out_c2p;
 wire \median_processor.input_storage[0] ;
 wire \median_processor.input_storage[10] ;
 wire \median_processor.input_storage[11] ;
 wire \median_processor.input_storage[12] ;
 wire \median_processor.input_storage[13] ;
 wire \median_processor.input_storage[14] ;
 wire \median_processor.input_storage[15] ;
 wire \median_processor.input_storage[16] ;
 wire \median_processor.input_storage[17] ;
 wire \median_processor.input_storage[18] ;
 wire \median_processor.input_storage[19] ;
 wire \median_processor.input_storage[1] ;
 wire \median_processor.input_storage[20] ;
 wire \median_processor.input_storage[21] ;
 wire \median_processor.input_storage[22] ;
 wire \median_processor.input_storage[23] ;
 wire \median_processor.input_storage[24] ;
 wire \median_processor.input_storage[25] ;
 wire \median_processor.input_storage[26] ;
 wire \median_processor.input_storage[27] ;
 wire \median_processor.input_storage[28] ;
 wire \median_processor.input_storage[29] ;
 wire \median_processor.input_storage[2] ;
 wire \median_processor.input_storage[30] ;
 wire \median_processor.input_storage[31] ;
 wire \median_processor.input_storage[32] ;
 wire \median_processor.input_storage[33] ;
 wire \median_processor.input_storage[34] ;
 wire \median_processor.input_storage[35] ;
 wire \median_processor.input_storage[36] ;
 wire \median_processor.input_storage[37] ;
 wire \median_processor.input_storage[38] ;
 wire \median_processor.input_storage[39] ;
 wire \median_processor.input_storage[3] ;
 wire \median_processor.input_storage[40] ;
 wire \median_processor.input_storage[41] ;
 wire \median_processor.input_storage[42] ;
 wire \median_processor.input_storage[43] ;
 wire \median_processor.input_storage[44] ;
 wire \median_processor.input_storage[45] ;
 wire \median_processor.input_storage[46] ;
 wire \median_processor.input_storage[47] ;
 wire \median_processor.input_storage[48] ;
 wire \median_processor.input_storage[49] ;
 wire \median_processor.input_storage[4] ;
 wire \median_processor.input_storage[50] ;
 wire \median_processor.input_storage[51] ;
 wire \median_processor.input_storage[52] ;
 wire \median_processor.input_storage[53] ;
 wire \median_processor.input_storage[54] ;
 wire \median_processor.input_storage[55] ;
 wire \median_processor.input_storage[56] ;
 wire \median_processor.input_storage[57] ;
 wire \median_processor.input_storage[58] ;
 wire \median_processor.input_storage[59] ;
 wire \median_processor.input_storage[5] ;
 wire \median_processor.input_storage[60] ;
 wire \median_processor.input_storage[61] ;
 wire \median_processor.input_storage[62] ;
 wire \median_processor.input_storage[63] ;
 wire \median_processor.input_storage[6] ;
 wire \median_processor.input_storage[7] ;
 wire \median_processor.input_storage[8] ;
 wire \median_processor.input_storage[9] ;
 wire \median_processor.median_processor.median_out[0] ;
 wire \median_processor.median_processor.median_out[1] ;
 wire \median_processor.median_processor.median_out[2] ;
 wire \median_processor.median_processor.median_out[3] ;
 wire \median_processor.median_processor.median_out[4] ;
 wire \median_processor.median_processor.median_out[5] ;
 wire \median_processor.median_processor.median_out[6] ;
 wire \median_processor.median_processor.median_out[7] ;
 wire \median_processor.rst ;
 wire \median_processor.wr_enable ;
 wire out_select_p2c_1;
 wire out_select_p2c_2;
 wire \rando_generator.lfsr_reg[10] ;
 wire \rando_generator.lfsr_reg[11] ;
 wire \rando_generator.lfsr_reg[12] ;
 wire \rando_generator.lfsr_reg[13] ;
 wire \rando_generator.lfsr_reg[14] ;
 wire \rando_generator.lfsr_reg[15] ;
 wire \rando_generator.lfsr_reg[16] ;
 wire \rando_generator.lfsr_reg[17] ;
 wire \rando_generator.lfsr_reg[18] ;
 wire \rando_generator.lfsr_reg[19] ;
 wire \rando_generator.lfsr_reg[1] ;
 wire \rando_generator.lfsr_reg[20] ;
 wire \rando_generator.lfsr_reg[21] ;
 wire \rando_generator.lfsr_reg[22] ;
 wire \rando_generator.lfsr_reg[23] ;
 wire \rando_generator.lfsr_reg[24] ;
 wire \rando_generator.lfsr_reg[25] ;
 wire \rando_generator.lfsr_reg[26] ;
 wire \rando_generator.lfsr_reg[27] ;
 wire \rando_generator.lfsr_reg[28] ;
 wire \rando_generator.lfsr_reg[29] ;
 wire \rando_generator.lfsr_reg[2] ;
 wire \rando_generator.lfsr_reg[30] ;
 wire \rando_generator.lfsr_reg[3] ;
 wire \rando_generator.lfsr_reg[4] ;
 wire \rando_generator.lfsr_reg[5] ;
 wire \rando_generator.lfsr_reg[6] ;
 wire \rando_generator.lfsr_reg[7] ;
 wire \rando_generator.lfsr_reg[8] ;
 wire \rando_generator.lfsr_reg[9] ;
 wire reg_addr_p2c_1;
 wire reg_addr_p2c_2;
 wire reg_addr_p2c_3;
 wire \shift_storage.shreg_in ;
 wire \shift_storage.shreg_out ;
 wire \shift_storage.storage[0] ;
 wire \shift_storage.storage[1000] ;
 wire \shift_storage.storage[1001] ;
 wire \shift_storage.storage[1002] ;
 wire \shift_storage.storage[1003] ;
 wire \shift_storage.storage[1004] ;
 wire \shift_storage.storage[1005] ;
 wire \shift_storage.storage[1006] ;
 wire \shift_storage.storage[1007] ;
 wire \shift_storage.storage[1008] ;
 wire \shift_storage.storage[1009] ;
 wire \shift_storage.storage[100] ;
 wire \shift_storage.storage[1010] ;
 wire \shift_storage.storage[1011] ;
 wire \shift_storage.storage[1012] ;
 wire \shift_storage.storage[1013] ;
 wire \shift_storage.storage[1014] ;
 wire \shift_storage.storage[1015] ;
 wire \shift_storage.storage[1016] ;
 wire \shift_storage.storage[1017] ;
 wire \shift_storage.storage[1018] ;
 wire \shift_storage.storage[1019] ;
 wire \shift_storage.storage[101] ;
 wire \shift_storage.storage[1020] ;
 wire \shift_storage.storage[1021] ;
 wire \shift_storage.storage[1022] ;
 wire \shift_storage.storage[1023] ;
 wire \shift_storage.storage[1024] ;
 wire \shift_storage.storage[1025] ;
 wire \shift_storage.storage[1026] ;
 wire \shift_storage.storage[1027] ;
 wire \shift_storage.storage[1028] ;
 wire \shift_storage.storage[1029] ;
 wire \shift_storage.storage[102] ;
 wire \shift_storage.storage[1030] ;
 wire \shift_storage.storage[1031] ;
 wire \shift_storage.storage[1032] ;
 wire \shift_storage.storage[1033] ;
 wire \shift_storage.storage[1034] ;
 wire \shift_storage.storage[1035] ;
 wire \shift_storage.storage[1036] ;
 wire \shift_storage.storage[1037] ;
 wire \shift_storage.storage[1038] ;
 wire \shift_storage.storage[1039] ;
 wire \shift_storage.storage[103] ;
 wire \shift_storage.storage[1040] ;
 wire \shift_storage.storage[1041] ;
 wire \shift_storage.storage[1042] ;
 wire \shift_storage.storage[1043] ;
 wire \shift_storage.storage[1044] ;
 wire \shift_storage.storage[1045] ;
 wire \shift_storage.storage[1046] ;
 wire \shift_storage.storage[1047] ;
 wire \shift_storage.storage[1048] ;
 wire \shift_storage.storage[1049] ;
 wire \shift_storage.storage[104] ;
 wire \shift_storage.storage[1050] ;
 wire \shift_storage.storage[1051] ;
 wire \shift_storage.storage[1052] ;
 wire \shift_storage.storage[1053] ;
 wire \shift_storage.storage[1054] ;
 wire \shift_storage.storage[1055] ;
 wire \shift_storage.storage[1056] ;
 wire \shift_storage.storage[1057] ;
 wire \shift_storage.storage[1058] ;
 wire \shift_storage.storage[1059] ;
 wire \shift_storage.storage[105] ;
 wire \shift_storage.storage[1060] ;
 wire \shift_storage.storage[1061] ;
 wire \shift_storage.storage[1062] ;
 wire \shift_storage.storage[1063] ;
 wire \shift_storage.storage[1064] ;
 wire \shift_storage.storage[1065] ;
 wire \shift_storage.storage[1066] ;
 wire \shift_storage.storage[1067] ;
 wire \shift_storage.storage[1068] ;
 wire \shift_storage.storage[1069] ;
 wire \shift_storage.storage[106] ;
 wire \shift_storage.storage[1070] ;
 wire \shift_storage.storage[1071] ;
 wire \shift_storage.storage[1072] ;
 wire \shift_storage.storage[1073] ;
 wire \shift_storage.storage[1074] ;
 wire \shift_storage.storage[1075] ;
 wire \shift_storage.storage[1076] ;
 wire \shift_storage.storage[1077] ;
 wire \shift_storage.storage[1078] ;
 wire \shift_storage.storage[1079] ;
 wire \shift_storage.storage[107] ;
 wire \shift_storage.storage[1080] ;
 wire \shift_storage.storage[1081] ;
 wire \shift_storage.storage[1082] ;
 wire \shift_storage.storage[1083] ;
 wire \shift_storage.storage[1084] ;
 wire \shift_storage.storage[1085] ;
 wire \shift_storage.storage[1086] ;
 wire \shift_storage.storage[1087] ;
 wire \shift_storage.storage[1088] ;
 wire \shift_storage.storage[1089] ;
 wire \shift_storage.storage[108] ;
 wire \shift_storage.storage[1090] ;
 wire \shift_storage.storage[1091] ;
 wire \shift_storage.storage[1092] ;
 wire \shift_storage.storage[1093] ;
 wire \shift_storage.storage[1094] ;
 wire \shift_storage.storage[1095] ;
 wire \shift_storage.storage[1096] ;
 wire \shift_storage.storage[1097] ;
 wire \shift_storage.storage[1098] ;
 wire \shift_storage.storage[1099] ;
 wire \shift_storage.storage[109] ;
 wire \shift_storage.storage[10] ;
 wire \shift_storage.storage[1100] ;
 wire \shift_storage.storage[1101] ;
 wire \shift_storage.storage[1102] ;
 wire \shift_storage.storage[1103] ;
 wire \shift_storage.storage[1104] ;
 wire \shift_storage.storage[1105] ;
 wire \shift_storage.storage[1106] ;
 wire \shift_storage.storage[1107] ;
 wire \shift_storage.storage[1108] ;
 wire \shift_storage.storage[1109] ;
 wire \shift_storage.storage[110] ;
 wire \shift_storage.storage[1110] ;
 wire \shift_storage.storage[1111] ;
 wire \shift_storage.storage[1112] ;
 wire \shift_storage.storage[1113] ;
 wire \shift_storage.storage[1114] ;
 wire \shift_storage.storage[1115] ;
 wire \shift_storage.storage[1116] ;
 wire \shift_storage.storage[1117] ;
 wire \shift_storage.storage[1118] ;
 wire \shift_storage.storage[1119] ;
 wire \shift_storage.storage[111] ;
 wire \shift_storage.storage[1120] ;
 wire \shift_storage.storage[1121] ;
 wire \shift_storage.storage[1122] ;
 wire \shift_storage.storage[1123] ;
 wire \shift_storage.storage[1124] ;
 wire \shift_storage.storage[1125] ;
 wire \shift_storage.storage[1126] ;
 wire \shift_storage.storage[1127] ;
 wire \shift_storage.storage[1128] ;
 wire \shift_storage.storage[1129] ;
 wire \shift_storage.storage[112] ;
 wire \shift_storage.storage[1130] ;
 wire \shift_storage.storage[1131] ;
 wire \shift_storage.storage[1132] ;
 wire \shift_storage.storage[1133] ;
 wire \shift_storage.storage[1134] ;
 wire \shift_storage.storage[1135] ;
 wire \shift_storage.storage[1136] ;
 wire \shift_storage.storage[1137] ;
 wire \shift_storage.storage[1138] ;
 wire \shift_storage.storage[1139] ;
 wire \shift_storage.storage[113] ;
 wire \shift_storage.storage[1140] ;
 wire \shift_storage.storage[1141] ;
 wire \shift_storage.storage[1142] ;
 wire \shift_storage.storage[1143] ;
 wire \shift_storage.storage[1144] ;
 wire \shift_storage.storage[1145] ;
 wire \shift_storage.storage[1146] ;
 wire \shift_storage.storage[1147] ;
 wire \shift_storage.storage[1148] ;
 wire \shift_storage.storage[1149] ;
 wire \shift_storage.storage[114] ;
 wire \shift_storage.storage[1150] ;
 wire \shift_storage.storage[1151] ;
 wire \shift_storage.storage[1152] ;
 wire \shift_storage.storage[1153] ;
 wire \shift_storage.storage[1154] ;
 wire \shift_storage.storage[1155] ;
 wire \shift_storage.storage[1156] ;
 wire \shift_storage.storage[1157] ;
 wire \shift_storage.storage[1158] ;
 wire \shift_storage.storage[1159] ;
 wire \shift_storage.storage[115] ;
 wire \shift_storage.storage[1160] ;
 wire \shift_storage.storage[1161] ;
 wire \shift_storage.storage[1162] ;
 wire \shift_storage.storage[1163] ;
 wire \shift_storage.storage[1164] ;
 wire \shift_storage.storage[1165] ;
 wire \shift_storage.storage[1166] ;
 wire \shift_storage.storage[1167] ;
 wire \shift_storage.storage[1168] ;
 wire \shift_storage.storage[1169] ;
 wire \shift_storage.storage[116] ;
 wire \shift_storage.storage[1170] ;
 wire \shift_storage.storage[1171] ;
 wire \shift_storage.storage[1172] ;
 wire \shift_storage.storage[1173] ;
 wire \shift_storage.storage[1174] ;
 wire \shift_storage.storage[1175] ;
 wire \shift_storage.storage[1176] ;
 wire \shift_storage.storage[1177] ;
 wire \shift_storage.storage[1178] ;
 wire \shift_storage.storage[1179] ;
 wire \shift_storage.storage[117] ;
 wire \shift_storage.storage[1180] ;
 wire \shift_storage.storage[1181] ;
 wire \shift_storage.storage[1182] ;
 wire \shift_storage.storage[1183] ;
 wire \shift_storage.storage[1184] ;
 wire \shift_storage.storage[1185] ;
 wire \shift_storage.storage[1186] ;
 wire \shift_storage.storage[1187] ;
 wire \shift_storage.storage[1188] ;
 wire \shift_storage.storage[1189] ;
 wire \shift_storage.storage[118] ;
 wire \shift_storage.storage[1190] ;
 wire \shift_storage.storage[1191] ;
 wire \shift_storage.storage[1192] ;
 wire \shift_storage.storage[1193] ;
 wire \shift_storage.storage[1194] ;
 wire \shift_storage.storage[1195] ;
 wire \shift_storage.storage[1196] ;
 wire \shift_storage.storage[1197] ;
 wire \shift_storage.storage[1198] ;
 wire \shift_storage.storage[1199] ;
 wire \shift_storage.storage[119] ;
 wire \shift_storage.storage[11] ;
 wire \shift_storage.storage[1200] ;
 wire \shift_storage.storage[1201] ;
 wire \shift_storage.storage[1202] ;
 wire \shift_storage.storage[1203] ;
 wire \shift_storage.storage[1204] ;
 wire \shift_storage.storage[1205] ;
 wire \shift_storage.storage[1206] ;
 wire \shift_storage.storage[1207] ;
 wire \shift_storage.storage[1208] ;
 wire \shift_storage.storage[1209] ;
 wire \shift_storage.storage[120] ;
 wire \shift_storage.storage[1210] ;
 wire \shift_storage.storage[1211] ;
 wire \shift_storage.storage[1212] ;
 wire \shift_storage.storage[1213] ;
 wire \shift_storage.storage[1214] ;
 wire \shift_storage.storage[1215] ;
 wire \shift_storage.storage[1216] ;
 wire \shift_storage.storage[1217] ;
 wire \shift_storage.storage[1218] ;
 wire \shift_storage.storage[1219] ;
 wire \shift_storage.storage[121] ;
 wire \shift_storage.storage[1220] ;
 wire \shift_storage.storage[1221] ;
 wire \shift_storage.storage[1222] ;
 wire \shift_storage.storage[1223] ;
 wire \shift_storage.storage[1224] ;
 wire \shift_storage.storage[1225] ;
 wire \shift_storage.storage[1226] ;
 wire \shift_storage.storage[1227] ;
 wire \shift_storage.storage[1228] ;
 wire \shift_storage.storage[1229] ;
 wire \shift_storage.storage[122] ;
 wire \shift_storage.storage[1230] ;
 wire \shift_storage.storage[1231] ;
 wire \shift_storage.storage[1232] ;
 wire \shift_storage.storage[1233] ;
 wire \shift_storage.storage[1234] ;
 wire \shift_storage.storage[1235] ;
 wire \shift_storage.storage[1236] ;
 wire \shift_storage.storage[1237] ;
 wire \shift_storage.storage[1238] ;
 wire \shift_storage.storage[1239] ;
 wire \shift_storage.storage[123] ;
 wire \shift_storage.storage[1240] ;
 wire \shift_storage.storage[1241] ;
 wire \shift_storage.storage[1242] ;
 wire \shift_storage.storage[1243] ;
 wire \shift_storage.storage[1244] ;
 wire \shift_storage.storage[1245] ;
 wire \shift_storage.storage[1246] ;
 wire \shift_storage.storage[1247] ;
 wire \shift_storage.storage[1248] ;
 wire \shift_storage.storage[1249] ;
 wire \shift_storage.storage[124] ;
 wire \shift_storage.storage[1250] ;
 wire \shift_storage.storage[1251] ;
 wire \shift_storage.storage[1252] ;
 wire \shift_storage.storage[1253] ;
 wire \shift_storage.storage[1254] ;
 wire \shift_storage.storage[1255] ;
 wire \shift_storage.storage[1256] ;
 wire \shift_storage.storage[1257] ;
 wire \shift_storage.storage[1258] ;
 wire \shift_storage.storage[1259] ;
 wire \shift_storage.storage[125] ;
 wire \shift_storage.storage[1260] ;
 wire \shift_storage.storage[1261] ;
 wire \shift_storage.storage[1262] ;
 wire \shift_storage.storage[1263] ;
 wire \shift_storage.storage[1264] ;
 wire \shift_storage.storage[1265] ;
 wire \shift_storage.storage[1266] ;
 wire \shift_storage.storage[1267] ;
 wire \shift_storage.storage[1268] ;
 wire \shift_storage.storage[1269] ;
 wire \shift_storage.storage[126] ;
 wire \shift_storage.storage[1270] ;
 wire \shift_storage.storage[1271] ;
 wire \shift_storage.storage[1272] ;
 wire \shift_storage.storage[1273] ;
 wire \shift_storage.storage[1274] ;
 wire \shift_storage.storage[1275] ;
 wire \shift_storage.storage[1276] ;
 wire \shift_storage.storage[1277] ;
 wire \shift_storage.storage[1278] ;
 wire \shift_storage.storage[1279] ;
 wire \shift_storage.storage[127] ;
 wire \shift_storage.storage[1280] ;
 wire \shift_storage.storage[1281] ;
 wire \shift_storage.storage[1282] ;
 wire \shift_storage.storage[1283] ;
 wire \shift_storage.storage[1284] ;
 wire \shift_storage.storage[1285] ;
 wire \shift_storage.storage[1286] ;
 wire \shift_storage.storage[1287] ;
 wire \shift_storage.storage[1288] ;
 wire \shift_storage.storage[1289] ;
 wire \shift_storage.storage[128] ;
 wire \shift_storage.storage[1290] ;
 wire \shift_storage.storage[1291] ;
 wire \shift_storage.storage[1292] ;
 wire \shift_storage.storage[1293] ;
 wire \shift_storage.storage[1294] ;
 wire \shift_storage.storage[1295] ;
 wire \shift_storage.storage[1296] ;
 wire \shift_storage.storage[1297] ;
 wire \shift_storage.storage[1298] ;
 wire \shift_storage.storage[1299] ;
 wire \shift_storage.storage[129] ;
 wire \shift_storage.storage[12] ;
 wire \shift_storage.storage[1300] ;
 wire \shift_storage.storage[1301] ;
 wire \shift_storage.storage[1302] ;
 wire \shift_storage.storage[1303] ;
 wire \shift_storage.storage[1304] ;
 wire \shift_storage.storage[1305] ;
 wire \shift_storage.storage[1306] ;
 wire \shift_storage.storage[1307] ;
 wire \shift_storage.storage[1308] ;
 wire \shift_storage.storage[1309] ;
 wire \shift_storage.storage[130] ;
 wire \shift_storage.storage[1310] ;
 wire \shift_storage.storage[1311] ;
 wire \shift_storage.storage[1312] ;
 wire \shift_storage.storage[1313] ;
 wire \shift_storage.storage[1314] ;
 wire \shift_storage.storage[1315] ;
 wire \shift_storage.storage[1316] ;
 wire \shift_storage.storage[1317] ;
 wire \shift_storage.storage[1318] ;
 wire \shift_storage.storage[1319] ;
 wire \shift_storage.storage[131] ;
 wire \shift_storage.storage[1320] ;
 wire \shift_storage.storage[1321] ;
 wire \shift_storage.storage[1322] ;
 wire \shift_storage.storage[1323] ;
 wire \shift_storage.storage[1324] ;
 wire \shift_storage.storage[1325] ;
 wire \shift_storage.storage[1326] ;
 wire \shift_storage.storage[1327] ;
 wire \shift_storage.storage[1328] ;
 wire \shift_storage.storage[1329] ;
 wire \shift_storage.storage[132] ;
 wire \shift_storage.storage[1330] ;
 wire \shift_storage.storage[1331] ;
 wire \shift_storage.storage[1332] ;
 wire \shift_storage.storage[1333] ;
 wire \shift_storage.storage[1334] ;
 wire \shift_storage.storage[1335] ;
 wire \shift_storage.storage[1336] ;
 wire \shift_storage.storage[1337] ;
 wire \shift_storage.storage[1338] ;
 wire \shift_storage.storage[1339] ;
 wire \shift_storage.storage[133] ;
 wire \shift_storage.storage[1340] ;
 wire \shift_storage.storage[1341] ;
 wire \shift_storage.storage[1342] ;
 wire \shift_storage.storage[1343] ;
 wire \shift_storage.storage[1344] ;
 wire \shift_storage.storage[1345] ;
 wire \shift_storage.storage[1346] ;
 wire \shift_storage.storage[1347] ;
 wire \shift_storage.storage[1348] ;
 wire \shift_storage.storage[1349] ;
 wire \shift_storage.storage[134] ;
 wire \shift_storage.storage[1350] ;
 wire \shift_storage.storage[1351] ;
 wire \shift_storage.storage[1352] ;
 wire \shift_storage.storage[1353] ;
 wire \shift_storage.storage[1354] ;
 wire \shift_storage.storage[1355] ;
 wire \shift_storage.storage[1356] ;
 wire \shift_storage.storage[1357] ;
 wire \shift_storage.storage[1358] ;
 wire \shift_storage.storage[1359] ;
 wire \shift_storage.storage[135] ;
 wire \shift_storage.storage[1360] ;
 wire \shift_storage.storage[1361] ;
 wire \shift_storage.storage[1362] ;
 wire \shift_storage.storage[1363] ;
 wire \shift_storage.storage[1364] ;
 wire \shift_storage.storage[1365] ;
 wire \shift_storage.storage[1366] ;
 wire \shift_storage.storage[1367] ;
 wire \shift_storage.storage[1368] ;
 wire \shift_storage.storage[1369] ;
 wire \shift_storage.storage[136] ;
 wire \shift_storage.storage[1370] ;
 wire \shift_storage.storage[1371] ;
 wire \shift_storage.storage[1372] ;
 wire \shift_storage.storage[1373] ;
 wire \shift_storage.storage[1374] ;
 wire \shift_storage.storage[1375] ;
 wire \shift_storage.storage[1376] ;
 wire \shift_storage.storage[1377] ;
 wire \shift_storage.storage[1378] ;
 wire \shift_storage.storage[1379] ;
 wire \shift_storage.storage[137] ;
 wire \shift_storage.storage[1380] ;
 wire \shift_storage.storage[1381] ;
 wire \shift_storage.storage[1382] ;
 wire \shift_storage.storage[1383] ;
 wire \shift_storage.storage[1384] ;
 wire \shift_storage.storage[1385] ;
 wire \shift_storage.storage[1386] ;
 wire \shift_storage.storage[1387] ;
 wire \shift_storage.storage[1388] ;
 wire \shift_storage.storage[1389] ;
 wire \shift_storage.storage[138] ;
 wire \shift_storage.storage[1390] ;
 wire \shift_storage.storage[1391] ;
 wire \shift_storage.storage[1392] ;
 wire \shift_storage.storage[1393] ;
 wire \shift_storage.storage[1394] ;
 wire \shift_storage.storage[1395] ;
 wire \shift_storage.storage[1396] ;
 wire \shift_storage.storage[1397] ;
 wire \shift_storage.storage[1398] ;
 wire \shift_storage.storage[1399] ;
 wire \shift_storage.storage[139] ;
 wire \shift_storage.storage[13] ;
 wire \shift_storage.storage[1400] ;
 wire \shift_storage.storage[1401] ;
 wire \shift_storage.storage[1402] ;
 wire \shift_storage.storage[1403] ;
 wire \shift_storage.storage[1404] ;
 wire \shift_storage.storage[1405] ;
 wire \shift_storage.storage[1406] ;
 wire \shift_storage.storage[1407] ;
 wire \shift_storage.storage[1408] ;
 wire \shift_storage.storage[1409] ;
 wire \shift_storage.storage[140] ;
 wire \shift_storage.storage[1410] ;
 wire \shift_storage.storage[1411] ;
 wire \shift_storage.storage[1412] ;
 wire \shift_storage.storage[1413] ;
 wire \shift_storage.storage[1414] ;
 wire \shift_storage.storage[1415] ;
 wire \shift_storage.storage[1416] ;
 wire \shift_storage.storage[1417] ;
 wire \shift_storage.storage[1418] ;
 wire \shift_storage.storage[1419] ;
 wire \shift_storage.storage[141] ;
 wire \shift_storage.storage[1420] ;
 wire \shift_storage.storage[1421] ;
 wire \shift_storage.storage[1422] ;
 wire \shift_storage.storage[1423] ;
 wire \shift_storage.storage[1424] ;
 wire \shift_storage.storage[1425] ;
 wire \shift_storage.storage[1426] ;
 wire \shift_storage.storage[1427] ;
 wire \shift_storage.storage[1428] ;
 wire \shift_storage.storage[1429] ;
 wire \shift_storage.storage[142] ;
 wire \shift_storage.storage[1430] ;
 wire \shift_storage.storage[1431] ;
 wire \shift_storage.storage[1432] ;
 wire \shift_storage.storage[1433] ;
 wire \shift_storage.storage[1434] ;
 wire \shift_storage.storage[1435] ;
 wire \shift_storage.storage[1436] ;
 wire \shift_storage.storage[1437] ;
 wire \shift_storage.storage[1438] ;
 wire \shift_storage.storage[1439] ;
 wire \shift_storage.storage[143] ;
 wire \shift_storage.storage[1440] ;
 wire \shift_storage.storage[1441] ;
 wire \shift_storage.storage[1442] ;
 wire \shift_storage.storage[1443] ;
 wire \shift_storage.storage[1444] ;
 wire \shift_storage.storage[1445] ;
 wire \shift_storage.storage[1446] ;
 wire \shift_storage.storage[1447] ;
 wire \shift_storage.storage[1448] ;
 wire \shift_storage.storage[1449] ;
 wire \shift_storage.storage[144] ;
 wire \shift_storage.storage[1450] ;
 wire \shift_storage.storage[1451] ;
 wire \shift_storage.storage[1452] ;
 wire \shift_storage.storage[1453] ;
 wire \shift_storage.storage[1454] ;
 wire \shift_storage.storage[1455] ;
 wire \shift_storage.storage[1456] ;
 wire \shift_storage.storage[1457] ;
 wire \shift_storage.storage[1458] ;
 wire \shift_storage.storage[1459] ;
 wire \shift_storage.storage[145] ;
 wire \shift_storage.storage[1460] ;
 wire \shift_storage.storage[1461] ;
 wire \shift_storage.storage[1462] ;
 wire \shift_storage.storage[1463] ;
 wire \shift_storage.storage[1464] ;
 wire \shift_storage.storage[1465] ;
 wire \shift_storage.storage[1466] ;
 wire \shift_storage.storage[1467] ;
 wire \shift_storage.storage[1468] ;
 wire \shift_storage.storage[1469] ;
 wire \shift_storage.storage[146] ;
 wire \shift_storage.storage[1470] ;
 wire \shift_storage.storage[1471] ;
 wire \shift_storage.storage[1472] ;
 wire \shift_storage.storage[1473] ;
 wire \shift_storage.storage[1474] ;
 wire \shift_storage.storage[1475] ;
 wire \shift_storage.storage[1476] ;
 wire \shift_storage.storage[1477] ;
 wire \shift_storage.storage[1478] ;
 wire \shift_storage.storage[1479] ;
 wire \shift_storage.storage[147] ;
 wire \shift_storage.storage[1480] ;
 wire \shift_storage.storage[1481] ;
 wire \shift_storage.storage[1482] ;
 wire \shift_storage.storage[1483] ;
 wire \shift_storage.storage[1484] ;
 wire \shift_storage.storage[1485] ;
 wire \shift_storage.storage[1486] ;
 wire \shift_storage.storage[1487] ;
 wire \shift_storage.storage[1488] ;
 wire \shift_storage.storage[1489] ;
 wire \shift_storage.storage[148] ;
 wire \shift_storage.storage[1490] ;
 wire \shift_storage.storage[1491] ;
 wire \shift_storage.storage[1492] ;
 wire \shift_storage.storage[1493] ;
 wire \shift_storage.storage[1494] ;
 wire \shift_storage.storage[1495] ;
 wire \shift_storage.storage[1496] ;
 wire \shift_storage.storage[1497] ;
 wire \shift_storage.storage[1498] ;
 wire \shift_storage.storage[1499] ;
 wire \shift_storage.storage[149] ;
 wire \shift_storage.storage[14] ;
 wire \shift_storage.storage[1500] ;
 wire \shift_storage.storage[1501] ;
 wire \shift_storage.storage[1502] ;
 wire \shift_storage.storage[1503] ;
 wire \shift_storage.storage[1504] ;
 wire \shift_storage.storage[1505] ;
 wire \shift_storage.storage[1506] ;
 wire \shift_storage.storage[1507] ;
 wire \shift_storage.storage[1508] ;
 wire \shift_storage.storage[1509] ;
 wire \shift_storage.storage[150] ;
 wire \shift_storage.storage[1510] ;
 wire \shift_storage.storage[1511] ;
 wire \shift_storage.storage[1512] ;
 wire \shift_storage.storage[1513] ;
 wire \shift_storage.storage[1514] ;
 wire \shift_storage.storage[1515] ;
 wire \shift_storage.storage[1516] ;
 wire \shift_storage.storage[1517] ;
 wire \shift_storage.storage[1518] ;
 wire \shift_storage.storage[1519] ;
 wire \shift_storage.storage[151] ;
 wire \shift_storage.storage[1520] ;
 wire \shift_storage.storage[1521] ;
 wire \shift_storage.storage[1522] ;
 wire \shift_storage.storage[1523] ;
 wire \shift_storage.storage[1524] ;
 wire \shift_storage.storage[1525] ;
 wire \shift_storage.storage[1526] ;
 wire \shift_storage.storage[1527] ;
 wire \shift_storage.storage[1528] ;
 wire \shift_storage.storage[1529] ;
 wire \shift_storage.storage[152] ;
 wire \shift_storage.storage[1530] ;
 wire \shift_storage.storage[1531] ;
 wire \shift_storage.storage[1532] ;
 wire \shift_storage.storage[1533] ;
 wire \shift_storage.storage[1534] ;
 wire \shift_storage.storage[1535] ;
 wire \shift_storage.storage[1536] ;
 wire \shift_storage.storage[1537] ;
 wire \shift_storage.storage[1538] ;
 wire \shift_storage.storage[1539] ;
 wire \shift_storage.storage[153] ;
 wire \shift_storage.storage[1540] ;
 wire \shift_storage.storage[1541] ;
 wire \shift_storage.storage[1542] ;
 wire \shift_storage.storage[1543] ;
 wire \shift_storage.storage[1544] ;
 wire \shift_storage.storage[1545] ;
 wire \shift_storage.storage[1546] ;
 wire \shift_storage.storage[1547] ;
 wire \shift_storage.storage[1548] ;
 wire \shift_storage.storage[1549] ;
 wire \shift_storage.storage[154] ;
 wire \shift_storage.storage[1550] ;
 wire \shift_storage.storage[1551] ;
 wire \shift_storage.storage[1552] ;
 wire \shift_storage.storage[1553] ;
 wire \shift_storage.storage[1554] ;
 wire \shift_storage.storage[1555] ;
 wire \shift_storage.storage[1556] ;
 wire \shift_storage.storage[1557] ;
 wire \shift_storage.storage[1558] ;
 wire \shift_storage.storage[1559] ;
 wire \shift_storage.storage[155] ;
 wire \shift_storage.storage[1560] ;
 wire \shift_storage.storage[1561] ;
 wire \shift_storage.storage[1562] ;
 wire \shift_storage.storage[1563] ;
 wire \shift_storage.storage[1564] ;
 wire \shift_storage.storage[1565] ;
 wire \shift_storage.storage[1566] ;
 wire \shift_storage.storage[1567] ;
 wire \shift_storage.storage[1568] ;
 wire \shift_storage.storage[1569] ;
 wire \shift_storage.storage[156] ;
 wire \shift_storage.storage[1570] ;
 wire \shift_storage.storage[1571] ;
 wire \shift_storage.storage[1572] ;
 wire \shift_storage.storage[1573] ;
 wire \shift_storage.storage[1574] ;
 wire \shift_storage.storage[1575] ;
 wire \shift_storage.storage[1576] ;
 wire \shift_storage.storage[1577] ;
 wire \shift_storage.storage[1578] ;
 wire \shift_storage.storage[1579] ;
 wire \shift_storage.storage[157] ;
 wire \shift_storage.storage[1580] ;
 wire \shift_storage.storage[1581] ;
 wire \shift_storage.storage[1582] ;
 wire \shift_storage.storage[1583] ;
 wire \shift_storage.storage[1584] ;
 wire \shift_storage.storage[1585] ;
 wire \shift_storage.storage[1586] ;
 wire \shift_storage.storage[1587] ;
 wire \shift_storage.storage[1588] ;
 wire \shift_storage.storage[1589] ;
 wire \shift_storage.storage[158] ;
 wire \shift_storage.storage[1590] ;
 wire \shift_storage.storage[1591] ;
 wire \shift_storage.storage[1592] ;
 wire \shift_storage.storage[1593] ;
 wire \shift_storage.storage[1594] ;
 wire \shift_storage.storage[1595] ;
 wire \shift_storage.storage[1596] ;
 wire \shift_storage.storage[1597] ;
 wire \shift_storage.storage[1598] ;
 wire \shift_storage.storage[159] ;
 wire \shift_storage.storage[15] ;
 wire \shift_storage.storage[160] ;
 wire \shift_storage.storage[161] ;
 wire \shift_storage.storage[162] ;
 wire \shift_storage.storage[163] ;
 wire \shift_storage.storage[164] ;
 wire \shift_storage.storage[165] ;
 wire \shift_storage.storage[166] ;
 wire \shift_storage.storage[167] ;
 wire \shift_storage.storage[168] ;
 wire \shift_storage.storage[169] ;
 wire \shift_storage.storage[16] ;
 wire \shift_storage.storage[170] ;
 wire \shift_storage.storage[171] ;
 wire \shift_storage.storage[172] ;
 wire \shift_storage.storage[173] ;
 wire \shift_storage.storage[174] ;
 wire \shift_storage.storage[175] ;
 wire \shift_storage.storage[176] ;
 wire \shift_storage.storage[177] ;
 wire \shift_storage.storage[178] ;
 wire \shift_storage.storage[179] ;
 wire \shift_storage.storage[17] ;
 wire \shift_storage.storage[180] ;
 wire \shift_storage.storage[181] ;
 wire \shift_storage.storage[182] ;
 wire \shift_storage.storage[183] ;
 wire \shift_storage.storage[184] ;
 wire \shift_storage.storage[185] ;
 wire \shift_storage.storage[186] ;
 wire \shift_storage.storage[187] ;
 wire \shift_storage.storage[188] ;
 wire \shift_storage.storage[189] ;
 wire \shift_storage.storage[18] ;
 wire \shift_storage.storage[190] ;
 wire \shift_storage.storage[191] ;
 wire \shift_storage.storage[192] ;
 wire \shift_storage.storage[193] ;
 wire \shift_storage.storage[194] ;
 wire \shift_storage.storage[195] ;
 wire \shift_storage.storage[196] ;
 wire \shift_storage.storage[197] ;
 wire \shift_storage.storage[198] ;
 wire \shift_storage.storage[199] ;
 wire \shift_storage.storage[19] ;
 wire \shift_storage.storage[1] ;
 wire \shift_storage.storage[200] ;
 wire \shift_storage.storage[201] ;
 wire \shift_storage.storage[202] ;
 wire \shift_storage.storage[203] ;
 wire \shift_storage.storage[204] ;
 wire \shift_storage.storage[205] ;
 wire \shift_storage.storage[206] ;
 wire \shift_storage.storage[207] ;
 wire \shift_storage.storage[208] ;
 wire \shift_storage.storage[209] ;
 wire \shift_storage.storage[20] ;
 wire \shift_storage.storage[210] ;
 wire \shift_storage.storage[211] ;
 wire \shift_storage.storage[212] ;
 wire \shift_storage.storage[213] ;
 wire \shift_storage.storage[214] ;
 wire \shift_storage.storage[215] ;
 wire \shift_storage.storage[216] ;
 wire \shift_storage.storage[217] ;
 wire \shift_storage.storage[218] ;
 wire \shift_storage.storage[219] ;
 wire \shift_storage.storage[21] ;
 wire \shift_storage.storage[220] ;
 wire \shift_storage.storage[221] ;
 wire \shift_storage.storage[222] ;
 wire \shift_storage.storage[223] ;
 wire \shift_storage.storage[224] ;
 wire \shift_storage.storage[225] ;
 wire \shift_storage.storage[226] ;
 wire \shift_storage.storage[227] ;
 wire \shift_storage.storage[228] ;
 wire \shift_storage.storage[229] ;
 wire \shift_storage.storage[22] ;
 wire \shift_storage.storage[230] ;
 wire \shift_storage.storage[231] ;
 wire \shift_storage.storage[232] ;
 wire \shift_storage.storage[233] ;
 wire \shift_storage.storage[234] ;
 wire \shift_storage.storage[235] ;
 wire \shift_storage.storage[236] ;
 wire \shift_storage.storage[237] ;
 wire \shift_storage.storage[238] ;
 wire \shift_storage.storage[239] ;
 wire \shift_storage.storage[23] ;
 wire \shift_storage.storage[240] ;
 wire \shift_storage.storage[241] ;
 wire \shift_storage.storage[242] ;
 wire \shift_storage.storage[243] ;
 wire \shift_storage.storage[244] ;
 wire \shift_storage.storage[245] ;
 wire \shift_storage.storage[246] ;
 wire \shift_storage.storage[247] ;
 wire \shift_storage.storage[248] ;
 wire \shift_storage.storage[249] ;
 wire \shift_storage.storage[24] ;
 wire \shift_storage.storage[250] ;
 wire \shift_storage.storage[251] ;
 wire \shift_storage.storage[252] ;
 wire \shift_storage.storage[253] ;
 wire \shift_storage.storage[254] ;
 wire \shift_storage.storage[255] ;
 wire \shift_storage.storage[256] ;
 wire \shift_storage.storage[257] ;
 wire \shift_storage.storage[258] ;
 wire \shift_storage.storage[259] ;
 wire \shift_storage.storage[25] ;
 wire \shift_storage.storage[260] ;
 wire \shift_storage.storage[261] ;
 wire \shift_storage.storage[262] ;
 wire \shift_storage.storage[263] ;
 wire \shift_storage.storage[264] ;
 wire \shift_storage.storage[265] ;
 wire \shift_storage.storage[266] ;
 wire \shift_storage.storage[267] ;
 wire \shift_storage.storage[268] ;
 wire \shift_storage.storage[269] ;
 wire \shift_storage.storage[26] ;
 wire \shift_storage.storage[270] ;
 wire \shift_storage.storage[271] ;
 wire \shift_storage.storage[272] ;
 wire \shift_storage.storage[273] ;
 wire \shift_storage.storage[274] ;
 wire \shift_storage.storage[275] ;
 wire \shift_storage.storage[276] ;
 wire \shift_storage.storage[277] ;
 wire \shift_storage.storage[278] ;
 wire \shift_storage.storage[279] ;
 wire \shift_storage.storage[27] ;
 wire \shift_storage.storage[280] ;
 wire \shift_storage.storage[281] ;
 wire \shift_storage.storage[282] ;
 wire \shift_storage.storage[283] ;
 wire \shift_storage.storage[284] ;
 wire \shift_storage.storage[285] ;
 wire \shift_storage.storage[286] ;
 wire \shift_storage.storage[287] ;
 wire \shift_storage.storage[288] ;
 wire \shift_storage.storage[289] ;
 wire \shift_storage.storage[28] ;
 wire \shift_storage.storage[290] ;
 wire \shift_storage.storage[291] ;
 wire \shift_storage.storage[292] ;
 wire \shift_storage.storage[293] ;
 wire \shift_storage.storage[294] ;
 wire \shift_storage.storage[295] ;
 wire \shift_storage.storage[296] ;
 wire \shift_storage.storage[297] ;
 wire \shift_storage.storage[298] ;
 wire \shift_storage.storage[299] ;
 wire \shift_storage.storage[29] ;
 wire \shift_storage.storage[2] ;
 wire \shift_storage.storage[300] ;
 wire \shift_storage.storage[301] ;
 wire \shift_storage.storage[302] ;
 wire \shift_storage.storage[303] ;
 wire \shift_storage.storage[304] ;
 wire \shift_storage.storage[305] ;
 wire \shift_storage.storage[306] ;
 wire \shift_storage.storage[307] ;
 wire \shift_storage.storage[308] ;
 wire \shift_storage.storage[309] ;
 wire \shift_storage.storage[30] ;
 wire \shift_storage.storage[310] ;
 wire \shift_storage.storage[311] ;
 wire \shift_storage.storage[312] ;
 wire \shift_storage.storage[313] ;
 wire \shift_storage.storage[314] ;
 wire \shift_storage.storage[315] ;
 wire \shift_storage.storage[316] ;
 wire \shift_storage.storage[317] ;
 wire \shift_storage.storage[318] ;
 wire \shift_storage.storage[319] ;
 wire \shift_storage.storage[31] ;
 wire \shift_storage.storage[320] ;
 wire \shift_storage.storage[321] ;
 wire \shift_storage.storage[322] ;
 wire \shift_storage.storage[323] ;
 wire \shift_storage.storage[324] ;
 wire \shift_storage.storage[325] ;
 wire \shift_storage.storage[326] ;
 wire \shift_storage.storage[327] ;
 wire \shift_storage.storage[328] ;
 wire \shift_storage.storage[329] ;
 wire \shift_storage.storage[32] ;
 wire \shift_storage.storage[330] ;
 wire \shift_storage.storage[331] ;
 wire \shift_storage.storage[332] ;
 wire \shift_storage.storage[333] ;
 wire \shift_storage.storage[334] ;
 wire \shift_storage.storage[335] ;
 wire \shift_storage.storage[336] ;
 wire \shift_storage.storage[337] ;
 wire \shift_storage.storage[338] ;
 wire \shift_storage.storage[339] ;
 wire \shift_storage.storage[33] ;
 wire \shift_storage.storage[340] ;
 wire \shift_storage.storage[341] ;
 wire \shift_storage.storage[342] ;
 wire \shift_storage.storage[343] ;
 wire \shift_storage.storage[344] ;
 wire \shift_storage.storage[345] ;
 wire \shift_storage.storage[346] ;
 wire \shift_storage.storage[347] ;
 wire \shift_storage.storage[348] ;
 wire \shift_storage.storage[349] ;
 wire \shift_storage.storage[34] ;
 wire \shift_storage.storage[350] ;
 wire \shift_storage.storage[351] ;
 wire \shift_storage.storage[352] ;
 wire \shift_storage.storage[353] ;
 wire \shift_storage.storage[354] ;
 wire \shift_storage.storage[355] ;
 wire \shift_storage.storage[356] ;
 wire \shift_storage.storage[357] ;
 wire \shift_storage.storage[358] ;
 wire \shift_storage.storage[359] ;
 wire \shift_storage.storage[35] ;
 wire \shift_storage.storage[360] ;
 wire \shift_storage.storage[361] ;
 wire \shift_storage.storage[362] ;
 wire \shift_storage.storage[363] ;
 wire \shift_storage.storage[364] ;
 wire \shift_storage.storage[365] ;
 wire \shift_storage.storage[366] ;
 wire \shift_storage.storage[367] ;
 wire \shift_storage.storage[368] ;
 wire \shift_storage.storage[369] ;
 wire \shift_storage.storage[36] ;
 wire \shift_storage.storage[370] ;
 wire \shift_storage.storage[371] ;
 wire \shift_storage.storage[372] ;
 wire \shift_storage.storage[373] ;
 wire \shift_storage.storage[374] ;
 wire \shift_storage.storage[375] ;
 wire \shift_storage.storage[376] ;
 wire \shift_storage.storage[377] ;
 wire \shift_storage.storage[378] ;
 wire \shift_storage.storage[379] ;
 wire \shift_storage.storage[37] ;
 wire \shift_storage.storage[380] ;
 wire \shift_storage.storage[381] ;
 wire \shift_storage.storage[382] ;
 wire \shift_storage.storage[383] ;
 wire \shift_storage.storage[384] ;
 wire \shift_storage.storage[385] ;
 wire \shift_storage.storage[386] ;
 wire \shift_storage.storage[387] ;
 wire \shift_storage.storage[388] ;
 wire \shift_storage.storage[389] ;
 wire \shift_storage.storage[38] ;
 wire \shift_storage.storage[390] ;
 wire \shift_storage.storage[391] ;
 wire \shift_storage.storage[392] ;
 wire \shift_storage.storage[393] ;
 wire \shift_storage.storage[394] ;
 wire \shift_storage.storage[395] ;
 wire \shift_storage.storage[396] ;
 wire \shift_storage.storage[397] ;
 wire \shift_storage.storage[398] ;
 wire \shift_storage.storage[399] ;
 wire \shift_storage.storage[39] ;
 wire \shift_storage.storage[3] ;
 wire \shift_storage.storage[400] ;
 wire \shift_storage.storage[401] ;
 wire \shift_storage.storage[402] ;
 wire \shift_storage.storage[403] ;
 wire \shift_storage.storage[404] ;
 wire \shift_storage.storage[405] ;
 wire \shift_storage.storage[406] ;
 wire \shift_storage.storage[407] ;
 wire \shift_storage.storage[408] ;
 wire \shift_storage.storage[409] ;
 wire \shift_storage.storage[40] ;
 wire \shift_storage.storage[410] ;
 wire \shift_storage.storage[411] ;
 wire \shift_storage.storage[412] ;
 wire \shift_storage.storage[413] ;
 wire \shift_storage.storage[414] ;
 wire \shift_storage.storage[415] ;
 wire \shift_storage.storage[416] ;
 wire \shift_storage.storage[417] ;
 wire \shift_storage.storage[418] ;
 wire \shift_storage.storage[419] ;
 wire \shift_storage.storage[41] ;
 wire \shift_storage.storage[420] ;
 wire \shift_storage.storage[421] ;
 wire \shift_storage.storage[422] ;
 wire \shift_storage.storage[423] ;
 wire \shift_storage.storage[424] ;
 wire \shift_storage.storage[425] ;
 wire \shift_storage.storage[426] ;
 wire \shift_storage.storage[427] ;
 wire \shift_storage.storage[428] ;
 wire \shift_storage.storage[429] ;
 wire \shift_storage.storage[42] ;
 wire \shift_storage.storage[430] ;
 wire \shift_storage.storage[431] ;
 wire \shift_storage.storage[432] ;
 wire \shift_storage.storage[433] ;
 wire \shift_storage.storage[434] ;
 wire \shift_storage.storage[435] ;
 wire \shift_storage.storage[436] ;
 wire \shift_storage.storage[437] ;
 wire \shift_storage.storage[438] ;
 wire \shift_storage.storage[439] ;
 wire \shift_storage.storage[43] ;
 wire \shift_storage.storage[440] ;
 wire \shift_storage.storage[441] ;
 wire \shift_storage.storage[442] ;
 wire \shift_storage.storage[443] ;
 wire \shift_storage.storage[444] ;
 wire \shift_storage.storage[445] ;
 wire \shift_storage.storage[446] ;
 wire \shift_storage.storage[447] ;
 wire \shift_storage.storage[448] ;
 wire \shift_storage.storage[449] ;
 wire \shift_storage.storage[44] ;
 wire \shift_storage.storage[450] ;
 wire \shift_storage.storage[451] ;
 wire \shift_storage.storage[452] ;
 wire \shift_storage.storage[453] ;
 wire \shift_storage.storage[454] ;
 wire \shift_storage.storage[455] ;
 wire \shift_storage.storage[456] ;
 wire \shift_storage.storage[457] ;
 wire \shift_storage.storage[458] ;
 wire \shift_storage.storage[459] ;
 wire \shift_storage.storage[45] ;
 wire \shift_storage.storage[460] ;
 wire \shift_storage.storage[461] ;
 wire \shift_storage.storage[462] ;
 wire \shift_storage.storage[463] ;
 wire \shift_storage.storage[464] ;
 wire \shift_storage.storage[465] ;
 wire \shift_storage.storage[466] ;
 wire \shift_storage.storage[467] ;
 wire \shift_storage.storage[468] ;
 wire \shift_storage.storage[469] ;
 wire \shift_storage.storage[46] ;
 wire \shift_storage.storage[470] ;
 wire \shift_storage.storage[471] ;
 wire \shift_storage.storage[472] ;
 wire \shift_storage.storage[473] ;
 wire \shift_storage.storage[474] ;
 wire \shift_storage.storage[475] ;
 wire \shift_storage.storage[476] ;
 wire \shift_storage.storage[477] ;
 wire \shift_storage.storage[478] ;
 wire \shift_storage.storage[479] ;
 wire \shift_storage.storage[47] ;
 wire \shift_storage.storage[480] ;
 wire \shift_storage.storage[481] ;
 wire \shift_storage.storage[482] ;
 wire \shift_storage.storage[483] ;
 wire \shift_storage.storage[484] ;
 wire \shift_storage.storage[485] ;
 wire \shift_storage.storage[486] ;
 wire \shift_storage.storage[487] ;
 wire \shift_storage.storage[488] ;
 wire \shift_storage.storage[489] ;
 wire \shift_storage.storage[48] ;
 wire \shift_storage.storage[490] ;
 wire \shift_storage.storage[491] ;
 wire \shift_storage.storage[492] ;
 wire \shift_storage.storage[493] ;
 wire \shift_storage.storage[494] ;
 wire \shift_storage.storage[495] ;
 wire \shift_storage.storage[496] ;
 wire \shift_storage.storage[497] ;
 wire \shift_storage.storage[498] ;
 wire \shift_storage.storage[499] ;
 wire \shift_storage.storage[49] ;
 wire \shift_storage.storage[4] ;
 wire \shift_storage.storage[500] ;
 wire \shift_storage.storage[501] ;
 wire \shift_storage.storage[502] ;
 wire \shift_storage.storage[503] ;
 wire \shift_storage.storage[504] ;
 wire \shift_storage.storage[505] ;
 wire \shift_storage.storage[506] ;
 wire \shift_storage.storage[507] ;
 wire \shift_storage.storage[508] ;
 wire \shift_storage.storage[509] ;
 wire \shift_storage.storage[50] ;
 wire \shift_storage.storage[510] ;
 wire \shift_storage.storage[511] ;
 wire \shift_storage.storage[512] ;
 wire \shift_storage.storage[513] ;
 wire \shift_storage.storage[514] ;
 wire \shift_storage.storage[515] ;
 wire \shift_storage.storage[516] ;
 wire \shift_storage.storage[517] ;
 wire \shift_storage.storage[518] ;
 wire \shift_storage.storage[519] ;
 wire \shift_storage.storage[51] ;
 wire \shift_storage.storage[520] ;
 wire \shift_storage.storage[521] ;
 wire \shift_storage.storage[522] ;
 wire \shift_storage.storage[523] ;
 wire \shift_storage.storage[524] ;
 wire \shift_storage.storage[525] ;
 wire \shift_storage.storage[526] ;
 wire \shift_storage.storage[527] ;
 wire \shift_storage.storage[528] ;
 wire \shift_storage.storage[529] ;
 wire \shift_storage.storage[52] ;
 wire \shift_storage.storage[530] ;
 wire \shift_storage.storage[531] ;
 wire \shift_storage.storage[532] ;
 wire \shift_storage.storage[533] ;
 wire \shift_storage.storage[534] ;
 wire \shift_storage.storage[535] ;
 wire \shift_storage.storage[536] ;
 wire \shift_storage.storage[537] ;
 wire \shift_storage.storage[538] ;
 wire \shift_storage.storage[539] ;
 wire \shift_storage.storage[53] ;
 wire \shift_storage.storage[540] ;
 wire \shift_storage.storage[541] ;
 wire \shift_storage.storage[542] ;
 wire \shift_storage.storage[543] ;
 wire \shift_storage.storage[544] ;
 wire \shift_storage.storage[545] ;
 wire \shift_storage.storage[546] ;
 wire \shift_storage.storage[547] ;
 wire \shift_storage.storage[548] ;
 wire \shift_storage.storage[549] ;
 wire \shift_storage.storage[54] ;
 wire \shift_storage.storage[550] ;
 wire \shift_storage.storage[551] ;
 wire \shift_storage.storage[552] ;
 wire \shift_storage.storage[553] ;
 wire \shift_storage.storage[554] ;
 wire \shift_storage.storage[555] ;
 wire \shift_storage.storage[556] ;
 wire \shift_storage.storage[557] ;
 wire \shift_storage.storage[558] ;
 wire \shift_storage.storage[559] ;
 wire \shift_storage.storage[55] ;
 wire \shift_storage.storage[560] ;
 wire \shift_storage.storage[561] ;
 wire \shift_storage.storage[562] ;
 wire \shift_storage.storage[563] ;
 wire \shift_storage.storage[564] ;
 wire \shift_storage.storage[565] ;
 wire \shift_storage.storage[566] ;
 wire \shift_storage.storage[567] ;
 wire \shift_storage.storage[568] ;
 wire \shift_storage.storage[569] ;
 wire \shift_storage.storage[56] ;
 wire \shift_storage.storage[570] ;
 wire \shift_storage.storage[571] ;
 wire \shift_storage.storage[572] ;
 wire \shift_storage.storage[573] ;
 wire \shift_storage.storage[574] ;
 wire \shift_storage.storage[575] ;
 wire \shift_storage.storage[576] ;
 wire \shift_storage.storage[577] ;
 wire \shift_storage.storage[578] ;
 wire \shift_storage.storage[579] ;
 wire \shift_storage.storage[57] ;
 wire \shift_storage.storage[580] ;
 wire \shift_storage.storage[581] ;
 wire \shift_storage.storage[582] ;
 wire \shift_storage.storage[583] ;
 wire \shift_storage.storage[584] ;
 wire \shift_storage.storage[585] ;
 wire \shift_storage.storage[586] ;
 wire \shift_storage.storage[587] ;
 wire \shift_storage.storage[588] ;
 wire \shift_storage.storage[589] ;
 wire \shift_storage.storage[58] ;
 wire \shift_storage.storage[590] ;
 wire \shift_storage.storage[591] ;
 wire \shift_storage.storage[592] ;
 wire \shift_storage.storage[593] ;
 wire \shift_storage.storage[594] ;
 wire \shift_storage.storage[595] ;
 wire \shift_storage.storage[596] ;
 wire \shift_storage.storage[597] ;
 wire \shift_storage.storage[598] ;
 wire \shift_storage.storage[599] ;
 wire \shift_storage.storage[59] ;
 wire \shift_storage.storage[5] ;
 wire \shift_storage.storage[600] ;
 wire \shift_storage.storage[601] ;
 wire \shift_storage.storage[602] ;
 wire \shift_storage.storage[603] ;
 wire \shift_storage.storage[604] ;
 wire \shift_storage.storage[605] ;
 wire \shift_storage.storage[606] ;
 wire \shift_storage.storage[607] ;
 wire \shift_storage.storage[608] ;
 wire \shift_storage.storage[609] ;
 wire \shift_storage.storage[60] ;
 wire \shift_storage.storage[610] ;
 wire \shift_storage.storage[611] ;
 wire \shift_storage.storage[612] ;
 wire \shift_storage.storage[613] ;
 wire \shift_storage.storage[614] ;
 wire \shift_storage.storage[615] ;
 wire \shift_storage.storage[616] ;
 wire \shift_storage.storage[617] ;
 wire \shift_storage.storage[618] ;
 wire \shift_storage.storage[619] ;
 wire \shift_storage.storage[61] ;
 wire \shift_storage.storage[620] ;
 wire \shift_storage.storage[621] ;
 wire \shift_storage.storage[622] ;
 wire \shift_storage.storage[623] ;
 wire \shift_storage.storage[624] ;
 wire \shift_storage.storage[625] ;
 wire \shift_storage.storage[626] ;
 wire \shift_storage.storage[627] ;
 wire \shift_storage.storage[628] ;
 wire \shift_storage.storage[629] ;
 wire \shift_storage.storage[62] ;
 wire \shift_storage.storage[630] ;
 wire \shift_storage.storage[631] ;
 wire \shift_storage.storage[632] ;
 wire \shift_storage.storage[633] ;
 wire \shift_storage.storage[634] ;
 wire \shift_storage.storage[635] ;
 wire \shift_storage.storage[636] ;
 wire \shift_storage.storage[637] ;
 wire \shift_storage.storage[638] ;
 wire \shift_storage.storage[639] ;
 wire \shift_storage.storage[63] ;
 wire \shift_storage.storage[640] ;
 wire \shift_storage.storage[641] ;
 wire \shift_storage.storage[642] ;
 wire \shift_storage.storage[643] ;
 wire \shift_storage.storage[644] ;
 wire \shift_storage.storage[645] ;
 wire \shift_storage.storage[646] ;
 wire \shift_storage.storage[647] ;
 wire \shift_storage.storage[648] ;
 wire \shift_storage.storage[649] ;
 wire \shift_storage.storage[64] ;
 wire \shift_storage.storage[650] ;
 wire \shift_storage.storage[651] ;
 wire \shift_storage.storage[652] ;
 wire \shift_storage.storage[653] ;
 wire \shift_storage.storage[654] ;
 wire \shift_storage.storage[655] ;
 wire \shift_storage.storage[656] ;
 wire \shift_storage.storage[657] ;
 wire \shift_storage.storage[658] ;
 wire \shift_storage.storage[659] ;
 wire \shift_storage.storage[65] ;
 wire \shift_storage.storage[660] ;
 wire \shift_storage.storage[661] ;
 wire \shift_storage.storage[662] ;
 wire \shift_storage.storage[663] ;
 wire \shift_storage.storage[664] ;
 wire \shift_storage.storage[665] ;
 wire \shift_storage.storage[666] ;
 wire \shift_storage.storage[667] ;
 wire \shift_storage.storage[668] ;
 wire \shift_storage.storage[669] ;
 wire \shift_storage.storage[66] ;
 wire \shift_storage.storage[670] ;
 wire \shift_storage.storage[671] ;
 wire \shift_storage.storage[672] ;
 wire \shift_storage.storage[673] ;
 wire \shift_storage.storage[674] ;
 wire \shift_storage.storage[675] ;
 wire \shift_storage.storage[676] ;
 wire \shift_storage.storage[677] ;
 wire \shift_storage.storage[678] ;
 wire \shift_storage.storage[679] ;
 wire \shift_storage.storage[67] ;
 wire \shift_storage.storage[680] ;
 wire \shift_storage.storage[681] ;
 wire \shift_storage.storage[682] ;
 wire \shift_storage.storage[683] ;
 wire \shift_storage.storage[684] ;
 wire \shift_storage.storage[685] ;
 wire \shift_storage.storage[686] ;
 wire \shift_storage.storage[687] ;
 wire \shift_storage.storage[688] ;
 wire \shift_storage.storage[689] ;
 wire \shift_storage.storage[68] ;
 wire \shift_storage.storage[690] ;
 wire \shift_storage.storage[691] ;
 wire \shift_storage.storage[692] ;
 wire \shift_storage.storage[693] ;
 wire \shift_storage.storage[694] ;
 wire \shift_storage.storage[695] ;
 wire \shift_storage.storage[696] ;
 wire \shift_storage.storage[697] ;
 wire \shift_storage.storage[698] ;
 wire \shift_storage.storage[699] ;
 wire \shift_storage.storage[69] ;
 wire \shift_storage.storage[6] ;
 wire \shift_storage.storage[700] ;
 wire \shift_storage.storage[701] ;
 wire \shift_storage.storage[702] ;
 wire \shift_storage.storage[703] ;
 wire \shift_storage.storage[704] ;
 wire \shift_storage.storage[705] ;
 wire \shift_storage.storage[706] ;
 wire \shift_storage.storage[707] ;
 wire \shift_storage.storage[708] ;
 wire \shift_storage.storage[709] ;
 wire \shift_storage.storage[70] ;
 wire \shift_storage.storage[710] ;
 wire \shift_storage.storage[711] ;
 wire \shift_storage.storage[712] ;
 wire \shift_storage.storage[713] ;
 wire \shift_storage.storage[714] ;
 wire \shift_storage.storage[715] ;
 wire \shift_storage.storage[716] ;
 wire \shift_storage.storage[717] ;
 wire \shift_storage.storage[718] ;
 wire \shift_storage.storage[719] ;
 wire \shift_storage.storage[71] ;
 wire \shift_storage.storage[720] ;
 wire \shift_storage.storage[721] ;
 wire \shift_storage.storage[722] ;
 wire \shift_storage.storage[723] ;
 wire \shift_storage.storage[724] ;
 wire \shift_storage.storage[725] ;
 wire \shift_storage.storage[726] ;
 wire \shift_storage.storage[727] ;
 wire \shift_storage.storage[728] ;
 wire \shift_storage.storage[729] ;
 wire \shift_storage.storage[72] ;
 wire \shift_storage.storage[730] ;
 wire \shift_storage.storage[731] ;
 wire \shift_storage.storage[732] ;
 wire \shift_storage.storage[733] ;
 wire \shift_storage.storage[734] ;
 wire \shift_storage.storage[735] ;
 wire \shift_storage.storage[736] ;
 wire \shift_storage.storage[737] ;
 wire \shift_storage.storage[738] ;
 wire \shift_storage.storage[739] ;
 wire \shift_storage.storage[73] ;
 wire \shift_storage.storage[740] ;
 wire \shift_storage.storage[741] ;
 wire \shift_storage.storage[742] ;
 wire \shift_storage.storage[743] ;
 wire \shift_storage.storage[744] ;
 wire \shift_storage.storage[745] ;
 wire \shift_storage.storage[746] ;
 wire \shift_storage.storage[747] ;
 wire \shift_storage.storage[748] ;
 wire \shift_storage.storage[749] ;
 wire \shift_storage.storage[74] ;
 wire \shift_storage.storage[750] ;
 wire \shift_storage.storage[751] ;
 wire \shift_storage.storage[752] ;
 wire \shift_storage.storage[753] ;
 wire \shift_storage.storage[754] ;
 wire \shift_storage.storage[755] ;
 wire \shift_storage.storage[756] ;
 wire \shift_storage.storage[757] ;
 wire \shift_storage.storage[758] ;
 wire \shift_storage.storage[759] ;
 wire \shift_storage.storage[75] ;
 wire \shift_storage.storage[760] ;
 wire \shift_storage.storage[761] ;
 wire \shift_storage.storage[762] ;
 wire \shift_storage.storage[763] ;
 wire \shift_storage.storage[764] ;
 wire \shift_storage.storage[765] ;
 wire \shift_storage.storage[766] ;
 wire \shift_storage.storage[767] ;
 wire \shift_storage.storage[768] ;
 wire \shift_storage.storage[769] ;
 wire \shift_storage.storage[76] ;
 wire \shift_storage.storage[770] ;
 wire \shift_storage.storage[771] ;
 wire \shift_storage.storage[772] ;
 wire \shift_storage.storage[773] ;
 wire \shift_storage.storage[774] ;
 wire \shift_storage.storage[775] ;
 wire \shift_storage.storage[776] ;
 wire \shift_storage.storage[777] ;
 wire \shift_storage.storage[778] ;
 wire \shift_storage.storage[779] ;
 wire \shift_storage.storage[77] ;
 wire \shift_storage.storage[780] ;
 wire \shift_storage.storage[781] ;
 wire \shift_storage.storage[782] ;
 wire \shift_storage.storage[783] ;
 wire \shift_storage.storage[784] ;
 wire \shift_storage.storage[785] ;
 wire \shift_storage.storage[786] ;
 wire \shift_storage.storage[787] ;
 wire \shift_storage.storage[788] ;
 wire \shift_storage.storage[789] ;
 wire \shift_storage.storage[78] ;
 wire \shift_storage.storage[790] ;
 wire \shift_storage.storage[791] ;
 wire \shift_storage.storage[792] ;
 wire \shift_storage.storage[793] ;
 wire \shift_storage.storage[794] ;
 wire \shift_storage.storage[795] ;
 wire \shift_storage.storage[796] ;
 wire \shift_storage.storage[797] ;
 wire \shift_storage.storage[798] ;
 wire \shift_storage.storage[799] ;
 wire \shift_storage.storage[79] ;
 wire \shift_storage.storage[7] ;
 wire \shift_storage.storage[800] ;
 wire \shift_storage.storage[801] ;
 wire \shift_storage.storage[802] ;
 wire \shift_storage.storage[803] ;
 wire \shift_storage.storage[804] ;
 wire \shift_storage.storage[805] ;
 wire \shift_storage.storage[806] ;
 wire \shift_storage.storage[807] ;
 wire \shift_storage.storage[808] ;
 wire \shift_storage.storage[809] ;
 wire \shift_storage.storage[80] ;
 wire \shift_storage.storage[810] ;
 wire \shift_storage.storage[811] ;
 wire \shift_storage.storage[812] ;
 wire \shift_storage.storage[813] ;
 wire \shift_storage.storage[814] ;
 wire \shift_storage.storage[815] ;
 wire \shift_storage.storage[816] ;
 wire \shift_storage.storage[817] ;
 wire \shift_storage.storage[818] ;
 wire \shift_storage.storage[819] ;
 wire \shift_storage.storage[81] ;
 wire \shift_storage.storage[820] ;
 wire \shift_storage.storage[821] ;
 wire \shift_storage.storage[822] ;
 wire \shift_storage.storage[823] ;
 wire \shift_storage.storage[824] ;
 wire \shift_storage.storage[825] ;
 wire \shift_storage.storage[826] ;
 wire \shift_storage.storage[827] ;
 wire \shift_storage.storage[828] ;
 wire \shift_storage.storage[829] ;
 wire \shift_storage.storage[82] ;
 wire \shift_storage.storage[830] ;
 wire \shift_storage.storage[831] ;
 wire \shift_storage.storage[832] ;
 wire \shift_storage.storage[833] ;
 wire \shift_storage.storage[834] ;
 wire \shift_storage.storage[835] ;
 wire \shift_storage.storage[836] ;
 wire \shift_storage.storage[837] ;
 wire \shift_storage.storage[838] ;
 wire \shift_storage.storage[839] ;
 wire \shift_storage.storage[83] ;
 wire \shift_storage.storage[840] ;
 wire \shift_storage.storage[841] ;
 wire \shift_storage.storage[842] ;
 wire \shift_storage.storage[843] ;
 wire \shift_storage.storage[844] ;
 wire \shift_storage.storage[845] ;
 wire \shift_storage.storage[846] ;
 wire \shift_storage.storage[847] ;
 wire \shift_storage.storage[848] ;
 wire \shift_storage.storage[849] ;
 wire \shift_storage.storage[84] ;
 wire \shift_storage.storage[850] ;
 wire \shift_storage.storage[851] ;
 wire \shift_storage.storage[852] ;
 wire \shift_storage.storage[853] ;
 wire \shift_storage.storage[854] ;
 wire \shift_storage.storage[855] ;
 wire \shift_storage.storage[856] ;
 wire \shift_storage.storage[857] ;
 wire \shift_storage.storage[858] ;
 wire \shift_storage.storage[859] ;
 wire \shift_storage.storage[85] ;
 wire \shift_storage.storage[860] ;
 wire \shift_storage.storage[861] ;
 wire \shift_storage.storage[862] ;
 wire \shift_storage.storage[863] ;
 wire \shift_storage.storage[864] ;
 wire \shift_storage.storage[865] ;
 wire \shift_storage.storage[866] ;
 wire \shift_storage.storage[867] ;
 wire \shift_storage.storage[868] ;
 wire \shift_storage.storage[869] ;
 wire \shift_storage.storage[86] ;
 wire \shift_storage.storage[870] ;
 wire \shift_storage.storage[871] ;
 wire \shift_storage.storage[872] ;
 wire \shift_storage.storage[873] ;
 wire \shift_storage.storage[874] ;
 wire \shift_storage.storage[875] ;
 wire \shift_storage.storage[876] ;
 wire \shift_storage.storage[877] ;
 wire \shift_storage.storage[878] ;
 wire \shift_storage.storage[879] ;
 wire \shift_storage.storage[87] ;
 wire \shift_storage.storage[880] ;
 wire \shift_storage.storage[881] ;
 wire \shift_storage.storage[882] ;
 wire \shift_storage.storage[883] ;
 wire \shift_storage.storage[884] ;
 wire \shift_storage.storage[885] ;
 wire \shift_storage.storage[886] ;
 wire \shift_storage.storage[887] ;
 wire \shift_storage.storage[888] ;
 wire \shift_storage.storage[889] ;
 wire \shift_storage.storage[88] ;
 wire \shift_storage.storage[890] ;
 wire \shift_storage.storage[891] ;
 wire \shift_storage.storage[892] ;
 wire \shift_storage.storage[893] ;
 wire \shift_storage.storage[894] ;
 wire \shift_storage.storage[895] ;
 wire \shift_storage.storage[896] ;
 wire \shift_storage.storage[897] ;
 wire \shift_storage.storage[898] ;
 wire \shift_storage.storage[899] ;
 wire \shift_storage.storage[89] ;
 wire \shift_storage.storage[8] ;
 wire \shift_storage.storage[900] ;
 wire \shift_storage.storage[901] ;
 wire \shift_storage.storage[902] ;
 wire \shift_storage.storage[903] ;
 wire \shift_storage.storage[904] ;
 wire \shift_storage.storage[905] ;
 wire \shift_storage.storage[906] ;
 wire \shift_storage.storage[907] ;
 wire \shift_storage.storage[908] ;
 wire \shift_storage.storage[909] ;
 wire \shift_storage.storage[90] ;
 wire \shift_storage.storage[910] ;
 wire \shift_storage.storage[911] ;
 wire \shift_storage.storage[912] ;
 wire \shift_storage.storage[913] ;
 wire \shift_storage.storage[914] ;
 wire \shift_storage.storage[915] ;
 wire \shift_storage.storage[916] ;
 wire \shift_storage.storage[917] ;
 wire \shift_storage.storage[918] ;
 wire \shift_storage.storage[919] ;
 wire \shift_storage.storage[91] ;
 wire \shift_storage.storage[920] ;
 wire \shift_storage.storage[921] ;
 wire \shift_storage.storage[922] ;
 wire \shift_storage.storage[923] ;
 wire \shift_storage.storage[924] ;
 wire \shift_storage.storage[925] ;
 wire \shift_storage.storage[926] ;
 wire \shift_storage.storage[927] ;
 wire \shift_storage.storage[928] ;
 wire \shift_storage.storage[929] ;
 wire \shift_storage.storage[92] ;
 wire \shift_storage.storage[930] ;
 wire \shift_storage.storage[931] ;
 wire \shift_storage.storage[932] ;
 wire \shift_storage.storage[933] ;
 wire \shift_storage.storage[934] ;
 wire \shift_storage.storage[935] ;
 wire \shift_storage.storage[936] ;
 wire \shift_storage.storage[937] ;
 wire \shift_storage.storage[938] ;
 wire \shift_storage.storage[939] ;
 wire \shift_storage.storage[93] ;
 wire \shift_storage.storage[940] ;
 wire \shift_storage.storage[941] ;
 wire \shift_storage.storage[942] ;
 wire \shift_storage.storage[943] ;
 wire \shift_storage.storage[944] ;
 wire \shift_storage.storage[945] ;
 wire \shift_storage.storage[946] ;
 wire \shift_storage.storage[947] ;
 wire \shift_storage.storage[948] ;
 wire \shift_storage.storage[949] ;
 wire \shift_storage.storage[94] ;
 wire \shift_storage.storage[950] ;
 wire \shift_storage.storage[951] ;
 wire \shift_storage.storage[952] ;
 wire \shift_storage.storage[953] ;
 wire \shift_storage.storage[954] ;
 wire \shift_storage.storage[955] ;
 wire \shift_storage.storage[956] ;
 wire \shift_storage.storage[957] ;
 wire \shift_storage.storage[958] ;
 wire \shift_storage.storage[959] ;
 wire \shift_storage.storage[95] ;
 wire \shift_storage.storage[960] ;
 wire \shift_storage.storage[961] ;
 wire \shift_storage.storage[962] ;
 wire \shift_storage.storage[963] ;
 wire \shift_storage.storage[964] ;
 wire \shift_storage.storage[965] ;
 wire \shift_storage.storage[966] ;
 wire \shift_storage.storage[967] ;
 wire \shift_storage.storage[968] ;
 wire \shift_storage.storage[969] ;
 wire \shift_storage.storage[96] ;
 wire \shift_storage.storage[970] ;
 wire \shift_storage.storage[971] ;
 wire \shift_storage.storage[972] ;
 wire \shift_storage.storage[973] ;
 wire \shift_storage.storage[974] ;
 wire \shift_storage.storage[975] ;
 wire \shift_storage.storage[976] ;
 wire \shift_storage.storage[977] ;
 wire \shift_storage.storage[978] ;
 wire \shift_storage.storage[979] ;
 wire \shift_storage.storage[97] ;
 wire \shift_storage.storage[980] ;
 wire \shift_storage.storage[981] ;
 wire \shift_storage.storage[982] ;
 wire \shift_storage.storage[983] ;
 wire \shift_storage.storage[984] ;
 wire \shift_storage.storage[985] ;
 wire \shift_storage.storage[986] ;
 wire \shift_storage.storage[987] ;
 wire \shift_storage.storage[988] ;
 wire \shift_storage.storage[989] ;
 wire \shift_storage.storage[98] ;
 wire \shift_storage.storage[990] ;
 wire \shift_storage.storage[991] ;
 wire \shift_storage.storage[992] ;
 wire \shift_storage.storage[993] ;
 wire \shift_storage.storage[994] ;
 wire \shift_storage.storage[995] ;
 wire \shift_storage.storage[996] ;
 wire \shift_storage.storage[997] ;
 wire \shift_storage.storage[998] ;
 wire \shift_storage.storage[999] ;
 wire \shift_storage.storage[99] ;
 wire \shift_storage.storage[9] ;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net995;
 wire net996;
 wire net997;
 wire net998;
 wire net999;
 wire net1000;
 wire net1001;
 wire net1002;
 wire net1003;
 wire net1004;
 wire net1005;
 wire net1006;
 wire net1007;
 wire net1008;
 wire net1009;
 wire net1010;
 wire net1011;
 wire net1012;
 wire net1013;
 wire net1014;
 wire net1015;
 wire net1016;
 wire net1017;
 wire net1018;
 wire net1019;
 wire net1020;
 wire net1021;
 wire net1022;
 wire net1023;
 wire net1024;
 wire net1025;
 wire net1026;
 wire net1027;
 wire net1028;
 wire net1029;
 wire net1030;
 wire net1031;
 wire net1032;
 wire net1033;
 wire net1034;
 wire net1035;
 wire net1036;
 wire net1037;
 wire net1038;
 wire net1039;
 wire net1040;
 wire net1041;
 wire net1042;
 wire net1043;
 wire net1044;
 wire net1045;
 wire net1046;
 wire net1047;
 wire net1048;
 wire net1049;
 wire net1050;
 wire net1051;
 wire net1052;
 wire net1053;
 wire net1054;
 wire net1055;
 wire net1056;
 wire net1057;
 wire net1058;
 wire net1059;
 wire net1060;
 wire net1061;
 wire net1062;
 wire net1063;
 wire net1064;
 wire net1065;
 wire net1066;
 wire net1067;
 wire net1068;
 wire net1069;
 wire net1070;
 wire net1071;
 wire net1072;
 wire net1073;
 wire net1074;
 wire net1075;
 wire net1076;
 wire net1077;
 wire net1078;
 wire net1079;
 wire net1080;
 wire net1081;
 wire net1082;
 wire net1083;
 wire net1084;
 wire net1085;
 wire net1086;
 wire net1087;
 wire net1088;
 wire net1089;
 wire net1090;
 wire net1091;
 wire net1092;
 wire net1093;
 wire net1094;
 wire net1095;
 wire net1096;
 wire net1097;
 wire net1098;
 wire net1099;
 wire net1100;
 wire net1101;
 wire net1102;
 wire net1103;
 wire net1104;
 wire net1105;
 wire net1106;
 wire net1107;
 wire net1108;
 wire net1109;
 wire net1110;
 wire net1111;
 wire net1112;
 wire net1113;
 wire net1114;
 wire net1115;
 wire net1116;
 wire net1117;
 wire net1118;
 wire net1119;
 wire net1120;
 wire net1121;
 wire net1122;
 wire net1123;
 wire net1124;
 wire net1125;
 wire net1126;
 wire net1127;
 wire net1128;
 wire net1129;
 wire net1130;
 wire net1131;
 wire net1132;
 wire net1133;
 wire net1134;
 wire net1135;
 wire net1136;
 wire net1137;
 wire net1138;
 wire net1139;
 wire net1140;
 wire net1141;
 wire net1142;
 wire net1143;
 wire net1144;
 wire net1145;
 wire net1146;
 wire net1147;
 wire net1148;
 wire net1149;
 wire net1150;
 wire net1151;
 wire net1152;
 wire net1153;
 wire net1154;
 wire net1155;
 wire net1156;
 wire net1157;
 wire net1158;
 wire net1159;
 wire net1160;
 wire net1161;
 wire net1162;
 wire net1163;
 wire net1164;
 wire net1165;
 wire net1166;
 wire net1167;
 wire net1168;
 wire net1169;
 wire net1170;
 wire net1171;
 wire net1172;
 wire net1173;
 wire net1174;
 wire net1175;
 wire net1176;
 wire net1177;
 wire net1178;
 wire net1179;
 wire net1180;
 wire net1181;
 wire net1182;
 wire net1183;
 wire net1184;
 wire net1185;
 wire net1186;
 wire net1187;
 wire net1188;
 wire net1189;
 wire net1190;
 wire net1191;
 wire net1192;
 wire net1193;
 wire net1194;
 wire net1195;
 wire net1196;
 wire net1197;
 wire net1198;
 wire net1199;
 wire net1200;
 wire net1201;
 wire net1202;
 wire net1203;
 wire net1204;
 wire net1205;
 wire net1206;
 wire net1207;
 wire net1208;
 wire net1209;
 wire net1210;
 wire net1211;
 wire net1212;
 wire net1213;
 wire net1214;
 wire net1215;
 wire net1216;
 wire net1217;
 wire net1218;
 wire net1219;
 wire net1220;
 wire net1221;
 wire net1222;
 wire net1223;
 wire net1224;
 wire net1225;
 wire net1226;
 wire net1227;
 wire net1228;
 wire net1229;
 wire net1230;
 wire net1231;
 wire net1232;
 wire net1233;
 wire net1234;
 wire net1235;
 wire net1236;
 wire net1237;
 wire net1238;
 wire net1239;
 wire net1240;
 wire net1241;
 wire net1242;
 wire net1243;
 wire net1244;
 wire net1245;
 wire net1246;
 wire net1247;
 wire net1248;
 wire net1249;
 wire net1250;
 wire net1251;
 wire net1252;
 wire net1253;
 wire net1254;
 wire net1255;
 wire net1256;
 wire net1257;
 wire net1258;
 wire net1259;
 wire net1260;
 wire net1261;
 wire net1262;
 wire net1263;
 wire net1264;
 wire net1265;
 wire net1266;
 wire net1267;
 wire net1268;
 wire net1269;
 wire net1270;
 wire net1271;
 wire net1272;
 wire net1273;
 wire net1274;
 wire net1275;
 wire net1276;
 wire net1277;
 wire net1278;
 wire net1279;
 wire net1280;
 wire net1281;
 wire net1282;
 wire net1283;
 wire net1284;
 wire net1285;
 wire net1286;
 wire net1287;
 wire net1288;
 wire net1289;
 wire net1290;
 wire net1291;
 wire net1292;
 wire net1293;
 wire net1294;
 wire net1295;
 wire net1296;
 wire net1297;
 wire net1298;
 wire net1299;
 wire net1300;
 wire net1301;
 wire net1302;
 wire net1303;
 wire net1304;
 wire net1305;
 wire net1306;
 wire net1307;
 wire net1308;
 wire net1309;
 wire net1310;
 wire net1311;
 wire net1312;
 wire net1313;
 wire net1314;
 wire net1315;
 wire net1316;
 wire net1317;
 wire net1318;
 wire net1319;
 wire net1320;
 wire net1321;
 wire net1322;
 wire net1323;
 wire net1324;
 wire net1325;
 wire net1326;
 wire net1327;
 wire net1328;
 wire net1329;
 wire net1330;
 wire net1331;
 wire net1332;
 wire net1333;
 wire net1334;
 wire net1335;
 wire net1336;
 wire net1337;
 wire net1338;
 wire net1339;
 wire net1340;
 wire net1341;
 wire net1342;
 wire net1343;
 wire net1344;
 wire net1345;
 wire net1346;
 wire net1347;
 wire net1348;
 wire net1349;
 wire net1350;
 wire net1351;
 wire net1352;
 wire net1353;
 wire net1354;
 wire net1355;
 wire net1356;
 wire net1357;
 wire net1358;
 wire net1359;
 wire net1360;
 wire net1361;
 wire net1362;
 wire net1363;
 wire net1364;
 wire net1365;
 wire net1366;
 wire net1367;
 wire net1368;
 wire net1369;
 wire net1370;
 wire net1371;
 wire net1372;
 wire net1373;
 wire net1374;
 wire net1375;
 wire net1376;
 wire net1377;
 wire net1378;
 wire net1379;
 wire net1380;
 wire net1381;
 wire net1382;
 wire net1383;
 wire net1384;
 wire net1385;
 wire net1386;
 wire net1387;
 wire net1388;
 wire net1389;
 wire net1390;
 wire net1391;
 wire net1392;
 wire net1393;
 wire net1394;
 wire net1395;
 wire net1396;
 wire net1397;
 wire net1398;
 wire net1399;
 wire net1400;
 wire net1401;
 wire net1402;
 wire net1403;
 wire net1404;
 wire net1405;
 wire net1406;
 wire net1407;
 wire net1408;
 wire net1409;
 wire net1410;
 wire net1411;
 wire net1412;
 wire net1413;
 wire net1414;
 wire net1415;
 wire net1416;
 wire net1417;
 wire net1418;
 wire net1419;
 wire net1420;
 wire net1421;
 wire net1422;
 wire net1423;
 wire net1424;
 wire net1425;
 wire net1426;
 wire net1427;
 wire net1428;
 wire net1429;
 wire net1430;
 wire net1431;
 wire net1432;
 wire net1433;
 wire net1434;
 wire net1435;
 wire net1436;
 wire net1437;
 wire net1438;
 wire net1439;
 wire net1440;
 wire net1441;
 wire net1442;
 wire net1443;
 wire net1444;
 wire net1445;
 wire net1446;
 wire net1447;
 wire net1448;
 wire net1449;
 wire net1450;
 wire net1451;
 wire net1452;
 wire net1453;
 wire net1454;
 wire net1455;
 wire net1456;
 wire net1457;
 wire net1458;
 wire net1459;
 wire net1460;
 wire net1461;
 wire net1462;
 wire net1463;
 wire net1464;
 wire net1465;
 wire net1466;
 wire net1467;
 wire net1468;
 wire net1469;
 wire net1470;
 wire net1471;
 wire net1472;
 wire net1473;
 wire net1474;
 wire net1475;
 wire net1476;
 wire net1477;
 wire net1478;
 wire net1479;
 wire net1480;
 wire net1481;
 wire net1482;
 wire net1483;
 wire net1484;
 wire net1485;
 wire net1486;
 wire net1487;
 wire net1488;
 wire net1489;
 wire net1490;
 wire net1491;
 wire net1492;
 wire net1493;
 wire net1494;
 wire net1495;
 wire net1496;
 wire net1497;
 wire net1498;
 wire net1499;
 wire net1500;
 wire net1501;
 wire net1502;
 wire net1503;
 wire net1504;
 wire net1505;
 wire net1506;
 wire net1507;
 wire net1508;
 wire net1509;
 wire net1510;
 wire net1511;
 wire net1512;
 wire net1513;
 wire net1514;
 wire net1515;
 wire net1516;
 wire net1517;
 wire net1518;
 wire net1519;
 wire net1520;
 wire net1521;
 wire net1522;
 wire net1523;
 wire net1524;
 wire net1525;
 wire net1526;
 wire net1527;
 wire net1528;
 wire net1529;
 wire net1530;
 wire net1531;
 wire net1532;
 wire net1533;
 wire net1534;
 wire net1535;
 wire net1536;
 wire net1537;
 wire net1538;
 wire net1539;
 wire net1540;
 wire net1541;
 wire net1542;
 wire net1543;
 wire net1544;
 wire net1545;
 wire net1546;
 wire net1547;
 wire net1548;
 wire net1549;
 wire net1550;
 wire net1551;
 wire net1552;
 wire net1553;
 wire net1554;
 wire net1555;
 wire net1556;
 wire net1557;
 wire net1558;
 wire net1559;
 wire net1560;
 wire net1561;
 wire net1562;
 wire net1563;
 wire net1564;
 wire net1565;
 wire net1566;
 wire net1567;
 wire net1568;
 wire net1569;
 wire net1570;
 wire net1571;
 wire net1572;
 wire net1573;
 wire net1574;
 wire net1575;
 wire net1576;
 wire net1577;
 wire net1578;
 wire net1579;
 wire net1580;
 wire net1581;
 wire net1582;
 wire net1583;
 wire net1584;
 wire net1585;
 wire net1586;
 wire net1587;
 wire net1588;
 wire net1589;
 wire net1590;
 wire net1591;
 wire net1592;
 wire net1593;
 wire net1594;
 wire net1595;
 wire net1596;
 wire net1597;
 wire net1598;
 wire net1599;
 wire net1600;
 wire net1601;
 wire net1602;
 wire net1603;
 wire net1604;
 wire net1605;
 wire net1606;
 wire net1607;
 wire net1608;
 wire net1609;
 wire net1610;
 wire net1611;
 wire net1612;
 wire net1613;
 wire net1614;
 wire net1615;
 wire net1616;
 wire net1617;
 wire net1618;
 wire net1619;
 wire net1620;
 wire net1621;
 wire net1622;
 wire net1623;
 wire net1624;
 wire net1625;
 wire net1626;
 wire net1627;
 wire net1628;
 wire net1629;
 wire net1630;
 wire net1631;
 wire net1632;
 wire net1633;
 wire net1634;
 wire net1635;
 wire net1636;
 wire net1637;
 wire net1638;
 wire net1639;
 wire net1640;
 wire net1641;
 wire net1642;
 wire net1643;
 wire net1644;
 wire net1645;
 wire net1646;
 wire net1647;
 wire net1648;
 wire net1649;
 wire net1650;
 wire net1651;
 wire net1652;
 wire net1653;
 wire net1654;
 wire net1655;
 wire net1656;
 wire net1657;
 wire net1658;
 wire net1659;
 wire net1660;
 wire net1661;
 wire net1662;
 wire net1663;
 wire net1664;
 wire net1665;
 wire net1666;
 wire net1667;
 wire net1668;
 wire net1669;
 wire net1670;
 wire net1671;
 wire net1672;
 wire net1673;
 wire net1674;
 wire net1675;
 wire net1676;
 wire net1677;
 wire net1678;
 wire net1679;
 wire net1680;
 wire net1681;
 wire net1682;
 wire net1683;
 wire net1684;
 wire net1685;
 wire net1686;
 wire net1687;
 wire net1688;
 wire net1689;
 wire net1690;
 wire net1691;
 wire net1692;
 wire net1693;
 wire net1694;
 wire net1695;
 wire net1696;
 wire net1697;
 wire net1698;
 wire net1699;
 wire net1700;
 wire net1701;
 wire net1702;
 wire net1703;
 wire net1704;
 wire net1705;
 wire net1706;
 wire net1707;
 wire net1708;
 wire net1709;
 wire net1710;
 wire net1711;
 wire net1712;
 wire net1713;
 wire net1714;
 wire net1715;
 wire net1716;
 wire net1717;
 wire net1718;
 wire net1719;
 wire net1720;
 wire net1721;
 wire net1722;
 wire net1723;
 wire net1724;
 wire net1725;
 wire net1726;
 wire net1727;
 wire net1728;
 wire net1729;
 wire net1730;
 wire net1731;
 wire net1732;
 wire net1733;
 wire net1734;
 wire net1735;
 wire net1736;
 wire net1737;
 wire net1738;
 wire net1739;
 wire net1740;
 wire net1741;
 wire net1742;
 wire net1743;
 wire net1744;
 wire net1745;
 wire net1746;
 wire net1747;
 wire net1748;
 wire net1749;
 wire net1750;
 wire net1751;
 wire net1752;
 wire net1753;
 wire net1754;
 wire net1755;
 wire net1756;
 wire net1757;
 wire net1758;
 wire net1759;
 wire net1760;
 wire net1761;
 wire net1762;
 wire net1763;
 wire net1764;
 wire net1765;
 wire net1766;
 wire net1767;
 wire net1768;
 wire net1769;
 wire net1770;
 wire net1771;
 wire net1772;
 wire net1773;
 wire net1774;
 wire net1775;
 wire net1776;
 wire net1777;
 wire net1778;
 wire net1779;
 wire net1780;
 wire net1781;
 wire net1782;
 wire net1783;
 wire net1784;
 wire net1785;
 wire net1786;
 wire net1787;
 wire net1788;
 wire net1789;
 wire net1790;
 wire net1791;
 wire net1792;
 wire net1793;
 wire net1794;
 wire net1795;
 wire net1796;
 wire net1797;
 wire net1798;
 wire net1799;
 wire net1800;
 wire net1801;
 wire net1802;
 wire net1803;
 wire net1804;
 wire net1805;
 wire net1806;
 wire net1807;
 wire net1808;
 wire net1809;
 wire net1810;
 wire net1811;
 wire net1812;
 wire net1813;
 wire net1814;
 wire net1815;
 wire net1816;
 wire net1817;
 wire net1818;
 wire net1819;
 wire net1820;
 wire net1821;
 wire net1822;
 wire net1823;
 wire net1824;
 wire net1825;
 wire net1826;
 wire net1827;
 wire net1828;
 wire net1829;
 wire net1830;
 wire net1831;
 wire net1832;
 wire net1833;
 wire net1834;
 wire net1835;
 wire net1836;
 wire net1837;
 wire net1838;
 wire net1839;
 wire net1840;
 wire net1841;
 wire net1842;
 wire net1843;
 wire net1844;
 wire net1845;
 wire net1846;
 wire net1847;
 wire net1848;
 wire net1849;
 wire net1850;
 wire net1851;
 wire net1852;
 wire net1853;
 wire net1854;
 wire net1855;
 wire net1856;
 wire net1857;
 wire net1858;
 wire net1859;
 wire net1860;
 wire net1861;
 wire net1862;
 wire net1863;
 wire net1864;
 wire net1865;
 wire net1866;
 wire net1867;
 wire net1868;
 wire net1869;
 wire net1870;
 wire net1871;
 wire net1872;
 wire net1873;
 wire net1874;
 wire net1875;
 wire net1876;
 wire net1877;
 wire net1878;
 wire net1879;
 wire net1880;
 wire net1881;
 wire net1882;
 wire net1883;
 wire net1884;
 wire net1885;
 wire net1886;
 wire net1887;
 wire net1888;
 wire net1889;
 wire net1890;
 wire net1891;
 wire net1892;
 wire net1893;
 wire net1894;
 wire net1895;
 wire net1896;
 wire net1897;
 wire net1898;
 wire net1899;
 wire net1900;
 wire net1901;
 wire net1902;
 wire net1903;
 wire net1904;
 wire net1905;
 wire net1906;
 wire net1907;
 wire net1908;
 wire net1909;
 wire net1910;
 wire net1911;
 wire net1912;
 wire net1913;
 wire net1914;
 wire net1915;
 wire net1916;
 wire net1917;
 wire net1918;
 wire net1919;
 wire net1920;
 wire net1921;
 wire net1922;
 wire net1923;
 wire net1924;
 wire net1925;
 wire net1926;
 wire net1927;
 wire net1928;
 wire net1929;
 wire net1930;
 wire net1931;
 wire net1932;
 wire net1933;
 wire net1934;
 wire net1935;
 wire net1936;
 wire net1937;
 wire net1938;
 wire net1939;
 wire net1940;
 wire net1941;
 wire net1942;
 wire net1943;
 wire net1944;
 wire net1945;
 wire net1946;
 wire net1947;
 wire net1948;
 wire net1949;
 wire net1950;
 wire net1951;
 wire net1952;
 wire net1953;
 wire net1954;
 wire net1955;
 wire net1956;
 wire net1957;
 wire net1958;
 wire net1959;
 wire net1960;
 wire net1961;
 wire net1962;
 wire net1963;
 wire net1964;
 wire net1965;
 wire net1966;
 wire net1967;
 wire net1968;
 wire net1969;
 wire net1970;
 wire net1971;
 wire net1972;
 wire net1973;
 wire net1974;
 wire net1975;
 wire net1976;
 wire net1977;
 wire net1978;
 wire net1979;
 wire net1980;
 wire net1981;
 wire net1982;
 wire net1983;
 wire net1984;
 wire net1985;
 wire net1986;
 wire net1987;
 wire net1988;
 wire net1989;
 wire net1990;
 wire net1991;
 wire net1992;
 wire net1993;
 wire net1994;
 wire net1995;
 wire net1996;
 wire net1997;
 wire net1998;
 wire net1999;
 wire net2000;
 wire net2001;
 wire net2002;
 wire net2003;
 wire net2004;
 wire net2005;
 wire net2006;
 wire net2007;
 wire net2008;
 wire net2009;
 wire net2010;
 wire net2011;
 wire net2012;
 wire net2013;
 wire net2014;
 wire net2015;
 wire net2016;
 wire net2017;
 wire net2018;
 wire net2019;
 wire net2020;
 wire net2021;
 wire net2022;
 wire net2023;
 wire net2024;
 wire net2025;
 wire net2026;
 wire net2027;
 wire net2028;
 wire net2029;
 wire net2030;
 wire net2031;
 wire net2032;
 wire net2033;
 wire net2034;
 wire net2035;
 wire net2036;
 wire net2037;
 wire net2038;
 wire net2039;
 wire net2040;
 wire net2041;
 wire net2042;
 wire net2043;
 wire net2044;
 wire net2045;
 wire net2046;
 wire net2047;
 wire net2048;
 wire net2049;
 wire net2050;
 wire net2051;
 wire net2052;
 wire net2053;
 wire net2054;
 wire net2055;
 wire net2056;
 wire net2057;
 wire net2058;
 wire net2059;
 wire net2060;
 wire net2061;
 wire net2062;
 wire net2063;
 wire net2064;
 wire net2065;
 wire net2066;
 wire net2067;
 wire net2068;
 wire net2069;
 wire net2070;
 wire net2071;
 wire net2072;
 wire net2073;
 wire net2074;
 wire net2075;
 wire net2076;
 wire net2077;
 wire net2078;
 wire net2079;
 wire net2080;
 wire net2081;
 wire net2082;
 wire net2083;
 wire net2084;
 wire net2085;
 wire net2086;
 wire net2087;
 wire net2088;
 wire net2089;
 wire net2090;
 wire net2091;
 wire net2092;
 wire net2093;
 wire net2094;
 wire net2095;
 wire net2096;
 wire net2097;
 wire net2098;
 wire net2099;
 wire net2100;
 wire net2101;
 wire net2102;
 wire net2103;
 wire net2104;
 wire net2105;
 wire net2106;
 wire net2107;
 wire net2108;
 wire net2109;
 wire net2110;
 wire net2111;
 wire net2112;
 wire net2113;
 wire net2114;
 wire net2115;
 wire net2116;
 wire net2117;
 wire net2118;
 wire net2119;
 wire net2120;
 wire net2121;
 wire net2122;
 wire net2123;
 wire net2124;
 wire net2125;
 wire net2126;
 wire net2127;
 wire net2128;
 wire net2129;
 wire net2130;
 wire net2131;
 wire net2132;
 wire net2133;
 wire net2134;
 wire net2135;
 wire net2136;
 wire net2137;
 wire net2138;
 wire net2139;
 wire net2140;
 wire net2141;
 wire net2142;
 wire net2143;
 wire net2144;
 wire net2145;
 wire net2146;
 wire net2147;
 wire net2148;
 wire net2149;
 wire net2150;
 wire net2151;
 wire net2152;
 wire net2153;
 wire net2154;
 wire net2155;
 wire net2156;
 wire net2157;
 wire net2158;
 wire net2159;
 wire net2160;
 wire net2161;
 wire net2162;
 wire net2163;
 wire net2164;
 wire net2165;
 wire net2166;
 wire net2167;
 wire net2168;
 wire net2169;
 wire net2170;
 wire net2171;
 wire net2172;
 wire net2173;
 wire net2174;
 wire net2175;
 wire net2176;
 wire net2177;
 wire net2178;
 wire net2179;
 wire net2180;
 wire net2181;
 wire net2182;
 wire net2183;
 wire net2184;
 wire net2185;
 wire net2186;
 wire net2187;
 wire net2188;
 wire net2189;
 wire net2190;
 wire net2191;
 wire net2192;
 wire net2193;
 wire net2194;
 wire net2195;
 wire net2196;
 wire net2197;
 wire net2198;
 wire net2199;
 wire net2200;
 wire net2201;
 wire net2202;
 wire net2203;
 wire net2204;
 wire net2205;
 wire net2206;
 wire net2207;
 wire net2208;
 wire net2209;
 wire net2210;
 wire net2211;
 wire net2212;
 wire net2213;
 wire net2214;
 wire net2215;
 wire net2216;
 wire net2217;
 wire net2218;
 wire net2219;
 wire net2220;
 wire net2221;
 wire net2222;
 wire net2223;
 wire net2224;
 wire net2225;
 wire net2226;
 wire net2227;
 wire net2228;
 wire net2229;
 wire net2230;
 wire net2231;
 wire net2232;
 wire net2233;
 wire net2234;
 wire net2235;
 wire net2236;
 wire net2237;
 wire net2238;
 wire net2239;
 wire net2240;
 wire net2241;
 wire net2242;
 wire net2243;
 wire net2244;
 wire net2245;
 wire net2246;
 wire net2247;
 wire net2248;
 wire net2249;
 wire net2250;
 wire net2251;
 wire net2252;
 wire net2253;
 wire net2254;
 wire net2255;
 wire net2256;
 wire net2257;
 wire net2258;
 wire net2259;
 wire net2260;
 wire net2261;
 wire net2262;
 wire net2263;
 wire net2264;
 wire net2265;
 wire net2266;
 wire net2267;
 wire net2268;
 wire net2269;
 wire net2270;
 wire net2271;
 wire net2272;
 wire net2273;
 wire net2274;
 wire net2275;
 wire net2276;
 wire net2277;
 wire net2278;
 wire net2279;
 wire net2280;
 wire net2281;
 wire net2282;
 wire net2283;
 wire net2284;
 wire net2285;
 wire net2286;
 wire net2287;
 wire net2288;
 wire net2289;
 wire net2290;
 wire net2291;
 wire net2292;
 wire net2293;
 wire net2294;
 wire net2295;
 wire net2296;
 wire net2297;
 wire net2298;
 wire net2299;
 wire net2300;
 wire net2301;
 wire net2302;
 wire net2303;
 wire net2304;
 wire net2305;
 wire net2306;
 wire net2307;
 wire net2308;
 wire net2309;
 wire net2310;
 wire net2311;
 wire net2312;
 wire net2313;
 wire net2314;
 wire net2315;
 wire net2316;
 wire net2317;
 wire net2318;
 wire net2319;
 wire net2320;
 wire net2321;
 wire net2322;
 wire net2323;
 wire net2324;
 wire net2325;
 wire net2326;
 wire net2327;
 wire net2328;
 wire net2329;
 wire net2330;
 wire net2331;
 wire net2332;
 wire net2333;
 wire net2334;
 wire net2335;
 wire net2336;
 wire net2337;
 wire net2338;
 wire net2339;
 wire net2340;
 wire net2341;
 wire net2342;
 wire net2343;
 wire net2344;
 wire net2345;
 wire net2346;
 wire net2347;
 wire net2348;
 wire net2349;
 wire net2350;
 wire net2351;
 wire net2352;
 wire net2353;
 wire net2354;
 wire net2355;
 wire net2356;
 wire net2357;
 wire net2358;
 wire net2359;
 wire net2360;
 wire net2361;
 wire net2362;
 wire net2363;
 wire net2364;
 wire net2365;
 wire net2366;
 wire net2367;
 wire net2368;
 wire net2369;
 wire net2370;
 wire net2371;
 wire net2372;
 wire net2373;
 wire net2374;
 wire net2375;
 wire net2376;
 wire net2377;
 wire net2378;
 wire net2379;
 wire net2380;
 wire net2381;
 wire net2382;
 wire net2383;
 wire net2384;
 wire net2385;
 wire net2386;
 wire net2387;
 wire net2388;
 wire net2389;
 wire net2390;
 wire net2391;
 wire net2392;
 wire net2393;
 wire net2394;
 wire net2395;
 wire net2396;
 wire net2397;
 wire net2398;
 wire net2399;
 wire net2400;
 wire net2401;
 wire net2402;
 wire net2403;
 wire net2404;
 wire net2405;
 wire net2406;
 wire net2407;
 wire net2408;
 wire net2409;
 wire net2410;
 wire net2411;
 wire net2412;
 wire net2413;
 wire net2414;
 wire net2415;
 wire net2416;
 wire net2417;
 wire net2418;
 wire net2419;
 wire net2420;
 wire net2421;
 wire net2422;
 wire net2423;
 wire net2424;
 wire net2425;
 wire net2426;
 wire net2427;
 wire net2428;
 wire net2429;
 wire net2430;
 wire net2431;
 wire net2432;
 wire net2433;
 wire net2434;
 wire net2435;
 wire net2436;
 wire net2437;
 wire net2438;
 wire net2439;
 wire net2440;
 wire net2441;
 wire net2442;
 wire net2443;
 wire net2444;
 wire net2445;
 wire net2446;
 wire net2447;
 wire net2448;
 wire net2449;
 wire net2450;
 wire net2451;
 wire net2452;
 wire net2453;
 wire net2454;
 wire net2455;
 wire net2456;
 wire net2457;
 wire net2458;
 wire net2459;
 wire net2460;
 wire net2461;
 wire net2462;
 wire net2463;
 wire net2464;
 wire net2465;
 wire net2466;
 wire net2467;
 wire net2468;
 wire net2469;
 wire net2470;
 wire net2471;
 wire net2472;
 wire net2473;
 wire net2474;
 wire net2475;
 wire net2476;
 wire net2477;
 wire net2478;
 wire clknet_leaf_1_clk_p2c;
 wire clknet_leaf_2_clk_p2c;
 wire clknet_leaf_3_clk_p2c;
 wire clknet_leaf_4_clk_p2c;
 wire clknet_leaf_5_clk_p2c;
 wire clknet_leaf_6_clk_p2c;
 wire clknet_leaf_7_clk_p2c;
 wire clknet_leaf_8_clk_p2c;
 wire clknet_leaf_9_clk_p2c;
 wire clknet_leaf_10_clk_p2c;
 wire clknet_leaf_11_clk_p2c;
 wire clknet_leaf_12_clk_p2c;
 wire clknet_leaf_13_clk_p2c;
 wire clknet_leaf_14_clk_p2c;
 wire clknet_leaf_15_clk_p2c;
 wire clknet_leaf_16_clk_p2c;
 wire clknet_leaf_17_clk_p2c;
 wire clknet_leaf_18_clk_p2c;
 wire clknet_leaf_19_clk_p2c;
 wire clknet_leaf_20_clk_p2c;
 wire clknet_leaf_21_clk_p2c;
 wire clknet_leaf_22_clk_p2c;
 wire clknet_leaf_23_clk_p2c;
 wire clknet_leaf_24_clk_p2c;
 wire clknet_leaf_25_clk_p2c;
 wire clknet_leaf_26_clk_p2c;
 wire clknet_leaf_27_clk_p2c;
 wire clknet_leaf_28_clk_p2c;
 wire clknet_leaf_29_clk_p2c;
 wire clknet_leaf_30_clk_p2c;
 wire clknet_leaf_31_clk_p2c;
 wire clknet_leaf_32_clk_p2c;
 wire clknet_leaf_33_clk_p2c;
 wire clknet_leaf_34_clk_p2c;
 wire clknet_leaf_35_clk_p2c;
 wire clknet_leaf_36_clk_p2c;
 wire clknet_leaf_37_clk_p2c;
 wire clknet_leaf_38_clk_p2c;
 wire clknet_leaf_39_clk_p2c;
 wire clknet_leaf_40_clk_p2c;
 wire clknet_leaf_41_clk_p2c;
 wire clknet_leaf_42_clk_p2c;
 wire clknet_leaf_43_clk_p2c;
 wire clknet_leaf_44_clk_p2c;
 wire clknet_leaf_45_clk_p2c;
 wire clknet_leaf_46_clk_p2c;
 wire clknet_leaf_47_clk_p2c;
 wire clknet_leaf_48_clk_p2c;
 wire clknet_leaf_49_clk_p2c;
 wire clknet_leaf_50_clk_p2c;
 wire clknet_leaf_51_clk_p2c;
 wire clknet_leaf_52_clk_p2c;
 wire clknet_leaf_53_clk_p2c;
 wire clknet_leaf_54_clk_p2c;
 wire clknet_leaf_55_clk_p2c;
 wire clknet_leaf_56_clk_p2c;
 wire clknet_leaf_57_clk_p2c;
 wire clknet_leaf_58_clk_p2c;
 wire clknet_leaf_59_clk_p2c;
 wire clknet_leaf_60_clk_p2c;
 wire clknet_leaf_61_clk_p2c;
 wire clknet_leaf_62_clk_p2c;
 wire clknet_leaf_63_clk_p2c;
 wire clknet_leaf_64_clk_p2c;
 wire clknet_leaf_65_clk_p2c;
 wire clknet_leaf_66_clk_p2c;
 wire clknet_leaf_67_clk_p2c;
 wire clknet_leaf_68_clk_p2c;
 wire clknet_leaf_69_clk_p2c;
 wire clknet_leaf_70_clk_p2c;
 wire clknet_leaf_71_clk_p2c;
 wire clknet_leaf_72_clk_p2c;
 wire clknet_leaf_73_clk_p2c;
 wire clknet_leaf_74_clk_p2c;
 wire clknet_leaf_75_clk_p2c;
 wire clknet_leaf_76_clk_p2c;
 wire clknet_leaf_77_clk_p2c;
 wire clknet_leaf_78_clk_p2c;
 wire clknet_leaf_79_clk_p2c;
 wire clknet_leaf_80_clk_p2c;
 wire clknet_leaf_81_clk_p2c;
 wire clknet_leaf_82_clk_p2c;
 wire clknet_leaf_83_clk_p2c;
 wire clknet_leaf_84_clk_p2c;
 wire clknet_leaf_85_clk_p2c;
 wire clknet_leaf_86_clk_p2c;
 wire clknet_leaf_87_clk_p2c;
 wire clknet_leaf_88_clk_p2c;
 wire clknet_leaf_89_clk_p2c;
 wire clknet_leaf_90_clk_p2c;
 wire clknet_leaf_91_clk_p2c;
 wire clknet_leaf_92_clk_p2c;
 wire clknet_leaf_93_clk_p2c;
 wire clknet_leaf_94_clk_p2c;
 wire clknet_leaf_95_clk_p2c;
 wire clknet_leaf_96_clk_p2c;
 wire clknet_leaf_97_clk_p2c;
 wire clknet_leaf_98_clk_p2c;
 wire clknet_leaf_99_clk_p2c;
 wire clknet_leaf_100_clk_p2c;
 wire clknet_leaf_101_clk_p2c;
 wire clknet_leaf_102_clk_p2c;
 wire clknet_leaf_103_clk_p2c;
 wire clknet_leaf_104_clk_p2c;
 wire clknet_leaf_105_clk_p2c;
 wire clknet_leaf_106_clk_p2c;
 wire clknet_leaf_107_clk_p2c;
 wire clknet_leaf_108_clk_p2c;
 wire clknet_leaf_109_clk_p2c;
 wire clknet_leaf_110_clk_p2c;
 wire clknet_leaf_111_clk_p2c;
 wire clknet_leaf_112_clk_p2c;
 wire clknet_leaf_113_clk_p2c;
 wire clknet_leaf_114_clk_p2c;
 wire clknet_leaf_115_clk_p2c;
 wire clknet_leaf_116_clk_p2c;
 wire clknet_leaf_117_clk_p2c;
 wire clknet_leaf_118_clk_p2c;
 wire clknet_leaf_119_clk_p2c;
 wire clknet_leaf_120_clk_p2c;
 wire clknet_leaf_121_clk_p2c;
 wire clknet_leaf_122_clk_p2c;
 wire clknet_leaf_123_clk_p2c;
 wire clknet_leaf_124_clk_p2c;
 wire clknet_leaf_125_clk_p2c;
 wire clknet_leaf_126_clk_p2c;
 wire clknet_leaf_127_clk_p2c;
 wire clknet_leaf_128_clk_p2c;
 wire clknet_leaf_129_clk_p2c;
 wire clknet_leaf_130_clk_p2c;
 wire clknet_leaf_131_clk_p2c;
 wire clknet_leaf_132_clk_p2c;
 wire clknet_leaf_133_clk_p2c;
 wire clknet_leaf_134_clk_p2c;
 wire clknet_leaf_135_clk_p2c;
 wire clknet_leaf_136_clk_p2c;
 wire clknet_leaf_137_clk_p2c;
 wire clknet_leaf_138_clk_p2c;
 wire clknet_leaf_139_clk_p2c;
 wire clknet_leaf_140_clk_p2c;
 wire clknet_leaf_141_clk_p2c;
 wire clknet_leaf_142_clk_p2c;
 wire clknet_leaf_143_clk_p2c;
 wire clknet_leaf_144_clk_p2c;
 wire clknet_leaf_145_clk_p2c;
 wire clknet_leaf_146_clk_p2c;
 wire clknet_leaf_147_clk_p2c;
 wire clknet_leaf_148_clk_p2c;
 wire clknet_leaf_149_clk_p2c;
 wire clknet_leaf_150_clk_p2c;
 wire clknet_leaf_151_clk_p2c;
 wire clknet_leaf_152_clk_p2c;
 wire clknet_leaf_153_clk_p2c;
 wire clknet_leaf_154_clk_p2c;
 wire clknet_leaf_155_clk_p2c;
 wire clknet_leaf_156_clk_p2c;
 wire clknet_leaf_157_clk_p2c;
 wire clknet_leaf_158_clk_p2c;
 wire clknet_leaf_159_clk_p2c;
 wire clknet_leaf_160_clk_p2c;
 wire clknet_leaf_161_clk_p2c;
 wire clknet_leaf_162_clk_p2c;
 wire clknet_leaf_163_clk_p2c;
 wire clknet_leaf_164_clk_p2c;
 wire clknet_leaf_165_clk_p2c;
 wire clknet_leaf_166_clk_p2c;
 wire clknet_leaf_167_clk_p2c;
 wire clknet_leaf_168_clk_p2c;
 wire clknet_leaf_169_clk_p2c;
 wire clknet_leaf_170_clk_p2c;
 wire clknet_leaf_171_clk_p2c;
 wire clknet_leaf_172_clk_p2c;
 wire clknet_leaf_173_clk_p2c;
 wire clknet_leaf_174_clk_p2c;
 wire clknet_leaf_175_clk_p2c;
 wire clknet_leaf_176_clk_p2c;
 wire clknet_leaf_177_clk_p2c;
 wire clknet_leaf_178_clk_p2c;
 wire clknet_leaf_179_clk_p2c;
 wire clknet_leaf_180_clk_p2c;
 wire clknet_leaf_181_clk_p2c;
 wire clknet_leaf_182_clk_p2c;
 wire clknet_leaf_183_clk_p2c;
 wire clknet_leaf_184_clk_p2c;
 wire clknet_leaf_185_clk_p2c;
 wire clknet_leaf_186_clk_p2c;
 wire clknet_leaf_187_clk_p2c;
 wire clknet_leaf_188_clk_p2c;
 wire clknet_leaf_189_clk_p2c;
 wire clknet_leaf_190_clk_p2c;
 wire clknet_leaf_191_clk_p2c;
 wire clknet_leaf_192_clk_p2c;
 wire clknet_leaf_193_clk_p2c;
 wire clknet_leaf_194_clk_p2c;
 wire clknet_leaf_195_clk_p2c;
 wire clknet_leaf_196_clk_p2c;
 wire clknet_leaf_197_clk_p2c;
 wire clknet_leaf_198_clk_p2c;
 wire clknet_leaf_199_clk_p2c;
 wire clknet_leaf_200_clk_p2c;
 wire clknet_leaf_201_clk_p2c;
 wire clknet_leaf_202_clk_p2c;
 wire clknet_leaf_203_clk_p2c;
 wire clknet_leaf_204_clk_p2c;
 wire clknet_leaf_205_clk_p2c;
 wire clknet_leaf_206_clk_p2c;
 wire clknet_leaf_207_clk_p2c;
 wire clknet_leaf_208_clk_p2c;
 wire clknet_leaf_209_clk_p2c;
 wire clknet_leaf_210_clk_p2c;
 wire clknet_leaf_211_clk_p2c;
 wire clknet_leaf_212_clk_p2c;
 wire clknet_leaf_213_clk_p2c;
 wire clknet_leaf_214_clk_p2c;
 wire clknet_leaf_215_clk_p2c;
 wire clknet_leaf_216_clk_p2c;
 wire clknet_leaf_217_clk_p2c;
 wire clknet_leaf_218_clk_p2c;
 wire clknet_leaf_219_clk_p2c;
 wire clknet_leaf_220_clk_p2c;
 wire clknet_leaf_221_clk_p2c;
 wire clknet_leaf_222_clk_p2c;
 wire clknet_leaf_223_clk_p2c;
 wire clknet_leaf_224_clk_p2c;
 wire clknet_leaf_225_clk_p2c;
 wire clknet_leaf_226_clk_p2c;
 wire clknet_leaf_227_clk_p2c;
 wire clknet_leaf_228_clk_p2c;
 wire clknet_leaf_229_clk_p2c;
 wire clknet_leaf_230_clk_p2c;
 wire clknet_leaf_231_clk_p2c;
 wire clknet_leaf_232_clk_p2c;
 wire clknet_leaf_233_clk_p2c;
 wire clknet_leaf_234_clk_p2c;
 wire clknet_leaf_235_clk_p2c;
 wire clknet_leaf_236_clk_p2c;
 wire clknet_leaf_237_clk_p2c;
 wire clknet_leaf_238_clk_p2c;
 wire clknet_leaf_239_clk_p2c;
 wire clknet_leaf_240_clk_p2c;
 wire clknet_leaf_241_clk_p2c;
 wire clknet_leaf_242_clk_p2c;
 wire clknet_leaf_243_clk_p2c;
 wire clknet_leaf_244_clk_p2c;
 wire clknet_leaf_245_clk_p2c;
 wire clknet_leaf_246_clk_p2c;
 wire clknet_leaf_247_clk_p2c;
 wire clknet_leaf_248_clk_p2c;
 wire clknet_leaf_249_clk_p2c;
 wire clknet_leaf_250_clk_p2c;
 wire clknet_leaf_251_clk_p2c;
 wire clknet_leaf_252_clk_p2c;
 wire clknet_leaf_253_clk_p2c;
 wire clknet_leaf_254_clk_p2c;
 wire clknet_leaf_255_clk_p2c;
 wire clknet_leaf_256_clk_p2c;
 wire clknet_leaf_257_clk_p2c;
 wire clknet_leaf_258_clk_p2c;
 wire clknet_leaf_259_clk_p2c;
 wire clknet_leaf_260_clk_p2c;
 wire clknet_leaf_261_clk_p2c;
 wire clknet_leaf_262_clk_p2c;
 wire clknet_leaf_263_clk_p2c;
 wire clknet_leaf_264_clk_p2c;
 wire clknet_leaf_265_clk_p2c;
 wire clknet_leaf_266_clk_p2c;
 wire clknet_leaf_267_clk_p2c;
 wire clknet_leaf_268_clk_p2c;
 wire clknet_leaf_269_clk_p2c;
 wire clknet_leaf_270_clk_p2c;
 wire clknet_leaf_271_clk_p2c;
 wire clknet_leaf_272_clk_p2c;
 wire clknet_leaf_273_clk_p2c;
 wire clknet_leaf_274_clk_p2c;
 wire clknet_leaf_275_clk_p2c;
 wire clknet_leaf_276_clk_p2c;
 wire clknet_leaf_277_clk_p2c;
 wire clknet_leaf_278_clk_p2c;
 wire clknet_leaf_279_clk_p2c;
 wire clknet_leaf_280_clk_p2c;
 wire clknet_leaf_281_clk_p2c;
 wire clknet_leaf_282_clk_p2c;
 wire clknet_leaf_283_clk_p2c;
 wire clknet_leaf_284_clk_p2c;
 wire clknet_leaf_285_clk_p2c;
 wire clknet_leaf_286_clk_p2c;
 wire clknet_leaf_287_clk_p2c;
 wire clknet_leaf_288_clk_p2c;
 wire clknet_leaf_289_clk_p2c;
 wire clknet_leaf_290_clk_p2c;
 wire clknet_leaf_291_clk_p2c;
 wire clknet_leaf_292_clk_p2c;
 wire clknet_leaf_293_clk_p2c;
 wire clknet_0_clk_p2c;
 wire clknet_4_0_0_clk_p2c;
 wire clknet_4_1_0_clk_p2c;
 wire clknet_4_2_0_clk_p2c;
 wire clknet_4_3_0_clk_p2c;
 wire clknet_4_4_0_clk_p2c;
 wire clknet_4_5_0_clk_p2c;
 wire clknet_4_6_0_clk_p2c;
 wire clknet_4_7_0_clk_p2c;
 wire clknet_4_8_0_clk_p2c;
 wire clknet_4_9_0_clk_p2c;
 wire clknet_4_10_0_clk_p2c;
 wire clknet_4_11_0_clk_p2c;
 wire clknet_4_12_0_clk_p2c;
 wire clknet_4_13_0_clk_p2c;
 wire clknet_4_14_0_clk_p2c;
 wire clknet_4_15_0_clk_p2c;
 wire clknet_5_0__leaf_clk_p2c;
 wire clknet_5_1__leaf_clk_p2c;
 wire clknet_5_2__leaf_clk_p2c;
 wire clknet_5_3__leaf_clk_p2c;
 wire clknet_5_4__leaf_clk_p2c;
 wire clknet_5_5__leaf_clk_p2c;
 wire clknet_5_6__leaf_clk_p2c;
 wire clknet_5_7__leaf_clk_p2c;
 wire clknet_5_8__leaf_clk_p2c;
 wire clknet_5_9__leaf_clk_p2c;
 wire clknet_5_10__leaf_clk_p2c;
 wire clknet_5_11__leaf_clk_p2c;
 wire clknet_5_12__leaf_clk_p2c;
 wire clknet_5_13__leaf_clk_p2c;
 wire clknet_5_14__leaf_clk_p2c;
 wire clknet_5_15__leaf_clk_p2c;
 wire clknet_5_16__leaf_clk_p2c;
 wire clknet_5_17__leaf_clk_p2c;
 wire clknet_5_18__leaf_clk_p2c;
 wire clknet_5_19__leaf_clk_p2c;
 wire clknet_5_20__leaf_clk_p2c;
 wire clknet_5_21__leaf_clk_p2c;
 wire clknet_5_22__leaf_clk_p2c;
 wire clknet_5_23__leaf_clk_p2c;
 wire clknet_5_24__leaf_clk_p2c;
 wire clknet_5_25__leaf_clk_p2c;
 wire clknet_5_26__leaf_clk_p2c;
 wire clknet_5_27__leaf_clk_p2c;
 wire clknet_5_28__leaf_clk_p2c;
 wire clknet_5_29__leaf_clk_p2c;
 wire clknet_5_30__leaf_clk_p2c;
 wire clknet_5_31__leaf_clk_p2c;

 sg13g2_buf_4 fanout608 (.X(net608),
    .A(net611));
 sg13g2_buf_1 fanout607 (.A(net618),
    .X(net607));
 sg13g2_buf_2 fanout606 (.A(net607),
    .X(net606));
 sg13g2_buf_2 fanout605 (.A(net606),
    .X(net605));
 sg13g2_nor2b_1 _06973_ (.A(net164),
    .B_N(net112),
    .Y(_01707_));
 sg13g2_buf_4 fanout604 (.X(net604),
    .A(net606));
 sg13g2_inv_1 _06975_ (.Y(_01709_),
    .A(net161));
 sg13g2_o21ai_1 _06976_ (.B1(_01709_),
    .Y(_01710_),
    .A1(net110),
    .A2(_01707_));
 sg13g2_buf_1 fanout603 (.A(net607),
    .X(net603));
 sg13g2_inv_2 _06978_ (.Y(_01712_),
    .A(net105));
 sg13g2_buf_4 fanout602 (.X(net602),
    .A(net603));
 sg13g2_buf_4 fanout601 (.X(net601),
    .A(net603));
 sg13g2_nand2b_1 _06981_ (.Y(_01715_),
    .B(net107),
    .A_N(net159));
 sg13g2_nand3b_1 _06982_ (.B(\median_processor.input_storage[49] ),
    .C(net112),
    .Y(_01716_),
    .A_N(net163));
 sg13g2_and3_1 _06983_ (.X(_01717_),
    .A(_01712_),
    .B(_01715_),
    .C(_01716_));
 sg13g2_buf_2 fanout600 (.A(net603),
    .X(net600));
 sg13g2_inv_2 _06985_ (.Y(_01719_),
    .A(net158));
 sg13g2_buf_4 fanout599 (.X(net599),
    .A(net600));
 sg13g2_nand2b_1 _06987_ (.Y(_01721_),
    .B(\median_processor.input_storage[26] ),
    .A_N(\median_processor.input_storage[50] ));
 sg13g2_a21oi_1 _06988_ (.A1(_01719_),
    .A2(net106),
    .Y(_01722_),
    .B1(_01721_));
 sg13g2_a21oi_1 _06989_ (.A1(_01710_),
    .A2(_01717_),
    .Y(_01723_),
    .B1(_01722_));
 sg13g2_buf_4 fanout598 (.X(net598),
    .A(net600));
 sg13g2_and3_1 _06991_ (.X(_01725_),
    .A(net158),
    .B(_01715_),
    .C(_01716_));
 sg13g2_a22oi_1 _06992_ (.Y(_01726_),
    .B1(_01710_),
    .B2(_01725_),
    .A2(_01712_),
    .A1(net157));
 sg13g2_buf_1 fanout597 (.A(net618),
    .X(net597));
 sg13g2_buf_2 fanout596 (.A(net597),
    .X(net596));
 sg13g2_buf_4 fanout595 (.X(net595),
    .A(net596));
 sg13g2_inv_2 _06996_ (.Y(_01730_),
    .A(net102));
 sg13g2_buf_1 fanout594 (.A(net597),
    .X(net594));
 sg13g2_buf_4 fanout593 (.X(net593),
    .A(net597));
 sg13g2_inv_2 _06999_ (.Y(_01733_),
    .A(net103));
 sg13g2_buf_2 fanout592 (.A(net597),
    .X(net592));
 sg13g2_buf_4 fanout591 (.X(net591),
    .A(net592));
 sg13g2_a22oi_1 _07002_ (.Y(_01736_),
    .B1(_01733_),
    .B2(net155),
    .A2(_01730_),
    .A1(net153));
 sg13g2_buf_2 fanout590 (.A(net597),
    .X(net590));
 sg13g2_buf_4 fanout589 (.X(net589),
    .A(net597));
 sg13g2_buf_1 fanout588 (.A(net775),
    .X(net588));
 sg13g2_buf_1 fanout587 (.A(net588),
    .X(net587));
 sg13g2_inv_2 _07007_ (.Y(_01741_),
    .A(net98));
 sg13g2_buf_2 fanout586 (.A(net587),
    .X(net586));
 sg13g2_a21oi_1 _07009_ (.A1(net147),
    .A2(net73),
    .Y(_01743_),
    .B1(net148));
 sg13g2_nand4_1 _07010_ (.B(_01726_),
    .C(_01736_),
    .A(_01723_),
    .Y(_01744_),
    .D(_01743_));
 sg13g2_nand2b_1 _07011_ (.Y(_01745_),
    .B(net104),
    .A_N(net155));
 sg13g2_a21oi_1 _07012_ (.A1(net153),
    .A2(_01745_),
    .Y(_01746_),
    .B1(_01730_));
 sg13g2_nor2_1 _07013_ (.A(net153),
    .B(_01745_),
    .Y(_01747_));
 sg13g2_or2_1 _07014_ (.X(_01748_),
    .B(_01747_),
    .A(_01746_));
 sg13g2_buf_4 fanout585 (.X(net585),
    .A(net586));
 sg13g2_buf_4 fanout584 (.X(net584),
    .A(net586));
 sg13g2_buf_2 fanout583 (.A(net587),
    .X(net583));
 sg13g2_nand2_1 _07018_ (.Y(_01752_),
    .A(net97),
    .B(net100));
 sg13g2_nor2_1 _07019_ (.A(net148),
    .B(_01752_),
    .Y(_01753_));
 sg13g2_a21oi_1 _07020_ (.A1(_01748_),
    .A2(_01743_),
    .Y(_01754_),
    .B1(_01753_));
 sg13g2_inv_2 _07021_ (.Y(_01755_),
    .A(net100));
 sg13g2_a21oi_1 _07022_ (.A1(net147),
    .A2(net73),
    .Y(_01756_),
    .B1(net72));
 sg13g2_nand4_1 _07023_ (.B(_01726_),
    .C(_01736_),
    .A(_01723_),
    .Y(_01757_),
    .D(_01756_));
 sg13g2_o21ai_1 _07024_ (.B1(_01741_),
    .Y(_01758_),
    .A1(net148),
    .A2(_01755_));
 sg13g2_inv_2 _07025_ (.Y(_01759_),
    .A(net146));
 sg13g2_a22oi_1 _07026_ (.Y(_01760_),
    .B1(_01758_),
    .B2(_01759_),
    .A2(_01756_),
    .A1(_01748_));
 sg13g2_and4_1 _07027_ (.A(_01744_),
    .B(_01754_),
    .C(_01757_),
    .D(_01760_),
    .X(_01761_));
 sg13g2_buf_4 fanout582 (.X(net582),
    .A(net583));
 sg13g2_buf_2 fanout581 (.A(net587),
    .X(net581));
 sg13g2_buf_2 fanout580 (.A(net581),
    .X(net580));
 sg13g2_inv_2 _07031_ (.Y(_01765_),
    .A(net113));
 sg13g2_nor2_1 _07032_ (.A(net97),
    .B(net71),
    .Y(_01766_));
 sg13g2_buf_4 fanout579 (.X(net579),
    .A(net580));
 sg13g2_buf_4 fanout578 (.X(net578),
    .A(net581));
 sg13g2_buf_4 fanout577 (.X(net577),
    .A(net581));
 sg13g2_nand2_2 _07036_ (.Y(_01770_),
    .A(net97),
    .B(net71));
 sg13g2_and3_1 _07037_ (.X(_01771_),
    .A(net72),
    .B(net116),
    .C(_01770_));
 sg13g2_buf_2 fanout576 (.A(net588),
    .X(net576));
 sg13g2_inv_2 _07039_ (.Y(_01773_),
    .A(\median_processor.input_storage[41] ));
 sg13g2_buf_4 fanout575 (.X(net575),
    .A(net576));
 sg13g2_buf_4 fanout574 (.X(net574),
    .A(net576));
 sg13g2_nor2b_1 _07042_ (.A(\median_processor.input_storage[40] ),
    .B_N(net111),
    .Y(_01776_));
 sg13g2_o21ai_1 _07043_ (.B1(\median_processor.input_storage[49] ),
    .Y(_01777_),
    .A1(net70),
    .A2(_01776_));
 sg13g2_buf_2 fanout573 (.A(net576),
    .X(net573));
 sg13g2_buf_4 fanout572 (.X(net572),
    .A(net576));
 sg13g2_inv_2 _07046_ (.Y(_01780_),
    .A(net125));
 sg13g2_inv_1 _07047_ (.Y(_01781_),
    .A(net124));
 sg13g2_buf_2 fanout571 (.A(net588),
    .X(net571));
 sg13g2_a221oi_1 _07049_ (.B2(_01776_),
    .C1(net69),
    .B1(net70),
    .A1(net107),
    .Y(_01783_),
    .A2(_01780_));
 sg13g2_buf_4 fanout570 (.X(net570),
    .A(net571));
 sg13g2_buf_2 fanout569 (.A(net571),
    .X(net569));
 sg13g2_nand2b_1 _07052_ (.Y(_01786_),
    .B(net125),
    .A_N(net107));
 sg13g2_a21oi_1 _07053_ (.A1(net105),
    .A2(net69),
    .Y(_01787_),
    .B1(_01786_));
 sg13g2_a21oi_1 _07054_ (.A1(_01777_),
    .A2(_01783_),
    .Y(_01788_),
    .B1(_01787_));
 sg13g2_buf_4 fanout568 (.X(net568),
    .A(net571));
 sg13g2_a221oi_1 _07056_ (.B2(_01776_),
    .C1(net105),
    .B1(net70),
    .A1(net107),
    .Y(_01790_),
    .A2(_01780_));
 sg13g2_a22oi_1 _07057_ (.Y(_01791_),
    .B1(_01777_),
    .B2(_01790_),
    .A2(net123),
    .A1(_01712_));
 sg13g2_buf_1 fanout567 (.A(net588),
    .X(net567));
 sg13g2_buf_2 fanout566 (.A(net567),
    .X(net566));
 sg13g2_nor2_1 _07060_ (.A(net118),
    .B(net121),
    .Y(_01794_));
 sg13g2_nand2_1 _07061_ (.Y(_01795_),
    .A(net104),
    .B(_01794_));
 sg13g2_inv_4 _07062_ (.A(net118),
    .Y(_01796_));
 sg13g2_nor2b_1 _07063_ (.A(net121),
    .B_N(net104),
    .Y(_01797_));
 sg13g2_buf_4 fanout565 (.X(net565),
    .A(net566));
 sg13g2_o21ai_1 _07065_ (.B1(net102),
    .Y(_01799_),
    .A1(net68),
    .A2(_01797_));
 sg13g2_nand4_1 _07066_ (.B(_01795_),
    .C(_01799_),
    .A(net116),
    .Y(_01800_),
    .D(_01770_));
 sg13g2_nand4_1 _07067_ (.B(_01795_),
    .C(_01799_),
    .A(net72),
    .Y(_01801_),
    .D(_01770_));
 sg13g2_a22oi_1 _07068_ (.Y(_01802_),
    .B1(_01800_),
    .B2(_01801_),
    .A2(_01791_),
    .A1(_01788_));
 sg13g2_buf_4 fanout564 (.X(net564),
    .A(net565));
 sg13g2_nand2_1 _07070_ (.Y(_01804_),
    .A(_01733_),
    .B(net121));
 sg13g2_buf_2 fanout563 (.A(net566),
    .X(net563));
 sg13g2_nand2_1 _07072_ (.Y(_01806_),
    .A(_01730_),
    .B(net119));
 sg13g2_nand2_1 _07073_ (.Y(_01807_),
    .A(net116),
    .B(_01770_));
 sg13g2_nand2_1 _07074_ (.Y(_01808_),
    .A(net72),
    .B(_01770_));
 sg13g2_nand2_1 _07075_ (.Y(_01809_),
    .A(_01795_),
    .B(_01799_));
 sg13g2_a221oi_1 _07076_ (.B2(_01808_),
    .C1(_01809_),
    .B1(_01807_),
    .A1(_01804_),
    .Y(_01810_),
    .A2(_01806_));
 sg13g2_or4_2 _07077_ (.A(_01766_),
    .B(_01771_),
    .C(_01802_),
    .D(_01810_),
    .X(_01811_));
 sg13g2_buf_4 fanout562 (.X(net562),
    .A(net563));
 sg13g2_buf_1 fanout561 (.A(net567),
    .X(net561));
 sg13g2_inv_1 _07080_ (.Y(_01814_),
    .A(net85));
 sg13g2_buf_4 fanout560 (.X(net560),
    .A(net561));
 sg13g2_buf_4 fanout559 (.X(net559),
    .A(net561));
 sg13g2_buf_2 fanout558 (.A(net567),
    .X(net558));
 sg13g2_nand2_1 _07084_ (.Y(_01818_),
    .A(net73),
    .B(net83));
 sg13g2_nand2_1 _07085_ (.Y(_01819_),
    .A(net67),
    .B(_01818_));
 sg13g2_nand2_1 _07086_ (.Y(_01820_),
    .A(net99),
    .B(_01818_));
 sg13g2_buf_4 fanout557 (.X(net557),
    .A(net567));
 sg13g2_inv_1 _07088_ (.Y(_01822_),
    .A(net86));
 sg13g2_buf_1 fanout556 (.A(net588),
    .X(net556));
 sg13g2_nand2_1 _07090_ (.Y(_01824_),
    .A(net101),
    .B(net64));
 sg13g2_buf_2 fanout555 (.A(net556),
    .X(net555));
 sg13g2_buf_2 fanout554 (.A(net555),
    .X(net554));
 sg13g2_buf_4 fanout553 (.X(net553),
    .A(net554));
 sg13g2_nand2_1 _07094_ (.Y(_01828_),
    .A(net94),
    .B(net95));
 sg13g2_o21ai_1 _07095_ (.B1(net110),
    .Y(_01829_),
    .A1(net111),
    .A2(_01828_));
 sg13g2_buf_4 fanout552 (.X(net552),
    .A(net555));
 sg13g2_inv_2 _07097_ (.Y(_01831_),
    .A(net92));
 sg13g2_inv_2 _07098_ (.Y(_01832_),
    .A(net94));
 sg13g2_nand2b_1 _07099_ (.Y(_01833_),
    .B(net95),
    .A_N(net111));
 sg13g2_buf_2 fanout551 (.A(net556),
    .X(net551));
 sg13g2_inv_1 _07101_ (.Y(_01835_),
    .A(net90));
 sg13g2_a221oi_1 _07102_ (.B2(_01833_),
    .C1(_01835_),
    .B1(_01832_),
    .A1(net108),
    .Y(_01836_),
    .A2(_01831_));
 sg13g2_buf_4 fanout550 (.X(net550),
    .A(net551));
 sg13g2_nand2b_1 _07104_ (.Y(_01838_),
    .B(net93),
    .A_N(net108));
 sg13g2_a21oi_1 _07105_ (.A1(net106),
    .A2(_01835_),
    .Y(_01839_),
    .B1(_01838_));
 sg13g2_a21oi_1 _07106_ (.A1(_01829_),
    .A2(_01836_),
    .Y(_01840_),
    .B1(_01839_));
 sg13g2_buf_4 fanout549 (.X(net549),
    .A(net551));
 sg13g2_a221oi_1 _07108_ (.B2(_01833_),
    .C1(net106),
    .B1(_01832_),
    .A1(net108),
    .Y(_01842_),
    .A2(_01831_));
 sg13g2_a22oi_1 _07109_ (.Y(_01843_),
    .B1(_01829_),
    .B2(_01842_),
    .A2(net90),
    .A1(_01712_));
 sg13g2_buf_2 fanout548 (.A(net556),
    .X(net548));
 sg13g2_buf_4 fanout547 (.X(net547),
    .A(net556));
 sg13g2_nand2_1 _07112_ (.Y(_01846_),
    .A(_01733_),
    .B(net87));
 sg13g2_nand4_1 _07113_ (.B(_01840_),
    .C(_01843_),
    .A(net64),
    .Y(_01847_),
    .D(_01846_));
 sg13g2_nand4_1 _07114_ (.B(_01840_),
    .C(_01843_),
    .A(net101),
    .Y(_01848_),
    .D(_01846_));
 sg13g2_nor2_1 _07115_ (.A(_01733_),
    .B(net88),
    .Y(_01849_));
 sg13g2_o21ai_1 _07116_ (.B1(_01849_),
    .Y(_01850_),
    .A1(net101),
    .A2(net64));
 sg13g2_and4_1 _07117_ (.A(_01824_),
    .B(_01847_),
    .C(_01848_),
    .D(_01850_),
    .X(_01851_));
 sg13g2_a21oi_2 _07118_ (.B1(_01851_),
    .Y(_01852_),
    .A2(_01820_),
    .A1(_01819_));
 sg13g2_nand3_1 _07119_ (.B(net67),
    .C(_01818_),
    .A(net99),
    .Y(_01853_));
 sg13g2_o21ai_1 _07120_ (.B1(_01853_),
    .Y(_01854_),
    .A1(net73),
    .A2(net82));
 sg13g2_buf_1 fanout546 (.A(net775),
    .X(net546));
 sg13g2_nor4_1 _07122_ (.A(_01761_),
    .B(_01811_),
    .C(_01852_),
    .D(_01854_),
    .Y(_01856_));
 sg13g2_a21o_1 _07123_ (.A2(_01820_),
    .A1(_01819_),
    .B1(_01851_),
    .X(_01857_));
 sg13g2_inv_1 _07124_ (.Y(_01858_),
    .A(_01854_));
 sg13g2_nand4_1 _07125_ (.B(_01754_),
    .C(_01757_),
    .A(_01744_),
    .Y(_01859_),
    .D(_01760_));
 sg13g2_buf_1 fanout545 (.A(net546),
    .X(net545));
 sg13g2_nor4_1 _07127_ (.A(_01766_),
    .B(_01771_),
    .C(_01802_),
    .D(_01810_),
    .Y(_01861_));
 sg13g2_buf_2 fanout544 (.A(net545),
    .X(net544));
 sg13g2_xnor2_1 _07129_ (.Y(_01863_),
    .A(_01859_),
    .B(net31));
 sg13g2_a21oi_1 _07130_ (.A1(_01857_),
    .A2(_01858_),
    .Y(_01864_),
    .B1(_01863_));
 sg13g2_buf_4 fanout543 (.X(net543),
    .A(net544));
 sg13g2_buf_4 fanout542 (.X(net542),
    .A(net544));
 sg13g2_buf_4 fanout541 (.X(net541),
    .A(net544));
 sg13g2_nand2b_1 _07134_ (.Y(_01868_),
    .B(net100),
    .A_N(net167));
 sg13g2_nor2_1 _07135_ (.A(net166),
    .B(net167),
    .Y(_01869_));
 sg13g2_a21oi_1 _07136_ (.A1(net100),
    .A2(_01869_),
    .Y(_01870_),
    .B1(net97));
 sg13g2_a21oi_1 _07137_ (.A1(net166),
    .A2(_01868_),
    .Y(_01871_),
    .B1(_01870_));
 sg13g2_buf_4 fanout540 (.X(net540),
    .A(net544));
 sg13g2_inv_1 _07139_ (.Y(_01873_),
    .A(net170));
 sg13g2_nand2_1 _07140_ (.Y(_01874_),
    .A(net102),
    .B(_01873_));
 sg13g2_buf_2 fanout539 (.A(net545),
    .X(net539));
 sg13g2_buf_4 fanout538 (.X(net538),
    .A(net539));
 sg13g2_inv_2 _07143_ (.Y(_01877_),
    .A(net171));
 sg13g2_nor2_1 _07144_ (.A(net103),
    .B(_01877_),
    .Y(_01878_));
 sg13g2_buf_2 fanout537 (.A(net545),
    .X(net537));
 sg13g2_buf_4 fanout536 (.X(net536),
    .A(net537));
 sg13g2_nor2_1 _07147_ (.A(\median_processor.input_storage[49] ),
    .B(net112),
    .Y(_01881_));
 sg13g2_buf_1 fanout535 (.A(net545),
    .X(net535));
 sg13g2_a21oi_1 _07149_ (.A1(\median_processor.input_storage[16] ),
    .A2(_01881_),
    .Y(_01883_),
    .B1(net177));
 sg13g2_inv_1 _07150_ (.Y(_01884_),
    .A(net112));
 sg13g2_inv_1 _07151_ (.Y(_01885_),
    .A(net110));
 sg13g2_a21oi_1 _07152_ (.A1(_01884_),
    .A2(net178),
    .Y(_01886_),
    .B1(_01885_));
 sg13g2_buf_4 fanout534 (.X(net534),
    .A(net535));
 sg13g2_buf_4 fanout533 (.X(net533),
    .A(net534));
 sg13g2_buf_2 fanout532 (.A(net535),
    .X(net532));
 sg13g2_buf_4 fanout531 (.X(net531),
    .A(net532));
 sg13g2_nor2b_1 _07157_ (.A(net107),
    .B_N(net175),
    .Y(_01891_));
 sg13g2_a21oi_1 _07158_ (.A1(_01712_),
    .A2(net173),
    .Y(_01892_),
    .B1(_01891_));
 sg13g2_o21ai_1 _07159_ (.B1(_01892_),
    .Y(_01893_),
    .A1(_01883_),
    .A2(_01886_));
 sg13g2_a22oi_1 _07160_ (.Y(_01894_),
    .B1(_01877_),
    .B2(net103),
    .A2(_01873_),
    .A1(net102));
 sg13g2_inv_2 _07161_ (.Y(_01895_),
    .A(net173));
 sg13g2_nand2_1 _07162_ (.Y(_01896_),
    .A(net105),
    .B(_01895_));
 sg13g2_nor2b_1 _07163_ (.A(net175),
    .B_N(net107),
    .Y(_01897_));
 sg13g2_o21ai_1 _07164_ (.B1(_01897_),
    .Y(_01898_),
    .A1(net105),
    .A2(_01895_));
 sg13g2_and3_1 _07165_ (.X(_01899_),
    .A(_01894_),
    .B(_01896_),
    .C(_01898_));
 sg13g2_buf_2 fanout530 (.A(net545),
    .X(net530));
 sg13g2_nand2b_1 _07167_ (.Y(_01901_),
    .B(net167),
    .A_N(net99));
 sg13g2_buf_4 fanout529 (.X(net529),
    .A(net530));
 sg13g2_nand2b_1 _07169_ (.Y(_01903_),
    .B(net169),
    .A_N(net102));
 sg13g2_xnor2_1 _07170_ (.Y(_01904_),
    .A(net98),
    .B(net165));
 sg13g2_nand4_1 _07171_ (.B(_01901_),
    .C(_01903_),
    .A(_01868_),
    .Y(_01905_),
    .D(_01904_));
 sg13g2_a221oi_1 _07172_ (.B2(_01899_),
    .C1(_01905_),
    .B1(_01893_),
    .A1(_01874_),
    .Y(_01906_),
    .A2(_01878_));
 sg13g2_xnor2_1 _07173_ (.Y(_01907_),
    .A(net112),
    .B(\median_processor.input_storage[16] ));
 sg13g2_xor2_1 _07174_ (.B(net177),
    .A(net110),
    .X(_01908_));
 sg13g2_nor3_1 _07175_ (.A(_01908_),
    .B(_01891_),
    .C(_01897_),
    .Y(_01909_));
 sg13g2_xor2_1 _07176_ (.B(net174),
    .A(net105),
    .X(_01910_));
 sg13g2_nor3_1 _07177_ (.A(_01905_),
    .B(_01910_),
    .C(_01878_),
    .Y(_01911_));
 sg13g2_nand4_1 _07178_ (.B(_01894_),
    .C(_01909_),
    .A(_01907_),
    .Y(_01912_),
    .D(_01911_));
 sg13g2_o21ai_1 _07179_ (.B1(_01912_),
    .Y(_01913_),
    .A1(_01871_),
    .A2(_01906_));
 sg13g2_buf_4 fanout528 (.X(net528),
    .A(net529));
 sg13g2_buf_4 fanout527 (.X(net527),
    .A(net530));
 sg13g2_buf_1 fanout526 (.A(net546),
    .X(net526));
 sg13g2_buf_2 fanout525 (.A(net526),
    .X(net525));
 sg13g2_inv_2 _07184_ (.Y(_01918_),
    .A(net140));
 sg13g2_buf_4 fanout524 (.X(net524),
    .A(net525));
 sg13g2_nor2b_1 _07186_ (.A(net137),
    .B_N(net103),
    .Y(_01920_));
 sg13g2_buf_2 fanout523 (.A(net526),
    .X(net523));
 sg13g2_inv_1 _07188_ (.Y(_01922_),
    .A(net131));
 sg13g2_a221oi_1 _07189_ (.B2(net63),
    .C1(net105),
    .B1(_01920_),
    .A1(_01918_),
    .Y(_01923_),
    .A2(net107));
 sg13g2_buf_4 fanout522 (.X(net522),
    .A(net526));
 sg13g2_buf_2 fanout521 (.A(net526),
    .X(net521));
 sg13g2_inv_2 _07192_ (.Y(_01926_),
    .A(net139));
 sg13g2_a221oi_1 _07193_ (.B2(net63),
    .C1(net62),
    .B1(_01920_),
    .A1(_01918_),
    .Y(_01927_),
    .A2(net107));
 sg13g2_buf_4 fanout520 (.X(net520),
    .A(net521));
 sg13g2_buf_4 fanout519 (.X(net519),
    .A(net520));
 sg13g2_o21ai_1 _07196_ (.B1(_01885_),
    .Y(_01930_),
    .A1(net144),
    .A2(_01884_));
 sg13g2_inv_1 _07197_ (.Y(_01931_),
    .A(\median_processor.input_storage[50] ));
 sg13g2_buf_2 fanout518 (.A(net521),
    .X(net518));
 sg13g2_buf_4 fanout517 (.X(net517),
    .A(net518));
 sg13g2_a21oi_1 _07200_ (.A1(net140),
    .A2(_01931_),
    .Y(_01934_),
    .B1(net143));
 sg13g2_nand2_1 _07201_ (.Y(_01935_),
    .A(net110),
    .B(net111));
 sg13g2_a21oi_1 _07202_ (.A1(\median_processor.input_storage[34] ),
    .A2(_01931_),
    .Y(_01936_),
    .B1(_01935_));
 sg13g2_inv_1 _07203_ (.Y(_01937_),
    .A(net145));
 sg13g2_a22oi_1 _07204_ (.Y(_01938_),
    .B1(_01936_),
    .B2(_01937_),
    .A2(_01934_),
    .A1(_01930_));
 sg13g2_o21ai_1 _07205_ (.B1(_01938_),
    .Y(_01939_),
    .A1(_01923_),
    .A2(_01927_));
 sg13g2_buf_2 fanout516 (.A(net546),
    .X(net516));
 sg13g2_inv_1 _07207_ (.Y(_01941_),
    .A(net137));
 sg13g2_nor2_1 _07208_ (.A(_01941_),
    .B(net104),
    .Y(_01942_));
 sg13g2_nor2_1 _07209_ (.A(net63),
    .B(net97),
    .Y(_01943_));
 sg13g2_buf_2 fanout515 (.A(net516),
    .X(net515));
 sg13g2_inv_4 _07211_ (.A(net132),
    .Y(_01945_));
 sg13g2_buf_4 fanout514 (.X(net514),
    .A(net516));
 sg13g2_buf_4 fanout513 (.X(net513),
    .A(net516));
 sg13g2_nand2_1 _07214_ (.Y(_01948_),
    .A(net135),
    .B(_01730_));
 sg13g2_o21ai_1 _07215_ (.B1(_01948_),
    .Y(_01949_),
    .A1(net61),
    .A2(net99));
 sg13g2_and2_1 _07216_ (.A(net63),
    .B(_01920_),
    .X(_01950_));
 sg13g2_nor3_1 _07217_ (.A(net62),
    .B(net105),
    .C(_01950_),
    .Y(_01951_));
 sg13g2_nor4_1 _07218_ (.A(_01942_),
    .B(_01943_),
    .C(_01949_),
    .D(_01951_),
    .Y(_01952_));
 sg13g2_and2_1 _07219_ (.A(net98),
    .B(net102),
    .X(_01953_));
 sg13g2_nor2b_1 _07220_ (.A(net135),
    .B_N(net98),
    .Y(_01954_));
 sg13g2_o21ai_1 _07221_ (.B1(_01920_),
    .Y(_01955_),
    .A1(_01953_),
    .A2(_01954_));
 sg13g2_nor2_1 _07222_ (.A(net131),
    .B(net135),
    .Y(_01956_));
 sg13g2_o21ai_1 _07223_ (.B1(net102),
    .Y(_01957_),
    .A1(_01956_),
    .A2(_01954_));
 sg13g2_nand3_1 _07224_ (.B(_01955_),
    .C(_01957_),
    .A(_01752_),
    .Y(_01958_));
 sg13g2_buf_1 fanout512 (.A(net546),
    .X(net512));
 sg13g2_o21ai_1 _07226_ (.B1(_01741_),
    .Y(_01960_),
    .A1(net133),
    .A2(net72));
 sg13g2_a21oi_1 _07227_ (.A1(_01955_),
    .A2(_01957_),
    .Y(_01961_),
    .B1(net72));
 sg13g2_a21o_1 _07228_ (.A2(_01960_),
    .A1(net63),
    .B1(_01961_),
    .X(_01962_));
 sg13g2_a221oi_1 _07229_ (.B2(net61),
    .C1(_01962_),
    .B1(_01958_),
    .A1(_01939_),
    .Y(_01963_),
    .A2(_01952_));
 sg13g2_buf_2 fanout511 (.A(net512),
    .X(net511));
 sg13g2_buf_4 fanout510 (.X(net510),
    .A(net511));
 sg13g2_nor2_1 _07232_ (.A(net29),
    .B(net28),
    .Y(_01966_));
 sg13g2_and2_1 _07233_ (.A(net29),
    .B(net28),
    .X(_01967_));
 sg13g2_nor2_1 _07234_ (.A(_01966_),
    .B(_01967_),
    .Y(_01968_));
 sg13g2_o21ai_1 _07235_ (.B1(_01968_),
    .Y(_01969_),
    .A1(_01856_),
    .A2(_01864_));
 sg13g2_nor2_1 _07236_ (.A(_01859_),
    .B(net31),
    .Y(_01970_));
 sg13g2_nor2_1 _07237_ (.A(net32),
    .B(_01811_),
    .Y(_01971_));
 sg13g2_a22oi_1 _07238_ (.Y(_01972_),
    .B1(_01967_),
    .B2(_01971_),
    .A2(_01966_),
    .A1(_01970_));
 sg13g2_or3_1 _07239_ (.A(net29),
    .B(net28),
    .C(_01863_),
    .X(_01973_));
 sg13g2_nor2_2 _07240_ (.A(_01852_),
    .B(_01854_),
    .Y(_01974_));
 sg13g2_mux2_1 _07241_ (.A0(_01972_),
    .A1(_01973_),
    .S(_01974_),
    .X(_01975_));
 sg13g2_buf_2 fanout509 (.A(net512),
    .X(net509));
 sg13g2_buf_4 fanout508 (.X(net508),
    .A(net509));
 sg13g2_buf_1 fanout507 (.A(net509),
    .X(net507));
 sg13g2_buf_4 fanout506 (.X(net506),
    .A(net509));
 sg13g2_nand2b_1 _07246_ (.Y(_01980_),
    .B(net108),
    .A_N(net195));
 sg13g2_and3_1 _07247_ (.X(_01981_),
    .A(net76),
    .B(_01980_),
    .C(_01881_));
 sg13g2_inv_4 _07248_ (.A(net194),
    .Y(_01982_));
 sg13g2_nand2b_1 _07249_ (.Y(_01983_),
    .B(net76),
    .A_N(net111));
 sg13g2_buf_1 fanout505 (.A(data_in_p2c_2),
    .X(net505));
 sg13g2_inv_4 _07251_ (.A(net74),
    .Y(_01985_));
 sg13g2_a221oi_1 _07252_ (.B2(net110),
    .C1(_01985_),
    .B1(_01983_),
    .A1(net108),
    .Y(_01986_),
    .A2(net60));
 sg13g2_buf_2 fanout504 (.A(net505),
    .X(net504));
 sg13g2_buf_2 fanout503 (.A(data_in_p2c_4),
    .X(net503));
 sg13g2_xnor2_1 _07255_ (.Y(_01989_),
    .A(net103),
    .B(net189));
 sg13g2_buf_1 fanout502 (.A(data_in_p2c_5),
    .X(net502));
 sg13g2_xnor2_1 _07257_ (.Y(_01991_),
    .A(net101),
    .B(net187));
 sg13g2_nand2b_1 _07258_ (.Y(_01992_),
    .B(net194),
    .A_N(net108));
 sg13g2_buf_2 fanout501 (.A(net502),
    .X(net501));
 sg13g2_buf_2 fanout500 (.A(data_in_p2c_6),
    .X(net500));
 sg13g2_nand2b_1 _07261_ (.Y(_01995_),
    .B(net192),
    .A_N(net106));
 sg13g2_nand4_1 _07262_ (.B(_01991_),
    .C(_01992_),
    .A(_01989_),
    .Y(_01996_),
    .D(_01995_));
 sg13g2_or3_1 _07263_ (.A(_01981_),
    .B(_01986_),
    .C(_01996_),
    .X(_01997_));
 sg13g2_inv_1 _07264_ (.Y(_01998_),
    .A(net186));
 sg13g2_inv_1 _07265_ (.Y(_01999_),
    .A(net189));
 sg13g2_buf_1 fanout499 (.A(data_in_p2c_7),
    .X(net499));
 sg13g2_nand2b_1 _07267_ (.Y(_02001_),
    .B(net106),
    .A_N(net192));
 sg13g2_a21oi_1 _07268_ (.A1(_01730_),
    .A2(net186),
    .Y(_02002_),
    .B1(_02001_));
 sg13g2_a221oi_1 _07269_ (.B2(_02001_),
    .C1(_01733_),
    .B1(net190),
    .A1(_01730_),
    .Y(_02003_),
    .A2(net186));
 sg13g2_a221oi_1 _07270_ (.B2(_02002_),
    .C1(_02003_),
    .B1(_01999_),
    .A1(net101),
    .Y(_02004_),
    .A2(_01998_));
 sg13g2_buf_2 fanout498 (.A(net499),
    .X(net498));
 sg13g2_inv_2 _07272_ (.Y(_02006_),
    .A(net185));
 sg13g2_buf_2 fanout497 (.A(out_select_p2c_1),
    .X(net497));
 sg13g2_buf_2 fanout496 (.A(net497),
    .X(net496));
 sg13g2_nand2_1 _07275_ (.Y(_02009_),
    .A(net73),
    .B(net182));
 sg13g2_nand2_1 _07276_ (.Y(_02010_),
    .A(net59),
    .B(_02009_));
 sg13g2_nand2_1 _07277_ (.Y(_02011_),
    .A(net99),
    .B(_02009_));
 sg13g2_buf_2 fanout495 (.A(out_select_p2c_2),
    .X(net495));
 sg13g2_xor2_1 _07279_ (.B(net183),
    .A(net99),
    .X(_02013_));
 sg13g2_xnor2_1 _07280_ (.Y(_02014_),
    .A(net111),
    .B(net76));
 sg13g2_xnor2_1 _07281_ (.Y(_02015_),
    .A(net110),
    .B(\median_processor.input_storage[9] ));
 sg13g2_nand4_1 _07282_ (.B(_02001_),
    .C(_02014_),
    .A(_01980_),
    .Y(_02016_),
    .D(_02015_));
 sg13g2_nor3_1 _07283_ (.A(_01996_),
    .B(_02013_),
    .C(_02016_),
    .Y(_02017_));
 sg13g2_a221oi_1 _07284_ (.B2(_02011_),
    .C1(_02017_),
    .B1(_02010_),
    .A1(_01997_),
    .Y(_02018_),
    .A2(_02004_));
 sg13g2_buf_2 fanout494 (.A(net495),
    .X(net494));
 sg13g2_nand3_1 _07286_ (.B(net59),
    .C(_02009_),
    .A(net99),
    .Y(_02020_));
 sg13g2_o21ai_1 _07287_ (.B1(_02020_),
    .Y(_02021_),
    .A1(net73),
    .A2(net182));
 sg13g2_or2_1 _07288_ (.X(_02022_),
    .B(_02021_),
    .A(_02018_));
 sg13g2_buf_1 fanout493 (.A(\median_processor.rst ),
    .X(net493));
 sg13g2_buf_1 fanout492 (.A(net493),
    .X(net492));
 sg13g2_buf_1 fanout491 (.A(net492),
    .X(net491));
 sg13g2_buf_2 fanout490 (.A(net491),
    .X(net490));
 sg13g2_buf_2 fanout489 (.A(net491),
    .X(net489));
 sg13g2_buf_2 fanout488 (.A(net489),
    .X(net488));
 sg13g2_nor2b_1 _07295_ (.A(net108),
    .B_N(net150),
    .Y(_02029_));
 sg13g2_nor3_1 _07296_ (.A(net196),
    .B(_02029_),
    .C(_01935_),
    .Y(_02030_));
 sg13g2_nand2b_1 _07297_ (.Y(_02031_),
    .B(net111),
    .A_N(net196));
 sg13g2_buf_2 fanout487 (.A(net491),
    .X(net487));
 sg13g2_a221oi_1 _07299_ (.B2(_02031_),
    .C1(\median_processor.input_storage[1] ),
    .B1(_01885_),
    .A1(net150),
    .Y(_02033_),
    .A2(_01931_));
 sg13g2_buf_1 fanout486 (.A(net492),
    .X(net486));
 sg13g2_nand2b_1 _07301_ (.Y(_02035_),
    .B(net103),
    .A_N(\median_processor.input_storage[4] ));
 sg13g2_o21ai_1 _07302_ (.B1(_02035_),
    .Y(_02036_),
    .A1(net150),
    .A2(_01931_));
 sg13g2_nor4_1 _07303_ (.A(net106),
    .B(_02030_),
    .C(_02033_),
    .D(_02036_),
    .Y(_02037_));
 sg13g2_buf_2 fanout485 (.A(net486),
    .X(net485));
 sg13g2_buf_2 fanout484 (.A(net485),
    .X(net484));
 sg13g2_inv_2 _07306_ (.Y(_02040_),
    .A(net128));
 sg13g2_nor4_1 _07307_ (.A(_02040_),
    .B(_02030_),
    .C(_02033_),
    .D(_02036_),
    .Y(_02041_));
 sg13g2_inv_2 _07308_ (.Y(_02042_),
    .A(net109));
 sg13g2_nand3_1 _07309_ (.B(_01712_),
    .C(_02035_),
    .A(net128),
    .Y(_02043_));
 sg13g2_o21ai_1 _07310_ (.B1(_02043_),
    .Y(_02044_),
    .A1(net58),
    .A2(net103));
 sg13g2_buf_1 fanout483 (.A(net492),
    .X(net483));
 sg13g2_buf_1 fanout482 (.A(net483),
    .X(net482));
 sg13g2_buf_1 fanout481 (.A(net483),
    .X(net481));
 sg13g2_buf_1 fanout480 (.A(net492),
    .X(net480));
 sg13g2_a22oi_1 _07315_ (.Y(_02049_),
    .B1(net72),
    .B2(net80),
    .A2(net73),
    .A1(net77));
 sg13g2_nand2_1 _07316_ (.Y(_02050_),
    .A(net101),
    .B(_02049_));
 sg13g2_nor4_1 _07317_ (.A(_02037_),
    .B(_02041_),
    .C(_02044_),
    .D(_02050_),
    .Y(_02051_));
 sg13g2_buf_1 fanout479 (.A(net480),
    .X(net479));
 sg13g2_inv_2 _07319_ (.Y(_02053_),
    .A(net89));
 sg13g2_nand2_1 _07320_ (.Y(_02054_),
    .A(_02053_),
    .B(_02049_));
 sg13g2_nor4_1 _07321_ (.A(_02037_),
    .B(_02041_),
    .C(_02044_),
    .D(_02054_),
    .Y(_02055_));
 sg13g2_nor2_1 _07322_ (.A(net80),
    .B(net72),
    .Y(_02056_));
 sg13g2_nor2_1 _07323_ (.A(net97),
    .B(_02056_),
    .Y(_02057_));
 sg13g2_inv_1 _07324_ (.Y(_02058_),
    .A(net77));
 sg13g2_a21oi_1 _07325_ (.A1(net97),
    .A2(_02056_),
    .Y(_02059_),
    .B1(net57));
 sg13g2_nand3_1 _07326_ (.B(net101),
    .C(_02049_),
    .A(_02053_),
    .Y(_02060_));
 sg13g2_o21ai_1 _07327_ (.B1(_02060_),
    .Y(_02061_),
    .A1(_02057_),
    .A2(_02059_));
 sg13g2_nor3_1 _07328_ (.A(_02051_),
    .B(_02055_),
    .C(_02061_),
    .Y(_02062_));
 sg13g2_buf_1 fanout478 (.A(net480),
    .X(net478));
 sg13g2_nor2b_1 _07330_ (.A(net26),
    .B_N(_02062_),
    .Y(_02064_));
 sg13g2_nand2b_1 _07331_ (.Y(_02065_),
    .B(net26),
    .A_N(net24));
 sg13g2_nand2b_1 _07332_ (.Y(_02066_),
    .B(_02065_),
    .A_N(_02064_));
 sg13g2_a21oi_1 _07333_ (.A1(_01969_),
    .A2(_01975_),
    .Y(_02067_),
    .B1(_02066_));
 sg13g2_nand2_1 _07334_ (.Y(_02068_),
    .A(_01857_),
    .B(_01858_));
 sg13g2_and2_1 _07335_ (.A(net32),
    .B(net29),
    .X(_02069_));
 sg13g2_and2_1 _07336_ (.A(_01861_),
    .B(_02069_),
    .X(_02070_));
 sg13g2_nor3_1 _07337_ (.A(net31),
    .B(_01852_),
    .C(_01854_),
    .Y(_02071_));
 sg13g2_nor2_1 _07338_ (.A(_01761_),
    .B(net29),
    .Y(_02072_));
 sg13g2_a22oi_1 _07339_ (.Y(_02073_),
    .B1(_02071_),
    .B2(_02072_),
    .A2(_02070_),
    .A1(_02068_));
 sg13g2_o21ai_1 _07340_ (.B1(net31),
    .Y(_02074_),
    .A1(_01852_),
    .A2(_01854_));
 sg13g2_xnor2_1 _07341_ (.Y(_02075_),
    .A(_01859_),
    .B(net29));
 sg13g2_nand3b_1 _07342_ (.B(_02074_),
    .C(_02075_),
    .Y(_02076_),
    .A_N(_02071_));
 sg13g2_nand3b_1 _07343_ (.B(net26),
    .C(net27),
    .Y(_02077_),
    .A_N(net24));
 sg13g2_a21oi_1 _07344_ (.A1(_02073_),
    .A2(_02076_),
    .Y(_02078_),
    .B1(_02077_));
 sg13g2_a21oi_1 _07345_ (.A1(_01761_),
    .A2(net29),
    .Y(_02079_),
    .B1(_01811_));
 sg13g2_o21ai_1 _07346_ (.B1(_02064_),
    .Y(_02080_),
    .A1(_02072_),
    .A2(_02079_));
 sg13g2_xnor2_1 _07347_ (.Y(_02081_),
    .A(net31),
    .B(_02075_));
 sg13g2_nor2_1 _07348_ (.A(_01974_),
    .B(_02081_),
    .Y(_02082_));
 sg13g2_and2_1 _07349_ (.A(_01974_),
    .B(_02081_),
    .X(_02083_));
 sg13g2_nor4_1 _07350_ (.A(_02080_),
    .B(net27),
    .C(_02082_),
    .D(_02083_),
    .Y(_02084_));
 sg13g2_or4_1 _07351_ (.A(_02072_),
    .B(_02079_),
    .C(net28),
    .D(_02065_),
    .X(_02085_));
 sg13g2_a21oi_1 _07352_ (.A1(_02069_),
    .A2(_02071_),
    .Y(_02086_),
    .B1(_02085_));
 sg13g2_nor2b_1 _07353_ (.A(_02080_),
    .B_N(net28),
    .Y(_02087_));
 sg13g2_mux2_1 _07354_ (.A0(_02086_),
    .A1(_02087_),
    .S(_02082_),
    .X(_02088_));
 sg13g2_or4_1 _07355_ (.A(_02067_),
    .B(_02078_),
    .C(_02084_),
    .D(_02088_),
    .X(_02089_));
 sg13g2_buf_1 fanout477 (.A(net480),
    .X(net477));
 sg13g2_buf_1 fanout476 (.A(net480),
    .X(net476));
 sg13g2_buf_1 fanout475 (.A(net492),
    .X(net475));
 sg13g2_nand2b_1 _07359_ (.Y(_02093_),
    .B(net127),
    .A_N(net164));
 sg13g2_o21ai_1 _07360_ (.B1(_02093_),
    .Y(_02094_),
    .A1(net161),
    .A2(net70));
 sg13g2_a22oi_1 _07361_ (.Y(_02095_),
    .B1(_01773_),
    .B2(net162),
    .A2(_01780_),
    .A1(net159));
 sg13g2_nand2b_1 _07362_ (.Y(_02096_),
    .B(net126),
    .A_N(net159));
 sg13g2_nand2b_1 _07363_ (.Y(_02097_),
    .B(net120),
    .A_N(net155));
 sg13g2_nand2b_1 _07364_ (.Y(_02098_),
    .B(net123),
    .A_N(net157));
 sg13g2_nand3_1 _07365_ (.B(_02097_),
    .C(_02098_),
    .A(_02096_),
    .Y(_02099_));
 sg13g2_a21oi_1 _07366_ (.A1(_02094_),
    .A2(_02095_),
    .Y(_02100_),
    .B1(_02099_));
 sg13g2_a221oi_1 _07367_ (.B2(net157),
    .C1(net155),
    .B1(_01781_),
    .A1(net152),
    .Y(_02101_),
    .A2(net68));
 sg13g2_nor2b_1 _07368_ (.A(net124),
    .B_N(net157),
    .Y(_02102_));
 sg13g2_inv_1 _07369_ (.Y(_02103_),
    .A(net122));
 sg13g2_a221oi_1 _07370_ (.B2(net155),
    .C1(_02103_),
    .B1(_02102_),
    .A1(net152),
    .Y(_02104_),
    .A2(net68));
 sg13g2_o21ai_1 _07371_ (.B1(net114),
    .Y(_02105_),
    .A1(_02101_),
    .A2(_02104_));
 sg13g2_nor2_1 _07372_ (.A(net152),
    .B(_01796_),
    .Y(_02106_));
 sg13g2_inv_1 _07373_ (.Y(_02107_),
    .A(net148));
 sg13g2_a21oi_1 _07374_ (.A1(net114),
    .A2(_02106_),
    .Y(_02108_),
    .B1(_02107_));
 sg13g2_o21ai_1 _07375_ (.B1(_02108_),
    .Y(_02109_),
    .A1(_02100_),
    .A2(_02105_));
 sg13g2_nor2_1 _07376_ (.A(net114),
    .B(_02106_),
    .Y(_02110_));
 sg13g2_nor2_1 _07377_ (.A(_02101_),
    .B(_02104_),
    .Y(_02111_));
 sg13g2_nand2_1 _07378_ (.Y(_02112_),
    .A(_02094_),
    .B(_02095_));
 sg13g2_nor3_1 _07379_ (.A(net114),
    .B(_02106_),
    .C(_02099_),
    .Y(_02113_));
 sg13g2_a221oi_1 _07380_ (.B2(_02113_),
    .C1(net71),
    .B1(_02112_),
    .A1(_02110_),
    .Y(_02114_),
    .A2(_02111_));
 sg13g2_a21oi_1 _07381_ (.A1(_02109_),
    .A2(_02114_),
    .Y(_02115_),
    .B1(_01759_));
 sg13g2_nor2_1 _07382_ (.A(net113),
    .B(net116),
    .Y(_02116_));
 sg13g2_or2_1 _07383_ (.X(_02117_),
    .B(_02100_),
    .A(_02111_));
 sg13g2_inv_1 _07384_ (.Y(_02118_),
    .A(net117));
 sg13g2_nor2_1 _07385_ (.A(net148),
    .B(_02118_),
    .Y(_02119_));
 sg13g2_nor3_1 _07386_ (.A(net113),
    .B(_02106_),
    .C(_02119_),
    .Y(_02120_));
 sg13g2_a22oi_1 _07387_ (.Y(_02121_),
    .B1(_02117_),
    .B2(_02120_),
    .A2(_02116_),
    .A1(net148));
 sg13g2_nor2b_1 _07388_ (.A(_02115_),
    .B_N(_02121_),
    .Y(_02122_));
 sg13g2_nor2b_1 _07389_ (.A(net166),
    .B_N(\median_processor.input_storage[47] ),
    .Y(_02123_));
 sg13g2_a21oi_1 _07390_ (.A1(net172),
    .A2(_02103_),
    .Y(_02124_),
    .B1(net68));
 sg13g2_a21oi_1 _07391_ (.A1(net172),
    .A2(_01794_),
    .Y(_02125_),
    .B1(net169));
 sg13g2_o21ai_1 _07392_ (.B1(net115),
    .Y(_02126_),
    .A1(_02124_),
    .A2(_02125_));
 sg13g2_nor3_1 _07393_ (.A(net114),
    .B(_02124_),
    .C(_02125_),
    .Y(_02127_));
 sg13g2_a21oi_1 _07394_ (.A1(net167),
    .A2(_02126_),
    .Y(_02128_),
    .B1(_02127_));
 sg13g2_nand2b_1 _07395_ (.Y(_02129_),
    .B(net119),
    .A_N(net169));
 sg13g2_a21oi_1 _07396_ (.A1(_02118_),
    .A2(_02129_),
    .Y(_02130_),
    .B1(net167));
 sg13g2_nand2b_1 _07397_ (.Y(_02131_),
    .B(net125),
    .A_N(net176));
 sg13g2_a21oi_1 _07398_ (.A1(net69),
    .A2(_02131_),
    .Y(_02132_),
    .B1(net173));
 sg13g2_nand2_1 _07399_ (.Y(_02133_),
    .A(net117),
    .B(net118));
 sg13g2_nor2_1 _07400_ (.A(net170),
    .B(_02133_),
    .Y(_02134_));
 sg13g2_nand3b_1 _07401_ (.B(net123),
    .C(net126),
    .Y(_02135_),
    .A_N(net176));
 sg13g2_nand2b_1 _07402_ (.Y(_02136_),
    .B(net120),
    .A_N(net172));
 sg13g2_nand3b_1 _07403_ (.B(_02135_),
    .C(_02136_),
    .Y(_02137_),
    .A_N(_02123_));
 sg13g2_nor4_1 _07404_ (.A(_02130_),
    .B(_02132_),
    .C(_02134_),
    .D(_02137_),
    .Y(_02138_));
 sg13g2_a22oi_1 _07405_ (.Y(_02139_),
    .B1(_01780_),
    .B2(net175),
    .A2(net69),
    .A1(net173));
 sg13g2_inv_1 _07406_ (.Y(_02140_),
    .A(net127));
 sg13g2_o21ai_1 _07407_ (.B1(net70),
    .Y(_02141_),
    .A1(net178),
    .A2(_02140_));
 sg13g2_nand2_1 _07408_ (.Y(_02142_),
    .A(\median_processor.input_storage[41] ),
    .B(net127));
 sg13g2_o21ai_1 _07409_ (.B1(\median_processor.input_storage[17] ),
    .Y(_02143_),
    .A1(net178),
    .A2(_02142_));
 sg13g2_nand3_1 _07410_ (.B(_02141_),
    .C(_02143_),
    .A(_02139_),
    .Y(_02144_));
 sg13g2_a22oi_1 _07411_ (.Y(_02145_),
    .B1(_02138_),
    .B2(_02144_),
    .A2(net71),
    .A1(net165));
 sg13g2_o21ai_1 _07412_ (.B1(_02145_),
    .Y(_02146_),
    .A1(_02123_),
    .A2(_02128_));
 sg13g2_buf_2 fanout474 (.A(net475),
    .X(net474));
 sg13g2_nand2_1 _07414_ (.Y(_02148_),
    .A(net31),
    .B(_02146_));
 sg13g2_nor2_1 _07415_ (.A(net31),
    .B(_02146_),
    .Y(_02149_));
 sg13g2_a21oi_1 _07416_ (.A1(_02122_),
    .A2(_02148_),
    .Y(_02150_),
    .B1(_02149_));
 sg13g2_nand3_1 _07417_ (.B(net121),
    .C(net123),
    .A(net62),
    .Y(_02151_));
 sg13g2_a21oi_1 _07418_ (.A1(net62),
    .A2(net123),
    .Y(_02152_),
    .B1(net121));
 sg13g2_a21oi_1 _07419_ (.A1(net137),
    .A2(_02151_),
    .Y(_02153_),
    .B1(_02152_));
 sg13g2_inv_4 _07420_ (.A(net135),
    .Y(_02154_));
 sg13g2_buf_1 fanout473 (.A(net474),
    .X(net473));
 sg13g2_nor2_1 _07422_ (.A(net130),
    .B(_01765_),
    .Y(_02156_));
 sg13g2_a221oi_1 _07423_ (.B2(_02154_),
    .C1(_02156_),
    .B1(net119),
    .A1(net61),
    .Y(_02157_),
    .A2(net114));
 sg13g2_nor2b_1 _07424_ (.A(_02153_),
    .B_N(_02157_),
    .Y(_02158_));
 sg13g2_o21ai_1 _07425_ (.B1(net70),
    .Y(_02159_),
    .A1(net144),
    .A2(_02140_));
 sg13g2_o21ai_1 _07426_ (.B1(net143),
    .Y(_02160_),
    .A1(net144),
    .A2(_02142_));
 sg13g2_a22oi_1 _07427_ (.Y(_02161_),
    .B1(_02159_),
    .B2(_02160_),
    .A2(net125),
    .A1(_01918_));
 sg13g2_a22oi_1 _07428_ (.Y(_02162_),
    .B1(_01780_),
    .B2(net140),
    .A2(_01781_),
    .A1(net138));
 sg13g2_o21ai_1 _07429_ (.B1(_02162_),
    .Y(_02163_),
    .A1(_01941_),
    .A2(net120));
 sg13g2_or2_1 _07430_ (.X(_02164_),
    .B(_02163_),
    .A(_02161_));
 sg13g2_nand2b_1 _07431_ (.Y(_02165_),
    .B(net135),
    .A_N(net118));
 sg13g2_nand2_1 _07432_ (.Y(_02166_),
    .A(net114),
    .B(_02165_));
 sg13g2_o21ai_1 _07433_ (.B1(net61),
    .Y(_02167_),
    .A1(net114),
    .A2(_02165_));
 sg13g2_a22oi_1 _07434_ (.Y(_02168_),
    .B1(_02166_),
    .B2(_02167_),
    .A2(net71),
    .A1(net131));
 sg13g2_nor2_1 _07435_ (.A(_02156_),
    .B(_02168_),
    .Y(_02169_));
 sg13g2_a21oi_2 _07436_ (.B1(_02169_),
    .Y(_02170_),
    .A2(_02164_),
    .A1(_02158_));
 sg13g2_buf_2 fanout472 (.A(net475),
    .X(net472));
 sg13g2_or2_1 _07438_ (.X(_02172_),
    .B(_02142_),
    .A(net196));
 sg13g2_nor2b_1 _07439_ (.A(net196),
    .B_N(net127),
    .Y(_02173_));
 sg13g2_inv_2 _07440_ (.Y(_02174_),
    .A(\median_processor.input_storage[1] ));
 sg13g2_o21ai_1 _07441_ (.B1(_02174_),
    .Y(_02175_),
    .A1(\median_processor.input_storage[41] ),
    .A2(_02173_));
 sg13g2_inv_2 _07442_ (.Y(_02176_),
    .A(net151));
 sg13g2_nor2_1 _07443_ (.A(_02176_),
    .B(net125),
    .Y(_02177_));
 sg13g2_a221oi_1 _07444_ (.B2(_02175_),
    .C1(_02177_),
    .B1(_02172_),
    .A1(net128),
    .Y(_02178_),
    .A2(net69));
 sg13g2_nor2b_1 _07445_ (.A(net150),
    .B_N(net126),
    .Y(_02179_));
 sg13g2_o21ai_1 _07446_ (.B1(_02179_),
    .Y(_02180_),
    .A1(_02040_),
    .A2(net123));
 sg13g2_o21ai_1 _07447_ (.B1(_02180_),
    .Y(_02181_),
    .A1(net128),
    .A2(_01781_));
 sg13g2_o21ai_1 _07448_ (.B1(net122),
    .Y(_02182_),
    .A1(_02178_),
    .A2(_02181_));
 sg13g2_nor3_1 _07449_ (.A(net122),
    .B(_02178_),
    .C(_02181_),
    .Y(_02183_));
 sg13g2_a21o_1 _07450_ (.A2(_02182_),
    .A1(net109),
    .B1(_02183_),
    .X(_02184_));
 sg13g2_inv_2 _07451_ (.Y(_02185_),
    .A(net81));
 sg13g2_nor2_1 _07452_ (.A(net77),
    .B(net71),
    .Y(_02186_));
 sg13g2_a221oi_1 _07453_ (.B2(_02053_),
    .C1(_02186_),
    .B1(net118),
    .A1(_02185_),
    .Y(_02187_),
    .A2(net117));
 sg13g2_nand2_1 _07454_ (.Y(_02188_),
    .A(net89),
    .B(net68));
 sg13g2_o21ai_1 _07455_ (.B1(net56),
    .Y(_02189_),
    .A1(net117),
    .A2(_02188_));
 sg13g2_nand2_1 _07456_ (.Y(_02190_),
    .A(net117),
    .B(_02188_));
 sg13g2_a22oi_1 _07457_ (.Y(_02191_),
    .B1(_02189_),
    .B2(_02190_),
    .A2(net71),
    .A1(net77));
 sg13g2_nor2_1 _07458_ (.A(_02186_),
    .B(_02191_),
    .Y(_02192_));
 sg13g2_a21o_1 _07459_ (.A2(_02187_),
    .A1(_02184_),
    .B1(_02192_),
    .X(_02193_));
 sg13g2_buf_1 fanout471 (.A(net472),
    .X(net471));
 sg13g2_inv_1 _07461_ (.Y(_02195_),
    .A(net82));
 sg13g2_nor2b_1 _07462_ (.A(net96),
    .B_N(net127),
    .Y(_02196_));
 sg13g2_nor2_1 _07463_ (.A(_01832_),
    .B(_02196_),
    .Y(_02197_));
 sg13g2_a21oi_1 _07464_ (.A1(_01832_),
    .A2(_02196_),
    .Y(_02198_),
    .B1(\median_processor.input_storage[41] ));
 sg13g2_nand2b_1 _07465_ (.Y(_02199_),
    .B(net126),
    .A_N(net92));
 sg13g2_o21ai_1 _07466_ (.B1(_02199_),
    .Y(_02200_),
    .A1(_02197_),
    .A2(_02198_));
 sg13g2_buf_1 fanout470 (.A(net493),
    .X(net470));
 sg13g2_nand2b_1 _07468_ (.Y(_02202_),
    .B(net92),
    .A_N(net126));
 sg13g2_nand2b_1 _07469_ (.Y(_02203_),
    .B(net90),
    .A_N(net123));
 sg13g2_nand2b_1 _07470_ (.Y(_02204_),
    .B(\median_processor.input_storage[61] ),
    .A_N(net118));
 sg13g2_nand2b_1 _07471_ (.Y(_02205_),
    .B(net87),
    .A_N(net120));
 sg13g2_nand4_1 _07472_ (.B(_02203_),
    .C(_02204_),
    .A(_02202_),
    .Y(_02206_),
    .D(_02205_));
 sg13g2_nor2_1 _07473_ (.A(net85),
    .B(_02206_),
    .Y(_02207_));
 sg13g2_a221oi_1 _07474_ (.B2(_02207_),
    .C1(\median_processor.input_storage[47] ),
    .B1(_02200_),
    .A1(net66),
    .Y(_02208_),
    .A2(net115));
 sg13g2_a221oi_1 _07475_ (.B2(_02207_),
    .C1(_02195_),
    .B1(_02200_),
    .A1(net66),
    .Y(_02209_),
    .A2(net115));
 sg13g2_nor2_1 _07476_ (.A(_02118_),
    .B(_02206_),
    .Y(_02210_));
 sg13g2_nor2b_1 _07477_ (.A(net90),
    .B_N(net123),
    .Y(_02211_));
 sg13g2_a21oi_1 _07478_ (.A1(net120),
    .A2(_02211_),
    .Y(_02212_),
    .B1(net64));
 sg13g2_a21oi_1 _07479_ (.A1(net120),
    .A2(_02211_),
    .Y(_02213_),
    .B1(net118));
 sg13g2_inv_2 _07480_ (.Y(_02214_),
    .A(net87));
 sg13g2_o21ai_1 _07481_ (.B1(_02214_),
    .Y(_02215_),
    .A1(net120),
    .A2(_02211_));
 sg13g2_o21ai_1 _07482_ (.B1(_02215_),
    .Y(_02216_),
    .A1(_02212_),
    .A2(_02213_));
 sg13g2_a22oi_1 _07483_ (.Y(_02217_),
    .B1(_01796_),
    .B2(\median_processor.input_storage[61] ),
    .A2(_02118_),
    .A1(net84));
 sg13g2_nand2b_1 _07484_ (.Y(_02218_),
    .B(net120),
    .A_N(net87));
 sg13g2_nand2b_1 _07485_ (.Y(_02219_),
    .B(net119),
    .A_N(net86));
 sg13g2_nand3_1 _07486_ (.B(_02218_),
    .C(_02219_),
    .A(_02199_),
    .Y(_02220_));
 sg13g2_nand2b_1 _07487_ (.Y(_02221_),
    .B(net96),
    .A_N(net127));
 sg13g2_xnor2_1 _07488_ (.Y(_02222_),
    .A(net94),
    .B(\median_processor.input_storage[41] ));
 sg13g2_nand3b_1 _07489_ (.B(_02221_),
    .C(_02222_),
    .Y(_02223_),
    .A_N(_02196_));
 sg13g2_nor2b_1 _07490_ (.A(net82),
    .B_N(net113),
    .Y(_02224_));
 sg13g2_xor2_1 _07491_ (.B(net117),
    .A(net84),
    .X(_02225_));
 sg13g2_or3_1 _07492_ (.A(_02224_),
    .B(_02211_),
    .C(_02225_),
    .X(_02226_));
 sg13g2_nor4_1 _07493_ (.A(_02206_),
    .B(_02220_),
    .C(_02223_),
    .D(_02226_),
    .Y(_02227_));
 sg13g2_a221oi_1 _07494_ (.B2(_02217_),
    .C1(_02227_),
    .B1(_02216_),
    .A1(_02200_),
    .Y(_02228_),
    .A2(_02210_));
 sg13g2_o21ai_1 _07495_ (.B1(_02228_),
    .Y(_02229_),
    .A1(_02208_),
    .A2(_02209_));
 sg13g2_o21ai_1 _07496_ (.B1(_02229_),
    .Y(_02230_),
    .A1(_02195_),
    .A2(net113));
 sg13g2_buf_2 fanout469 (.A(net470),
    .X(net469));
 sg13g2_xnor2_1 _07498_ (.Y(_02232_),
    .A(_02193_),
    .B(_02230_));
 sg13g2_nor3_1 _07499_ (.A(_02150_),
    .B(_02170_),
    .C(_02232_),
    .Y(_02233_));
 sg13g2_and3_1 _07500_ (.X(_02234_),
    .A(net20),
    .B(_02230_),
    .C(_02170_));
 sg13g2_inv_1 _07501_ (.Y(_02235_),
    .A(_02170_));
 sg13g2_nor3_1 _07502_ (.A(net20),
    .B(_02230_),
    .C(_02235_),
    .Y(_02236_));
 sg13g2_mux2_1 _07503_ (.A0(_02234_),
    .A1(_02236_),
    .S(_02150_),
    .X(_02237_));
 sg13g2_nand2_1 _07504_ (.Y(_02238_),
    .A(net191),
    .B(net69));
 sg13g2_o21ai_1 _07505_ (.B1(net70),
    .Y(_02239_),
    .A1(\median_processor.input_storage[8] ),
    .A2(_02140_));
 sg13g2_o21ai_1 _07506_ (.B1(net74),
    .Y(_02240_),
    .A1(net76),
    .A2(_02142_));
 sg13g2_a21oi_1 _07507_ (.A1(_02239_),
    .A2(_02240_),
    .Y(_02241_),
    .B1(net125));
 sg13g2_nand3_1 _07508_ (.B(_02239_),
    .C(_02240_),
    .A(net125),
    .Y(_02242_));
 sg13g2_o21ai_1 _07509_ (.B1(_02242_),
    .Y(_02243_),
    .A1(net195),
    .A2(_02241_));
 sg13g2_nor2_1 _07510_ (.A(net192),
    .B(net69),
    .Y(_02244_));
 sg13g2_a21oi_1 _07511_ (.A1(_02238_),
    .A2(_02243_),
    .Y(_02245_),
    .B1(_02244_));
 sg13g2_o21ai_1 _07512_ (.B1(net113),
    .Y(_02246_),
    .A1(net59),
    .A2(net117));
 sg13g2_a21o_1 _07513_ (.A2(_02116_),
    .A1(net183),
    .B1(net180),
    .X(_02247_));
 sg13g2_a22oi_1 _07514_ (.Y(_02248_),
    .B1(_02246_),
    .B2(_02247_),
    .A2(net68),
    .A1(net186));
 sg13g2_o21ai_1 _07515_ (.B1(_02248_),
    .Y(_02249_),
    .A1(_01999_),
    .A2(net122));
 sg13g2_inv_1 _07516_ (.Y(_02250_),
    .A(net181));
 sg13g2_buf_2 fanout468 (.A(net469),
    .X(net468));
 sg13g2_nor2_1 _07518_ (.A(net190),
    .B(_02103_),
    .Y(_02252_));
 sg13g2_o21ai_1 _07519_ (.B1(_02118_),
    .Y(_02253_),
    .A1(net186),
    .A2(net68));
 sg13g2_o21ai_1 _07520_ (.B1(net183),
    .Y(_02254_),
    .A1(net187),
    .A2(_02133_));
 sg13g2_nand2_1 _07521_ (.Y(_02255_),
    .A(_02253_),
    .B(_02254_));
 sg13g2_a21oi_1 _07522_ (.A1(net180),
    .A2(net71),
    .Y(_02256_),
    .B1(_02255_));
 sg13g2_a221oi_1 _07523_ (.B2(_02252_),
    .C1(_02256_),
    .B1(_02248_),
    .A1(net55),
    .Y(_02257_),
    .A2(net113));
 sg13g2_o21ai_1 _07524_ (.B1(_02257_),
    .Y(_02258_),
    .A1(_02245_),
    .A2(_02249_));
 sg13g2_buf_2 fanout467 (.A(net468),
    .X(net467));
 sg13g2_xnor2_1 _07526_ (.Y(_02260_),
    .A(_01811_),
    .B(_02258_));
 sg13g2_nand2b_2 _07527_ (.Y(_02261_),
    .B(_02121_),
    .A_N(_02115_));
 sg13g2_buf_1 fanout466 (.A(net467),
    .X(net466));
 sg13g2_xnor2_1 _07529_ (.Y(_02263_),
    .A(_02146_),
    .B(_02261_));
 sg13g2_xor2_1 _07530_ (.B(_02263_),
    .A(_02260_),
    .X(_02264_));
 sg13g2_o21ai_1 _07531_ (.B1(_02264_),
    .Y(_02265_),
    .A1(_02233_),
    .A2(_02237_));
 sg13g2_or2_1 _07532_ (.X(_02266_),
    .B(_02263_),
    .A(_02260_));
 sg13g2_nor3_1 _07533_ (.A(net19),
    .B(_02146_),
    .C(_02261_),
    .Y(_02267_));
 sg13g2_and2_1 _07534_ (.A(_01811_),
    .B(_02258_),
    .X(_02268_));
 sg13g2_inv_1 _07535_ (.Y(_02269_),
    .A(_02146_));
 sg13g2_nor2_1 _07536_ (.A(_02269_),
    .B(_02122_),
    .Y(_02270_));
 sg13g2_a22oi_1 _07537_ (.Y(_02271_),
    .B1(_02268_),
    .B2(_02270_),
    .A2(_02267_),
    .A1(net31));
 sg13g2_or2_1 _07538_ (.X(_02272_),
    .B(_02230_),
    .A(_02193_));
 sg13g2_mux2_1 _07539_ (.A0(_02232_),
    .A1(_02272_),
    .S(_02235_),
    .X(_02273_));
 sg13g2_a21o_1 _07540_ (.A2(_02271_),
    .A1(_02266_),
    .B1(_02273_),
    .X(_02274_));
 sg13g2_nor3_1 _07541_ (.A(_02146_),
    .B(_02261_),
    .C(_02170_),
    .Y(_02275_));
 sg13g2_nand4_1 _07542_ (.B(_02230_),
    .C(_02268_),
    .A(net20),
    .Y(_02276_),
    .D(_02275_));
 sg13g2_nand3_1 _07543_ (.B(_02274_),
    .C(_02276_),
    .A(_02265_),
    .Y(_02277_));
 sg13g2_buf_2 fanout465 (.A(net467),
    .X(net465));
 sg13g2_nand2_1 _07545_ (.Y(_02279_),
    .A(net127),
    .B(net11));
 sg13g2_nand2_1 _07546_ (.Y(_02280_),
    .A(net111),
    .B(net12));
 sg13g2_o21ai_1 _07547_ (.B1(_02280_),
    .Y(_02281_),
    .A1(net12),
    .A2(_02279_));
 sg13g2_nor2b_1 _07548_ (.A(net75),
    .B_N(net96),
    .Y(_02282_));
 sg13g2_o21ai_1 _07549_ (.B1(net94),
    .Y(_02283_),
    .A1(_01985_),
    .A2(_02282_));
 sg13g2_inv_2 _07550_ (.Y(_02284_),
    .A(net193));
 sg13g2_a221oi_1 _07551_ (.B2(_02282_),
    .C1(_02284_),
    .B1(_01985_),
    .A1(net92),
    .Y(_02285_),
    .A2(net60));
 sg13g2_nand2b_1 _07552_ (.Y(_02286_),
    .B(net194),
    .A_N(net92));
 sg13g2_a21oi_1 _07553_ (.A1(net91),
    .A2(_02284_),
    .Y(_02287_),
    .B1(_02286_));
 sg13g2_a21o_1 _07554_ (.A2(_02285_),
    .A1(_02283_),
    .B1(_02287_),
    .X(_02288_));
 sg13g2_a221oi_1 _07555_ (.B2(_02282_),
    .C1(net91),
    .B1(_01985_),
    .A1(net92),
    .Y(_02289_),
    .A2(net60));
 sg13g2_nor2_1 _07556_ (.A(net91),
    .B(_02284_),
    .Y(_02290_));
 sg13g2_a21o_1 _07557_ (.A2(_02289_),
    .A1(_02283_),
    .B1(_02290_),
    .X(_02291_));
 sg13g2_nor2b_1 _07558_ (.A(net87),
    .B_N(net189),
    .Y(_02292_));
 sg13g2_o21ai_1 _07559_ (.B1(net65),
    .Y(_02293_),
    .A1(net188),
    .A2(_02292_));
 sg13g2_buf_1 fanout464 (.A(net470),
    .X(net464));
 sg13g2_nand2_1 _07561_ (.Y(_02295_),
    .A(net188),
    .B(_02292_));
 sg13g2_nand2b_1 _07562_ (.Y(_02296_),
    .B(net180),
    .A_N(net83));
 sg13g2_and2_1 _07563_ (.A(net59),
    .B(_02296_),
    .X(_02297_));
 sg13g2_nand3_1 _07564_ (.B(_02295_),
    .C(_02297_),
    .A(_02293_),
    .Y(_02298_));
 sg13g2_nor3_1 _07565_ (.A(_02288_),
    .B(_02291_),
    .C(_02298_),
    .Y(_02299_));
 sg13g2_and2_1 _07566_ (.A(net84),
    .B(_02296_),
    .X(_02300_));
 sg13g2_nand3_1 _07567_ (.B(_02295_),
    .C(_02300_),
    .A(_02293_),
    .Y(_02301_));
 sg13g2_nor3_1 _07568_ (.A(_02288_),
    .B(_02291_),
    .C(_02301_),
    .Y(_02302_));
 sg13g2_nand2b_1 _07569_ (.Y(_02303_),
    .B(net87),
    .A_N(net190));
 sg13g2_o21ai_1 _07570_ (.B1(_02303_),
    .Y(_02304_),
    .A1(net65),
    .A2(net188));
 sg13g2_nand4_1 _07571_ (.B(_02295_),
    .C(_02304_),
    .A(_02293_),
    .Y(_02305_),
    .D(_02297_));
 sg13g2_nand4_1 _07572_ (.B(_02295_),
    .C(_02304_),
    .A(_02293_),
    .Y(_02306_),
    .D(_02300_));
 sg13g2_nand3_1 _07573_ (.B(net59),
    .C(_02296_),
    .A(net84),
    .Y(_02307_));
 sg13g2_nand3_1 _07574_ (.B(_02306_),
    .C(_02307_),
    .A(_02305_),
    .Y(_02308_));
 sg13g2_nand2_1 _07575_ (.Y(_02309_),
    .A(net83),
    .B(net55));
 sg13g2_inv_1 _07576_ (.Y(_02310_),
    .A(_02309_));
 sg13g2_or4_2 _07577_ (.A(_02299_),
    .B(_02302_),
    .C(_02308_),
    .D(_02310_),
    .X(_02311_));
 sg13g2_buf_2 fanout463 (.A(net464),
    .X(net463));
 sg13g2_nor2_1 _07579_ (.A(_02040_),
    .B(net91),
    .Y(_02313_));
 sg13g2_nor2b_1 _07580_ (.A(net196),
    .B_N(net95),
    .Y(_02314_));
 sg13g2_o21ai_1 _07581_ (.B1(\median_processor.input_storage[1] ),
    .Y(_02315_),
    .A1(net196),
    .A2(_01828_));
 sg13g2_o21ai_1 _07582_ (.B1(_02315_),
    .Y(_02316_),
    .A1(net94),
    .A2(_02314_));
 sg13g2_a21oi_1 _07583_ (.A1(net151),
    .A2(_01831_),
    .Y(_02317_),
    .B1(_02316_));
 sg13g2_a221oi_1 _07584_ (.B2(_02176_),
    .C1(_02317_),
    .B1(net93),
    .A1(_02040_),
    .Y(_02318_),
    .A2(net90));
 sg13g2_nand2_1 _07585_ (.Y(_02319_),
    .A(net77),
    .B(_02195_));
 sg13g2_a22oi_1 _07586_ (.Y(_02320_),
    .B1(net64),
    .B2(net89),
    .A2(net67),
    .A1(net80));
 sg13g2_nand2_1 _07587_ (.Y(_02321_),
    .A(net109),
    .B(_02214_));
 sg13g2_nand3_1 _07588_ (.B(_02320_),
    .C(_02321_),
    .A(_02319_),
    .Y(_02322_));
 sg13g2_nor3_1 _07589_ (.A(_02313_),
    .B(_02318_),
    .C(_02322_),
    .Y(_02323_));
 sg13g2_nand2_1 _07590_ (.Y(_02324_),
    .A(_02053_),
    .B(net86));
 sg13g2_o21ai_1 _07591_ (.B1(net80),
    .Y(_02325_),
    .A1(net66),
    .A2(_02324_));
 sg13g2_nand2_1 _07592_ (.Y(_02326_),
    .A(net66),
    .B(_02324_));
 sg13g2_nand2_1 _07593_ (.Y(_02327_),
    .A(_02325_),
    .B(_02326_));
 sg13g2_o21ai_1 _07594_ (.B1(_02327_),
    .Y(_02328_),
    .A1(net77),
    .A2(_02195_));
 sg13g2_and3_1 _07595_ (.X(_02329_),
    .A(net58),
    .B(net88),
    .C(_02319_));
 sg13g2_a22oi_1 _07596_ (.Y(_02330_),
    .B1(_02320_),
    .B2(_02329_),
    .A2(_02328_),
    .A1(_02319_));
 sg13g2_nand2b_1 _07597_ (.Y(_02331_),
    .B(_02330_),
    .A_N(_02323_));
 sg13g2_and2_1 _07598_ (.A(_02311_),
    .B(_02331_),
    .X(_02332_));
 sg13g2_buf_1 fanout462 (.A(net463),
    .X(net462));
 sg13g2_inv_2 _07600_ (.Y(_02334_),
    .A(_02230_));
 sg13g2_nor2b_1 _07601_ (.A(net90),
    .B_N(net139),
    .Y(_02335_));
 sg13g2_nand2_1 _07602_ (.Y(_02336_),
    .A(_02214_),
    .B(_02335_));
 sg13g2_o21ai_1 _07603_ (.B1(net136),
    .Y(_02337_),
    .A1(_02214_),
    .A2(_02335_));
 sg13g2_nand2_1 _07604_ (.Y(_02338_),
    .A(_02336_),
    .B(_02337_));
 sg13g2_a221oi_1 _07605_ (.B2(_02154_),
    .C1(net82),
    .B1(net86),
    .A1(_01945_),
    .Y(_02339_),
    .A2(net85));
 sg13g2_nand2b_1 _07606_ (.Y(_02340_),
    .B(net88),
    .A_N(net136));
 sg13g2_nand2b_1 _07607_ (.Y(_02341_),
    .B(net91),
    .A_N(net139));
 sg13g2_nand2b_1 _07608_ (.Y(_02342_),
    .B(net93),
    .A_N(net141));
 sg13g2_nand3_1 _07609_ (.B(_02341_),
    .C(_02342_),
    .A(_02340_),
    .Y(_02343_));
 sg13g2_nor2b_1 _07610_ (.A(_02343_),
    .B_N(_02339_),
    .Y(_02344_));
 sg13g2_nand2b_1 _07611_ (.Y(_02345_),
    .B(net95),
    .A_N(net144));
 sg13g2_o21ai_1 _07612_ (.B1(_02345_),
    .Y(_02346_),
    .A1(net142),
    .A2(_01832_));
 sg13g2_a22oi_1 _07613_ (.Y(_02347_),
    .B1(_01832_),
    .B2(net142),
    .A2(_01831_),
    .A1(net141));
 sg13g2_nand2_1 _07614_ (.Y(_02348_),
    .A(_02346_),
    .B(_02347_));
 sg13g2_nor2b_1 _07615_ (.A(net86),
    .B_N(net134),
    .Y(_02349_));
 sg13g2_a21oi_1 _07616_ (.A1(net66),
    .A2(_02349_),
    .Y(_02350_),
    .B1(net132));
 sg13g2_nor2_1 _07617_ (.A(net66),
    .B(_02349_),
    .Y(_02351_));
 sg13g2_nor3_1 _07618_ (.A(net82),
    .B(_02350_),
    .C(_02351_),
    .Y(_02352_));
 sg13g2_a221oi_1 _07619_ (.B2(_02348_),
    .C1(_02352_),
    .B1(_02344_),
    .A1(_02338_),
    .Y(_02353_),
    .A2(_02339_));
 sg13g2_nand2b_1 _07620_ (.Y(_02354_),
    .B(net86),
    .A_N(net134));
 sg13g2_o21ai_1 _07621_ (.B1(_02354_),
    .Y(_02355_),
    .A1(net132),
    .A2(net66));
 sg13g2_inv_1 _07622_ (.Y(_02356_),
    .A(_02355_));
 sg13g2_nor2_1 _07623_ (.A(_02355_),
    .B(_02343_),
    .Y(_02357_));
 sg13g2_o21ai_1 _07624_ (.B1(net82),
    .Y(_02358_),
    .A1(_02350_),
    .A2(_02351_));
 sg13g2_a221oi_1 _07625_ (.B2(_02357_),
    .C1(_02358_),
    .B1(_02348_),
    .A1(_02356_),
    .Y(_02359_),
    .A2(_02338_));
 sg13g2_a21oi_2 _07626_ (.B1(_02359_),
    .Y(_02360_),
    .A2(_02353_),
    .A1(_01922_));
 sg13g2_buf_1 fanout461 (.A(net464),
    .X(net461));
 sg13g2_nor2_2 _07628_ (.A(_02334_),
    .B(_02360_),
    .Y(_02362_));
 sg13g2_nor2b_1 _07629_ (.A(_02230_),
    .B_N(_02360_),
    .Y(_02363_));
 sg13g2_inv_2 _07630_ (.Y(_02364_),
    .A(net167));
 sg13g2_nand2_1 _07631_ (.Y(_02365_),
    .A(net64),
    .B(net169));
 sg13g2_nand2_1 _07632_ (.Y(_02366_),
    .A(net90),
    .B(_01895_));
 sg13g2_nor2_1 _07633_ (.A(_01831_),
    .B(net176),
    .Y(_02367_));
 sg13g2_nand2b_1 _07634_ (.Y(_02368_),
    .B(net95),
    .A_N(net179));
 sg13g2_nand3b_1 _07635_ (.B(net95),
    .C(net94),
    .Y(_02369_),
    .A_N(net179));
 sg13g2_a22oi_1 _07636_ (.Y(_02370_),
    .B1(_02369_),
    .B2(net177),
    .A2(_02368_),
    .A1(_01832_));
 sg13g2_a22oi_1 _07637_ (.Y(_02371_),
    .B1(net176),
    .B2(_01831_),
    .A2(net174),
    .A1(_01835_));
 sg13g2_o21ai_1 _07638_ (.B1(_02371_),
    .Y(_02372_),
    .A1(_02367_),
    .A2(_02370_));
 sg13g2_a22oi_1 _07639_ (.Y(_02373_),
    .B1(_02366_),
    .B2(_02372_),
    .A2(net171),
    .A1(_02214_));
 sg13g2_a21o_1 _07640_ (.A2(_01877_),
    .A1(net88),
    .B1(_02373_),
    .X(_02374_));
 sg13g2_inv_2 _07641_ (.Y(_02375_),
    .A(net165));
 sg13g2_buf_1 fanout460 (.A(net461),
    .X(net460));
 sg13g2_nand2_1 _07643_ (.Y(_02377_),
    .A(net82),
    .B(net54));
 sg13g2_o21ai_1 _07644_ (.B1(_02377_),
    .Y(_02378_),
    .A1(net64),
    .A2(net169));
 sg13g2_a221oi_1 _07645_ (.B2(_02374_),
    .C1(_02378_),
    .B1(_02365_),
    .A1(net85),
    .Y(_02379_),
    .A2(_02364_));
 sg13g2_nand3_1 _07646_ (.B(net168),
    .C(_02377_),
    .A(net67),
    .Y(_02380_));
 sg13g2_o21ai_1 _07647_ (.B1(_02380_),
    .Y(_02381_),
    .A1(net82),
    .A2(net54));
 sg13g2_or2_1 _07648_ (.X(_02382_),
    .B(_02381_),
    .A(_02379_));
 sg13g2_buf_1 fanout459 (.A(net470),
    .X(net459));
 sg13g2_nand2_1 _07650_ (.Y(_02384_),
    .A(net146),
    .B(_02195_));
 sg13g2_nor2_1 _07651_ (.A(net152),
    .B(net64),
    .Y(_02385_));
 sg13g2_a21oi_1 _07652_ (.A1(net84),
    .A2(_02385_),
    .Y(_02386_),
    .B1(_02107_));
 sg13g2_nor2_1 _07653_ (.A(net84),
    .B(_02385_),
    .Y(_02387_));
 sg13g2_nand2_1 _07654_ (.Y(_02388_),
    .A(_01759_),
    .B(net83));
 sg13g2_o21ai_1 _07655_ (.B1(_02388_),
    .Y(_02389_),
    .A1(_02386_),
    .A2(_02387_));
 sg13g2_nand2_1 _07656_ (.Y(_02390_),
    .A(net160),
    .B(_01831_));
 sg13g2_inv_1 _07657_ (.Y(_02391_),
    .A(net163));
 sg13g2_a21oi_1 _07658_ (.A1(_02391_),
    .A2(net95),
    .Y(_02392_),
    .B1(_01709_));
 sg13g2_nor2_1 _07659_ (.A(net162),
    .B(net164),
    .Y(_02393_));
 sg13g2_a21oi_1 _07660_ (.A1(net95),
    .A2(_02393_),
    .Y(_02394_),
    .B1(\median_processor.input_storage[57] ));
 sg13g2_nand2b_1 _07661_ (.Y(_02395_),
    .B(net93),
    .A_N(net160));
 sg13g2_o21ai_1 _07662_ (.B1(_02395_),
    .Y(_02396_),
    .A1(_02392_),
    .A2(_02394_));
 sg13g2_a22oi_1 _07663_ (.Y(_02397_),
    .B1(_02390_),
    .B2(_02396_),
    .A2(net90),
    .A1(_01719_));
 sg13g2_a21oi_1 _07664_ (.A1(net157),
    .A2(_01835_),
    .Y(_02398_),
    .B1(_02397_));
 sg13g2_a22oi_1 _07665_ (.Y(_02399_),
    .B1(net65),
    .B2(net152),
    .A2(net66),
    .A1(net148));
 sg13g2_nand2_1 _07666_ (.Y(_02400_),
    .A(_02384_),
    .B(_02399_));
 sg13g2_a21oi_1 _07667_ (.A1(net156),
    .A2(_02214_),
    .Y(_02401_),
    .B1(_02400_));
 sg13g2_nor3_1 _07668_ (.A(net156),
    .B(_02214_),
    .C(_02400_),
    .Y(_02402_));
 sg13g2_a221oi_1 _07669_ (.B2(_02401_),
    .C1(_02402_),
    .B1(_02398_),
    .A1(_02384_),
    .Y(_02403_),
    .A2(_02389_));
 sg13g2_buf_1 fanout458 (.A(net459),
    .X(net458));
 sg13g2_buf_2 fanout457 (.A(net458),
    .X(net457));
 sg13g2_xnor2_1 _07672_ (.Y(_02406_),
    .A(net17),
    .B(_02403_));
 sg13g2_nor3_1 _07673_ (.A(_02362_),
    .B(_02363_),
    .C(_02406_),
    .Y(_02407_));
 sg13g2_and2_1 _07674_ (.A(net17),
    .B(net18),
    .X(_02408_));
 sg13g2_nor2_1 _07675_ (.A(net17),
    .B(_02403_),
    .Y(_02409_));
 sg13g2_a22oi_1 _07676_ (.Y(_02410_),
    .B1(_02409_),
    .B2(_02363_),
    .A2(_02408_),
    .A1(_02362_));
 sg13g2_nand2b_1 _07677_ (.Y(_02411_),
    .B(_02410_),
    .A_N(_02407_));
 sg13g2_or2_1 _07678_ (.X(_02412_),
    .B(_02403_),
    .A(net17));
 sg13g2_mux2_1 _07679_ (.A0(_02406_),
    .A1(_02412_),
    .S(_02360_),
    .X(_02413_));
 sg13g2_nand3b_1 _07680_ (.B(_02409_),
    .C(_02334_),
    .Y(_02414_),
    .A_N(_02360_));
 sg13g2_o21ai_1 _07681_ (.B1(_02414_),
    .Y(_02415_),
    .A1(_02334_),
    .A2(_02413_));
 sg13g2_nor2_1 _07682_ (.A(_02311_),
    .B(_02331_),
    .Y(_02416_));
 sg13g2_nor2_1 _07683_ (.A(_02332_),
    .B(_02416_),
    .Y(_02417_));
 sg13g2_nand3_1 _07684_ (.B(_02416_),
    .C(_02409_),
    .A(_02362_),
    .Y(_02418_));
 sg13g2_nand2_1 _07685_ (.Y(_02419_),
    .A(_02068_),
    .B(_02418_));
 sg13g2_a221oi_1 _07686_ (.B2(_02417_),
    .C1(_02419_),
    .B1(_02415_),
    .A1(_02332_),
    .Y(_02420_),
    .A2(_02411_));
 sg13g2_nor2_1 _07687_ (.A(_02362_),
    .B(_02363_),
    .Y(_02421_));
 sg13g2_and2_1 _07688_ (.A(_02332_),
    .B(_02408_),
    .X(_02422_));
 sg13g2_a21o_1 _07689_ (.A2(_02409_),
    .A1(_02416_),
    .B1(_02422_),
    .X(_02423_));
 sg13g2_a22oi_1 _07690_ (.Y(_02424_),
    .B1(_02416_),
    .B2(_02362_),
    .A2(_02363_),
    .A1(_02332_));
 sg13g2_o21ai_1 _07691_ (.B1(_01974_),
    .Y(_02425_),
    .A1(_02406_),
    .A2(_02424_));
 sg13g2_a221oi_1 _07692_ (.B2(_02417_),
    .C1(_02425_),
    .B1(_02411_),
    .A1(_02421_),
    .Y(_02426_),
    .A2(_02423_));
 sg13g2_nor2_2 _07693_ (.A(_02420_),
    .B(_02426_),
    .Y(_02427_));
 sg13g2_buf_1 fanout456 (.A(net458),
    .X(net456));
 sg13g2_nand2_1 _07695_ (.Y(_02429_),
    .A(net149),
    .B(net59));
 sg13g2_o21ai_1 _07696_ (.B1(_02429_),
    .Y(_02430_),
    .A1(_01759_),
    .A2(net180));
 sg13g2_nor2b_1 _07697_ (.A(net190),
    .B_N(net156),
    .Y(_02431_));
 sg13g2_a21oi_1 _07698_ (.A1(net154),
    .A2(_02431_),
    .Y(_02432_),
    .B1(_01998_));
 sg13g2_nor2_1 _07699_ (.A(net154),
    .B(_02431_),
    .Y(_02433_));
 sg13g2_nor2_1 _07700_ (.A(_02432_),
    .B(_02433_),
    .Y(_02434_));
 sg13g2_nand2b_1 _07701_ (.Y(_02435_),
    .B(net183),
    .A_N(net149));
 sg13g2_a21oi_1 _07702_ (.A1(net146),
    .A2(net55),
    .Y(_02436_),
    .B1(_02435_));
 sg13g2_a21oi_1 _07703_ (.A1(_01759_),
    .A2(net180),
    .Y(_02437_),
    .B1(_02436_));
 sg13g2_o21ai_1 _07704_ (.B1(_02437_),
    .Y(_02438_),
    .A1(_02430_),
    .A2(_02434_));
 sg13g2_buf_2 fanout455 (.A(net459),
    .X(net455));
 sg13g2_xnor2_1 _07706_ (.Y(_02440_),
    .A(net156),
    .B(net190));
 sg13g2_xor2_1 _07707_ (.B(net188),
    .A(net154),
    .X(_02441_));
 sg13g2_xor2_1 _07708_ (.B(net180),
    .A(net146),
    .X(_02442_));
 sg13g2_nor2_1 _07709_ (.A(_02441_),
    .B(_02442_),
    .Y(_02443_));
 sg13g2_and4_1 _07710_ (.A(_02429_),
    .B(_02435_),
    .C(_02440_),
    .D(_02443_),
    .X(_02444_));
 sg13g2_xnor2_1 _07711_ (.Y(_02445_),
    .A(net163),
    .B(net75));
 sg13g2_nand2b_1 _07712_ (.Y(_02446_),
    .B(net194),
    .A_N(net160));
 sg13g2_nand2_1 _07713_ (.Y(_02447_),
    .A(net160),
    .B(net60));
 sg13g2_xor2_1 _07714_ (.B(net74),
    .A(net161),
    .X(_02448_));
 sg13g2_xor2_1 _07715_ (.B(net191),
    .A(net158),
    .X(_02449_));
 sg13g2_nor2_1 _07716_ (.A(_02448_),
    .B(_02449_),
    .Y(_02450_));
 sg13g2_nand4_1 _07717_ (.B(_02446_),
    .C(_02447_),
    .A(_02445_),
    .Y(_02451_),
    .D(_02450_));
 sg13g2_nand2b_1 _07718_ (.Y(_02452_),
    .B(net75),
    .A_N(net163));
 sg13g2_nand3_1 _07719_ (.B(_02452_),
    .C(_02446_),
    .A(_01985_),
    .Y(_02453_));
 sg13g2_nand3b_1 _07720_ (.B(net74),
    .C(net75),
    .Y(_02454_),
    .A_N(net163));
 sg13g2_nand3_1 _07721_ (.B(_02446_),
    .C(_02454_),
    .A(net161),
    .Y(_02455_));
 sg13g2_nand4_1 _07722_ (.B(_02447_),
    .C(_02453_),
    .A(net191),
    .Y(_02456_),
    .D(_02455_));
 sg13g2_nand2_1 _07723_ (.Y(_02457_),
    .A(net161),
    .B(_02454_));
 sg13g2_a221oi_1 _07724_ (.B2(_02452_),
    .C1(net158),
    .B1(_01985_),
    .A1(net160),
    .Y(_02458_),
    .A2(net60));
 sg13g2_a21oi_1 _07725_ (.A1(_02284_),
    .A2(_02446_),
    .Y(_02459_),
    .B1(net158));
 sg13g2_a21oi_1 _07726_ (.A1(_02457_),
    .A2(_02458_),
    .Y(_02460_),
    .B1(_02459_));
 sg13g2_nand4_1 _07727_ (.B(_02451_),
    .C(_02456_),
    .A(_02444_),
    .Y(_02461_),
    .D(_02460_));
 sg13g2_buf_1 fanout454 (.A(net470),
    .X(net454));
 sg13g2_nand2_2 _07729_ (.Y(_02463_),
    .A(_02438_),
    .B(_02461_));
 sg13g2_buf_1 fanout453 (.A(net454),
    .X(net453));
 sg13g2_nand2b_1 _07731_ (.Y(_02465_),
    .B(net89),
    .A_N(net154));
 sg13g2_nand2_1 _07732_ (.Y(_02466_),
    .A(net149),
    .B(_02465_));
 sg13g2_o21ai_1 _07733_ (.B1(net56),
    .Y(_02467_),
    .A1(net149),
    .A2(_02465_));
 sg13g2_a22oi_1 _07734_ (.Y(_02468_),
    .B1(_02466_),
    .B2(_02467_),
    .A2(net77),
    .A1(_01759_));
 sg13g2_a21oi_1 _07735_ (.A1(net146),
    .A2(net57),
    .Y(_02469_),
    .B1(_02468_));
 sg13g2_nor2_1 _07736_ (.A(net77),
    .B(net80),
    .Y(_02470_));
 sg13g2_a21oi_1 _07737_ (.A1(net149),
    .A2(_02470_),
    .Y(_02471_),
    .B1(net146));
 sg13g2_a21oi_1 _07738_ (.A1(net56),
    .A2(net149),
    .Y(_02472_),
    .B1(net57));
 sg13g2_nand2_1 _07739_ (.Y(_02473_),
    .A(_02053_),
    .B(net152));
 sg13g2_o21ai_1 _07740_ (.B1(_02473_),
    .Y(_02474_),
    .A1(_02471_),
    .A2(_02472_));
 sg13g2_nor2_1 _07741_ (.A(net196),
    .B(_02391_),
    .Y(_02475_));
 sg13g2_nand2_1 _07742_ (.Y(_02476_),
    .A(net162),
    .B(_02475_));
 sg13g2_o21ai_1 _07743_ (.B1(_02174_),
    .Y(_02477_),
    .A1(net162),
    .A2(_02475_));
 sg13g2_nor2_1 _07744_ (.A(_02176_),
    .B(net160),
    .Y(_02478_));
 sg13g2_a221oi_1 _07745_ (.B2(_02477_),
    .C1(_02478_),
    .B1(_02476_),
    .A1(net128),
    .Y(_02479_),
    .A2(_01719_));
 sg13g2_nor2b_1 _07746_ (.A(net150),
    .B_N(net160),
    .Y(_02480_));
 sg13g2_o21ai_1 _07747_ (.B1(_02480_),
    .Y(_02481_),
    .A1(_02040_),
    .A2(net158));
 sg13g2_o21ai_1 _07748_ (.B1(_02481_),
    .Y(_02482_),
    .A1(net128),
    .A2(_01719_));
 sg13g2_nor4_1 _07749_ (.A(_02042_),
    .B(_02474_),
    .C(_02479_),
    .D(_02482_),
    .Y(_02483_));
 sg13g2_nor4_1 _07750_ (.A(net156),
    .B(_02474_),
    .C(_02479_),
    .D(_02482_),
    .Y(_02484_));
 sg13g2_nor3_1 _07751_ (.A(net156),
    .B(net58),
    .C(_02474_),
    .Y(_02485_));
 sg13g2_nor4_2 _07752_ (.A(_02469_),
    .B(_02483_),
    .C(_02484_),
    .Y(_02486_),
    .D(_02485_));
 sg13g2_buf_1 fanout452 (.A(net453),
    .X(net452));
 sg13g2_and2_1 _07754_ (.A(_02463_),
    .B(_02486_),
    .X(_02488_));
 sg13g2_nor2_1 _07755_ (.A(_02463_),
    .B(_02486_),
    .Y(_02489_));
 sg13g2_nand2_1 _07756_ (.Y(_02490_),
    .A(net155),
    .B(_01877_));
 sg13g2_nand2_1 _07757_ (.Y(_02491_),
    .A(\median_processor.input_storage[21] ),
    .B(_02490_));
 sg13g2_nand2_1 _07758_ (.Y(_02492_),
    .A(net147),
    .B(net54));
 sg13g2_nand2_1 _07759_ (.Y(_02493_),
    .A(_02107_),
    .B(_02492_));
 sg13g2_nand2_1 _07760_ (.Y(_02494_),
    .A(\median_processor.input_storage[22] ),
    .B(_02492_));
 sg13g2_nor2_1 _07761_ (.A(\median_processor.input_storage[21] ),
    .B(_02490_),
    .Y(_02495_));
 sg13g2_a221oi_1 _07762_ (.B2(_02494_),
    .C1(_02495_),
    .B1(_02493_),
    .A1(net153),
    .Y(_02496_),
    .A2(_02491_));
 sg13g2_nand3_1 _07763_ (.B(\median_processor.input_storage[22] ),
    .C(_02492_),
    .A(_02107_),
    .Y(_02497_));
 sg13g2_o21ai_1 _07764_ (.B1(_02497_),
    .Y(_02498_),
    .A1(net147),
    .A2(net54));
 sg13g2_and2_1 _07765_ (.A(\median_processor.input_storage[17] ),
    .B(net179),
    .X(_02499_));
 sg13g2_nand2b_1 _07766_ (.Y(_02500_),
    .B(net175),
    .A_N(net159));
 sg13g2_nand2_1 _07767_ (.Y(_02501_),
    .A(_01895_),
    .B(_02500_));
 sg13g2_nand2_1 _07768_ (.Y(_02502_),
    .A(net157),
    .B(_02500_));
 sg13g2_inv_2 _07769_ (.Y(_02503_),
    .A(\median_processor.input_storage[17] ));
 sg13g2_nand2b_1 _07770_ (.Y(_02504_),
    .B(net178),
    .A_N(net163));
 sg13g2_a21oi_1 _07771_ (.A1(_02503_),
    .A2(_02504_),
    .Y(_02505_),
    .B1(net161));
 sg13g2_a221oi_1 _07772_ (.B2(_02502_),
    .C1(_02505_),
    .B1(_02501_),
    .A1(_02391_),
    .Y(_02506_),
    .A2(_02499_));
 sg13g2_nor2b_1 _07773_ (.A(net175),
    .B_N(net159),
    .Y(_02507_));
 sg13g2_o21ai_1 _07774_ (.B1(_02507_),
    .Y(_02508_),
    .A1(\median_processor.input_storage[27] ),
    .A2(_01895_));
 sg13g2_o21ai_1 _07775_ (.B1(_02508_),
    .Y(_02509_),
    .A1(_01719_),
    .A2(net173));
 sg13g2_xnor2_1 _07776_ (.Y(_02510_),
    .A(net155),
    .B(net171));
 sg13g2_xnor2_1 _07777_ (.Y(_02511_),
    .A(net147),
    .B(net165));
 sg13g2_xnor2_1 _07778_ (.Y(_02512_),
    .A(net153),
    .B(net169));
 sg13g2_xnor2_1 _07779_ (.Y(_02513_),
    .A(\median_processor.input_storage[30] ),
    .B(net167));
 sg13g2_nand4_1 _07780_ (.B(_02511_),
    .C(_02512_),
    .A(_02510_),
    .Y(_02514_),
    .D(_02513_));
 sg13g2_xor2_1 _07781_ (.B(net178),
    .A(net163),
    .X(_02515_));
 sg13g2_xor2_1 _07782_ (.B(net175),
    .A(net159),
    .X(_02516_));
 sg13g2_xor2_1 _07783_ (.B(net173),
    .A(net157),
    .X(_02517_));
 sg13g2_xor2_1 _07784_ (.B(net177),
    .A(net161),
    .X(_02518_));
 sg13g2_nor4_1 _07785_ (.A(_02515_),
    .B(_02516_),
    .C(_02517_),
    .D(_02518_),
    .Y(_02519_));
 sg13g2_nor2_1 _07786_ (.A(_02514_),
    .B(_02519_),
    .Y(_02520_));
 sg13g2_o21ai_1 _07787_ (.B1(_02520_),
    .Y(_02521_),
    .A1(_02506_),
    .A2(_02509_));
 sg13g2_o21ai_1 _07788_ (.B1(_02521_),
    .Y(_02522_),
    .A1(_02496_),
    .A2(_02498_));
 sg13g2_buf_2 fanout451 (.A(net453),
    .X(net451));
 sg13g2_buf_2 fanout450 (.A(net454),
    .X(net450));
 sg13g2_nand2_1 _07791_ (.Y(_02525_),
    .A(_02107_),
    .B(net132));
 sg13g2_o21ai_1 _07792_ (.B1(net147),
    .Y(_02526_),
    .A1(net63),
    .A2(_02525_));
 sg13g2_nand2_1 _07793_ (.Y(_02527_),
    .A(net63),
    .B(_02525_));
 sg13g2_nand2b_1 _07794_ (.Y(_02528_),
    .B(\median_processor.input_storage[26] ),
    .A_N(net140));
 sg13g2_nor2_1 _07795_ (.A(net138),
    .B(_02528_),
    .Y(_02529_));
 sg13g2_a21oi_1 _07796_ (.A1(\median_processor.input_storage[28] ),
    .A2(_01941_),
    .Y(_02530_),
    .B1(_02529_));
 sg13g2_nor2b_1 _07797_ (.A(net164),
    .B_N(net144),
    .Y(_02531_));
 sg13g2_nor2b_1 _07798_ (.A(net159),
    .B_N(net140),
    .Y(_02532_));
 sg13g2_a221oi_1 _07799_ (.B2(_02531_),
    .C1(_02532_),
    .B1(net143),
    .A1(_01719_),
    .Y(_02533_),
    .A2(net138));
 sg13g2_o21ai_1 _07800_ (.B1(_01709_),
    .Y(_02534_),
    .A1(net143),
    .A2(_02531_));
 sg13g2_nand2_1 _07801_ (.Y(_02535_),
    .A(net138),
    .B(_02528_));
 sg13g2_nand2b_1 _07802_ (.Y(_02536_),
    .B(net148),
    .A_N(net133));
 sg13g2_nand2b_1 _07803_ (.Y(_02537_),
    .B(net146),
    .A_N(net131));
 sg13g2_nand2b_1 _07804_ (.Y(_02538_),
    .B(net152),
    .A_N(net135));
 sg13g2_nand3_1 _07805_ (.B(_02537_),
    .C(_02538_),
    .A(_02536_),
    .Y(_02539_));
 sg13g2_a221oi_1 _07806_ (.B2(net157),
    .C1(_02539_),
    .B1(_02535_),
    .A1(_02533_),
    .Y(_02540_),
    .A2(_02534_));
 sg13g2_nand2b_1 _07807_ (.Y(_02541_),
    .B(net137),
    .A_N(net155));
 sg13g2_o21ai_1 _07808_ (.B1(_02541_),
    .Y(_02542_),
    .A1(net152),
    .A2(_02154_));
 sg13g2_nor2b_1 _07809_ (.A(_02539_),
    .B_N(_02542_),
    .Y(_02543_));
 sg13g2_a221oi_1 _07810_ (.B2(_02540_),
    .C1(_02543_),
    .B1(_02530_),
    .A1(_02526_),
    .Y(_02544_),
    .A2(_02527_));
 sg13g2_buf_2 fanout449 (.A(net454),
    .X(net449));
 sg13g2_nand2_1 _07812_ (.Y(_02546_),
    .A(net23),
    .B(net35));
 sg13g2_o21ai_1 _07813_ (.B1(net32),
    .Y(_02547_),
    .A1(net23),
    .A2(net35));
 sg13g2_nand2_1 _07814_ (.Y(_02548_),
    .A(_02546_),
    .B(_02547_));
 sg13g2_mux2_1 _07815_ (.A0(_02488_),
    .A1(_02489_),
    .S(_02548_),
    .X(_02549_));
 sg13g2_xor2_1 _07816_ (.B(net35),
    .A(net23),
    .X(_02550_));
 sg13g2_xnor2_1 _07817_ (.Y(_02551_),
    .A(net32),
    .B(_02550_));
 sg13g2_xnor2_1 _07818_ (.Y(_02552_),
    .A(_02261_),
    .B(_02551_));
 sg13g2_nor3_1 _07819_ (.A(_02122_),
    .B(net18),
    .C(_02551_),
    .Y(_02553_));
 sg13g2_a21o_1 _07820_ (.A2(_02552_),
    .A1(net18),
    .B1(_02553_),
    .X(_02554_));
 sg13g2_nor4_1 _07821_ (.A(_01859_),
    .B(_02122_),
    .C(net23),
    .D(net35),
    .Y(_02555_));
 sg13g2_nor3_1 _07822_ (.A(net32),
    .B(_02261_),
    .C(_02546_),
    .Y(_02556_));
 sg13g2_o21ai_1 _07823_ (.B1(net18),
    .Y(_02557_),
    .A1(_02555_),
    .A2(_02556_));
 sg13g2_xnor2_1 _07824_ (.Y(_02558_),
    .A(net32),
    .B(_02261_));
 sg13g2_or3_1 _07825_ (.A(net18),
    .B(_02546_),
    .C(_02558_),
    .X(_02559_));
 sg13g2_a221oi_1 _07826_ (.B2(_01759_),
    .C1(_01859_),
    .B1(_02121_),
    .A1(_02109_),
    .Y(_02560_),
    .A2(_02114_));
 sg13g2_o21ai_1 _07827_ (.B1(_02550_),
    .Y(_02561_),
    .A1(net18),
    .A2(_02560_));
 sg13g2_a21o_1 _07828_ (.A2(_02558_),
    .A1(net18),
    .B1(_02561_),
    .X(_02562_));
 sg13g2_nand3_1 _07829_ (.B(_02559_),
    .C(_02562_),
    .A(_02557_),
    .Y(_02563_));
 sg13g2_nor2_1 _07830_ (.A(_02488_),
    .B(_02489_),
    .Y(_02564_));
 sg13g2_nand2_1 _07831_ (.Y(_02565_),
    .A(_02463_),
    .B(_02486_));
 sg13g2_nor2_1 _07832_ (.A(net32),
    .B(_02546_),
    .Y(_02566_));
 sg13g2_a21oi_1 _07833_ (.A1(net32),
    .A2(_02550_),
    .Y(_02567_),
    .B1(_02566_));
 sg13g2_nor4_1 _07834_ (.A(_02261_),
    .B(net18),
    .C(_02565_),
    .D(_02567_),
    .Y(_02568_));
 sg13g2_a221oi_1 _07835_ (.B2(_02564_),
    .C1(_02568_),
    .B1(_02563_),
    .A1(_02549_),
    .Y(_02569_),
    .A2(_02554_));
 sg13g2_buf_1 fanout448 (.A(net454),
    .X(net448));
 sg13g2_xnor2_1 _07837_ (.Y(_02571_),
    .A(_02360_),
    .B(net35));
 sg13g2_nor2_1 _07838_ (.A(_01941_),
    .B(net172),
    .Y(_02572_));
 sg13g2_nor2_1 _07839_ (.A(_02154_),
    .B(net169),
    .Y(_02573_));
 sg13g2_nand2_1 _07840_ (.Y(_02574_),
    .A(net133),
    .B(_02364_));
 sg13g2_a21oi_1 _07841_ (.A1(net133),
    .A2(_01869_),
    .Y(_02575_),
    .B1(net131));
 sg13g2_a21oi_1 _07842_ (.A1(net166),
    .A2(_02574_),
    .Y(_02576_),
    .B1(_02575_));
 sg13g2_nand2_1 _07843_ (.Y(_02577_),
    .A(net177),
    .B(net178));
 sg13g2_o21ai_1 _07844_ (.B1(net143),
    .Y(_02578_),
    .A1(net144),
    .A2(_02577_));
 sg13g2_inv_2 _07845_ (.Y(_02579_),
    .A(net175));
 sg13g2_nand2b_1 _07846_ (.Y(_02580_),
    .B(net178),
    .A_N(net144));
 sg13g2_nor2b_1 _07847_ (.A(net173),
    .B_N(net138),
    .Y(_02581_));
 sg13g2_a221oi_1 _07848_ (.B2(_02580_),
    .C1(_02581_),
    .B1(_02503_),
    .A1(net140),
    .Y(_02582_),
    .A2(_02579_));
 sg13g2_nand2b_1 _07849_ (.Y(_02583_),
    .B(net175),
    .A_N(net140));
 sg13g2_o21ai_1 _07850_ (.B1(_01895_),
    .Y(_02584_),
    .A1(net138),
    .A2(_02583_));
 sg13g2_nand2_1 _07851_ (.Y(_02585_),
    .A(net138),
    .B(_02583_));
 sg13g2_nor2_1 _07852_ (.A(net137),
    .B(_01877_),
    .Y(_02586_));
 sg13g2_a221oi_1 _07853_ (.B2(_02585_),
    .C1(_02586_),
    .B1(_02584_),
    .A1(_02578_),
    .Y(_02587_),
    .A2(_02582_));
 sg13g2_nor4_2 _07854_ (.A(_02572_),
    .B(_02573_),
    .C(_02576_),
    .Y(_02588_),
    .D(_02587_));
 sg13g2_xor2_1 _07855_ (.B(net167),
    .A(net132),
    .X(_02589_));
 sg13g2_xor2_1 _07856_ (.B(net165),
    .A(net131),
    .X(_02590_));
 sg13g2_nor2_1 _07857_ (.A(net135),
    .B(_01873_),
    .Y(_02591_));
 sg13g2_nor3_1 _07858_ (.A(_02589_),
    .B(_02590_),
    .C(_02591_),
    .Y(_02592_));
 sg13g2_xor2_1 _07859_ (.B(net176),
    .A(net140),
    .X(_02593_));
 sg13g2_xor2_1 _07860_ (.B(net177),
    .A(net143),
    .X(_02594_));
 sg13g2_nor4_1 _07861_ (.A(_02589_),
    .B(_02590_),
    .C(_02593_),
    .D(_02594_),
    .Y(_02595_));
 sg13g2_xor2_1 _07862_ (.B(net173),
    .A(net138),
    .X(_02596_));
 sg13g2_xor2_1 _07863_ (.B(net171),
    .A(net137),
    .X(_02597_));
 sg13g2_xor2_1 _07864_ (.B(net169),
    .A(net134),
    .X(_02598_));
 sg13g2_xor2_1 _07865_ (.B(net178),
    .A(net144),
    .X(_02599_));
 sg13g2_nor4_1 _07866_ (.A(_02596_),
    .B(_02597_),
    .C(_02598_),
    .D(_02599_),
    .Y(_02600_));
 sg13g2_nand2_1 _07867_ (.Y(_02601_),
    .A(_02595_),
    .B(_02600_));
 sg13g2_o21ai_1 _07868_ (.B1(_02601_),
    .Y(_02602_),
    .A1(_02576_),
    .A2(_02592_));
 sg13g2_buf_2 fanout447 (.A(net448),
    .X(net447));
 sg13g2_nor2_2 _07870_ (.A(_02588_),
    .B(_02602_),
    .Y(_02604_));
 sg13g2_buf_2 fanout446 (.A(net448),
    .X(net446));
 sg13g2_nand3_1 _07872_ (.B(_02571_),
    .C(_02604_),
    .A(net27),
    .Y(_02606_));
 sg13g2_and2_1 _07873_ (.A(_01922_),
    .B(_02353_),
    .X(_02607_));
 sg13g2_nor3_1 _07874_ (.A(_02359_),
    .B(_02607_),
    .C(_02544_),
    .Y(_02608_));
 sg13g2_or2_1 _07875_ (.X(_02609_),
    .B(_02602_),
    .A(_02588_));
 sg13g2_buf_1 fanout445 (.A(net470),
    .X(net445));
 sg13g2_xnor2_1 _07877_ (.Y(_02611_),
    .A(net27),
    .B(_02609_));
 sg13g2_nand2_1 _07878_ (.Y(_02612_),
    .A(_02608_),
    .B(_02611_));
 sg13g2_nand2_1 _07879_ (.Y(_02613_),
    .A(_02176_),
    .B(net141));
 sg13g2_o21ai_1 _07880_ (.B1(_02613_),
    .Y(_02614_),
    .A1(net128),
    .A2(net62));
 sg13g2_nor2b_1 _07881_ (.A(net196),
    .B_N(net145),
    .Y(_02615_));
 sg13g2_nand2_1 _07882_ (.Y(_02616_),
    .A(net142),
    .B(_02615_));
 sg13g2_o21ai_1 _07883_ (.B1(_02174_),
    .Y(_02617_),
    .A1(net142),
    .A2(_02615_));
 sg13g2_a22oi_1 _07884_ (.Y(_02618_),
    .B1(_02616_),
    .B2(_02617_),
    .A2(_01918_),
    .A1(net150));
 sg13g2_nor2_1 _07885_ (.A(net58),
    .B(net136),
    .Y(_02619_));
 sg13g2_a221oi_1 _07886_ (.B2(net129),
    .C1(_02619_),
    .B1(net62),
    .A1(net89),
    .Y(_02620_),
    .A2(_02154_));
 sg13g2_o21ai_1 _07887_ (.B1(_02620_),
    .Y(_02621_),
    .A1(_02614_),
    .A2(_02618_));
 sg13g2_nand3_1 _07888_ (.B(net134),
    .C(net136),
    .A(net58),
    .Y(_02622_));
 sg13g2_a21oi_1 _07889_ (.A1(net58),
    .A2(net136),
    .Y(_02623_),
    .B1(net134));
 sg13g2_a21oi_1 _07890_ (.A1(net89),
    .A2(_02622_),
    .Y(_02624_),
    .B1(_02623_));
 sg13g2_a221oi_1 _07891_ (.B2(net56),
    .C1(_02624_),
    .B1(net132),
    .A1(net57),
    .Y(_02625_),
    .A2(net130));
 sg13g2_nand2_1 _07892_ (.Y(_02626_),
    .A(net80),
    .B(net61));
 sg13g2_nand2_1 _07893_ (.Y(_02627_),
    .A(net130),
    .B(_02626_));
 sg13g2_o21ai_1 _07894_ (.B1(net57),
    .Y(_02628_),
    .A1(net130),
    .A2(_02626_));
 sg13g2_a22oi_1 _07895_ (.Y(_02629_),
    .B1(_02627_),
    .B2(_02628_),
    .A2(_02625_),
    .A1(_02621_));
 sg13g2_buf_2 fanout444 (.A(net445),
    .X(net444));
 sg13g2_xor2_1 _07897_ (.B(_02629_),
    .A(_02170_),
    .X(_02631_));
 sg13g2_nand2b_1 _07898_ (.Y(_02632_),
    .B(net136),
    .A_N(net190));
 sg13g2_nand2_1 _07899_ (.Y(_02633_),
    .A(net186),
    .B(_02632_));
 sg13g2_nand2b_1 _07900_ (.Y(_02634_),
    .B(net130),
    .A_N(net180));
 sg13g2_nand2_1 _07901_ (.Y(_02635_),
    .A(net61),
    .B(_02634_));
 sg13g2_nand2_1 _07902_ (.Y(_02636_),
    .A(net183),
    .B(_02634_));
 sg13g2_nor2_1 _07903_ (.A(net186),
    .B(_02632_),
    .Y(_02637_));
 sg13g2_a221oi_1 _07904_ (.B2(_02636_),
    .C1(_02637_),
    .B1(_02635_),
    .A1(net134),
    .Y(_02638_),
    .A2(_02633_));
 sg13g2_nand3_1 _07905_ (.B(net183),
    .C(_02634_),
    .A(net61),
    .Y(_02639_));
 sg13g2_o21ai_1 _07906_ (.B1(_02639_),
    .Y(_02640_),
    .A1(net130),
    .A2(net55));
 sg13g2_or2_1 _07907_ (.X(_02641_),
    .B(_02640_),
    .A(_02638_));
 sg13g2_buf_2 fanout443 (.A(net444),
    .X(net443));
 sg13g2_nand2_1 _07909_ (.Y(_02643_),
    .A(net62),
    .B(net191));
 sg13g2_nand2b_1 _07910_ (.Y(_02644_),
    .B(net76),
    .A_N(net145));
 sg13g2_a21oi_1 _07911_ (.A1(net142),
    .A2(_02644_),
    .Y(_02645_),
    .B1(_01985_));
 sg13g2_nor2_1 _07912_ (.A(net142),
    .B(_02644_),
    .Y(_02646_));
 sg13g2_a22oi_1 _07913_ (.Y(_02647_),
    .B1(net60),
    .B2(net141),
    .A2(_02284_),
    .A1(net139));
 sg13g2_o21ai_1 _07914_ (.B1(_02647_),
    .Y(_02648_),
    .A1(_02645_),
    .A2(_02646_));
 sg13g2_nor2_1 _07915_ (.A(net141),
    .B(net60),
    .Y(_02649_));
 sg13g2_o21ai_1 _07916_ (.B1(_02649_),
    .Y(_02650_),
    .A1(net62),
    .A2(net191));
 sg13g2_xnor2_1 _07917_ (.Y(_02651_),
    .A(net130),
    .B(net180));
 sg13g2_xnor2_1 _07918_ (.Y(_02652_),
    .A(net136),
    .B(net189));
 sg13g2_xnor2_1 _07919_ (.Y(_02653_),
    .A(net134),
    .B(net187));
 sg13g2_xnor2_1 _07920_ (.Y(_02654_),
    .A(net132),
    .B(net183));
 sg13g2_nand4_1 _07921_ (.B(_02652_),
    .C(_02653_),
    .A(_02651_),
    .Y(_02655_),
    .D(_02654_));
 sg13g2_xor2_1 _07922_ (.B(net74),
    .A(net142),
    .X(_02656_));
 sg13g2_xor2_1 _07923_ (.B(net195),
    .A(net141),
    .X(_02657_));
 sg13g2_xor2_1 _07924_ (.B(net192),
    .A(net139),
    .X(_02658_));
 sg13g2_xor2_1 _07925_ (.B(net75),
    .A(net145),
    .X(_02659_));
 sg13g2_nor4_1 _07926_ (.A(_02656_),
    .B(_02657_),
    .C(_02658_),
    .D(_02659_),
    .Y(_02660_));
 sg13g2_nor2_1 _07927_ (.A(_02655_),
    .B(_02660_),
    .Y(_02661_));
 sg13g2_nand4_1 _07928_ (.B(_02648_),
    .C(_02650_),
    .A(_02643_),
    .Y(_02662_),
    .D(_02661_));
 sg13g2_and2_1 _07929_ (.A(_02641_),
    .B(_02662_),
    .X(_02663_));
 sg13g2_buf_1 fanout442 (.A(net445),
    .X(net442));
 sg13g2_nand2b_1 _07931_ (.Y(_02665_),
    .B(net22),
    .A_N(_02631_));
 sg13g2_a21oi_1 _07932_ (.A1(_02606_),
    .A2(_02612_),
    .Y(_02666_),
    .B1(_02665_));
 sg13g2_nand2b_1 _07933_ (.Y(_02667_),
    .B(_02629_),
    .A_N(_02170_));
 sg13g2_nand3_1 _07934_ (.B(net35),
    .C(_02604_),
    .A(net27),
    .Y(_02668_));
 sg13g2_or3_1 _07935_ (.A(net27),
    .B(net35),
    .C(_02604_),
    .X(_02669_));
 sg13g2_mux2_1 _07936_ (.A0(_02668_),
    .A1(_02669_),
    .S(_02360_),
    .X(_02670_));
 sg13g2_nand2_1 _07937_ (.Y(_02671_),
    .A(_02571_),
    .B(_02611_));
 sg13g2_nor2b_1 _07938_ (.A(_02663_),
    .B_N(_02631_),
    .Y(_02672_));
 sg13g2_a221oi_1 _07939_ (.B2(_02671_),
    .C1(_02672_),
    .B1(_02670_),
    .A1(net22),
    .Y(_02673_),
    .A2(_02667_));
 sg13g2_nand2b_1 _07940_ (.Y(_02674_),
    .B(_02170_),
    .A_N(_02629_));
 sg13g2_o21ai_1 _07941_ (.B1(_02544_),
    .Y(_02675_),
    .A1(_02588_),
    .A2(_02602_));
 sg13g2_nor3_1 _07942_ (.A(net35),
    .B(_02588_),
    .C(_02602_),
    .Y(_02676_));
 sg13g2_a21oi_1 _07943_ (.A1(net27),
    .A2(_02675_),
    .Y(_02677_),
    .B1(_02676_));
 sg13g2_mux2_1 _07944_ (.A0(_02674_),
    .A1(_02667_),
    .S(_02677_),
    .X(_02678_));
 sg13g2_xnor2_1 _07945_ (.Y(_02679_),
    .A(_02571_),
    .B(_02611_));
 sg13g2_nor3_1 _07946_ (.A(net22),
    .B(_02678_),
    .C(_02679_),
    .Y(_02680_));
 sg13g2_nor2b_1 _07947_ (.A(_02674_),
    .B_N(_02676_),
    .Y(_02681_));
 sg13g2_and4_1 _07948_ (.A(net27),
    .B(_02360_),
    .C(net22),
    .D(_02681_),
    .X(_02682_));
 sg13g2_nor3_2 _07949_ (.A(_02673_),
    .B(_02680_),
    .C(_02682_),
    .Y(_02683_));
 sg13g2_nor2b_1 _07950_ (.A(_02666_),
    .B_N(_02683_),
    .Y(_02684_));
 sg13g2_buf_1 fanout441 (.A(net442),
    .X(net441));
 sg13g2_nor2b_1 _07952_ (.A(net190),
    .B_N(net171),
    .Y(_02686_));
 sg13g2_o21ai_1 _07953_ (.B1(_01998_),
    .Y(_02687_),
    .A1(net170),
    .A2(_02686_));
 sg13g2_nand2_1 _07954_ (.Y(_02688_),
    .A(net170),
    .B(_02686_));
 sg13g2_a22oi_1 _07955_ (.Y(_02689_),
    .B1(_02687_),
    .B2(_02688_),
    .A2(_02364_),
    .A1(net184));
 sg13g2_inv_1 _07956_ (.Y(_02690_),
    .A(net76));
 sg13g2_nor2b_1 _07957_ (.A(net192),
    .B_N(net174),
    .Y(_02691_));
 sg13g2_a221oi_1 _07958_ (.B2(_02690_),
    .C1(_02691_),
    .B1(_02499_),
    .A1(net60),
    .Y(_02692_),
    .A2(net176));
 sg13g2_nor2b_1 _07959_ (.A(net76),
    .B_N(net179),
    .Y(_02693_));
 sg13g2_o21ai_1 _07960_ (.B1(_01985_),
    .Y(_02694_),
    .A1(net177),
    .A2(_02693_));
 sg13g2_nor2_1 _07961_ (.A(_01982_),
    .B(net176),
    .Y(_02695_));
 sg13g2_nand2_1 _07962_ (.Y(_02696_),
    .A(_02284_),
    .B(net174));
 sg13g2_nand2b_1 _07963_ (.Y(_02697_),
    .B(net183),
    .A_N(net168));
 sg13g2_nand2b_1 _07964_ (.Y(_02698_),
    .B(net187),
    .A_N(net170));
 sg13g2_nand2b_1 _07965_ (.Y(_02699_),
    .B(net192),
    .A_N(net174));
 sg13g2_nand2b_1 _07966_ (.Y(_02700_),
    .B(net189),
    .A_N(net171));
 sg13g2_nand4_1 _07967_ (.B(_02698_),
    .C(_02699_),
    .A(_02697_),
    .Y(_02701_),
    .D(_02700_));
 sg13g2_a221oi_1 _07968_ (.B2(_02696_),
    .C1(_02701_),
    .B1(_02695_),
    .A1(_02692_),
    .Y(_02702_),
    .A2(_02694_));
 sg13g2_nand2_1 _07969_ (.Y(_02703_),
    .A(_02006_),
    .B(net168));
 sg13g2_o21ai_1 _07970_ (.B1(_02703_),
    .Y(_02704_),
    .A1(net182),
    .A2(net53));
 sg13g2_or3_2 _07971_ (.A(_02689_),
    .B(_02702_),
    .C(_02704_),
    .X(_02705_));
 sg13g2_buf_2 fanout440 (.A(net442),
    .X(net440));
 sg13g2_nor2_1 _07973_ (.A(net78),
    .B(net53),
    .Y(_02707_));
 sg13g2_nand2_1 _07974_ (.Y(_02708_),
    .A(net182),
    .B(net53));
 sg13g2_o21ai_1 _07975_ (.B1(_02708_),
    .Y(_02709_),
    .A1(_02705_),
    .A2(_02707_));
 sg13g2_and2_1 _07976_ (.A(net80),
    .B(_02709_),
    .X(_02710_));
 sg13g2_nand2b_1 _07977_ (.Y(_02711_),
    .B(net179),
    .A_N(net197));
 sg13g2_nand3b_1 _07978_ (.B(net177),
    .C(net179),
    .Y(_02712_),
    .A_N(net197));
 sg13g2_a22oi_1 _07979_ (.Y(_02713_),
    .B1(_02712_),
    .B2(\median_processor.input_storage[1] ),
    .A2(_02711_),
    .A1(_02503_));
 sg13g2_nor2_1 _07980_ (.A(net150),
    .B(_02579_),
    .Y(_02714_));
 sg13g2_nand2_1 _07981_ (.Y(_02715_),
    .A(net150),
    .B(_02579_));
 sg13g2_o21ai_1 _07982_ (.B1(_02715_),
    .Y(_02716_),
    .A1(_02713_),
    .A2(_02714_));
 sg13g2_nand2_1 _07983_ (.Y(_02717_),
    .A(_02040_),
    .B(net174));
 sg13g2_nor2_1 _07984_ (.A(_02040_),
    .B(net174),
    .Y(_02718_));
 sg13g2_a21o_1 _07985_ (.A2(_02717_),
    .A1(_02716_),
    .B1(_02718_),
    .X(_02719_));
 sg13g2_nor2_1 _07986_ (.A(_02053_),
    .B(net170),
    .Y(_02720_));
 sg13g2_nor2_1 _07987_ (.A(net58),
    .B(net171),
    .Y(_02721_));
 sg13g2_or2_1 _07988_ (.X(_02722_),
    .B(_02721_),
    .A(_02720_));
 sg13g2_nand2_1 _07989_ (.Y(_02723_),
    .A(net58),
    .B(net171));
 sg13g2_nand2_1 _07990_ (.Y(_02724_),
    .A(_02053_),
    .B(net170));
 sg13g2_o21ai_1 _07991_ (.B1(_02724_),
    .Y(_02725_),
    .A1(_02723_),
    .A2(_02720_));
 sg13g2_inv_1 _07992_ (.Y(_02726_),
    .A(_02725_));
 sg13g2_o21ai_1 _07993_ (.B1(_02726_),
    .Y(_02727_),
    .A1(_02719_),
    .A2(_02722_));
 sg13g2_buf_1 fanout439 (.A(net470),
    .X(net439));
 sg13g2_nand2_1 _07995_ (.Y(_02729_),
    .A(net168),
    .B(_02727_));
 sg13g2_nor3_2 _07996_ (.A(_02689_),
    .B(_02702_),
    .C(_02704_),
    .Y(_02730_));
 sg13g2_nand2_1 _07997_ (.Y(_02731_),
    .A(_02364_),
    .B(_02730_));
 sg13g2_o21ai_1 _07998_ (.B1(net53),
    .Y(_02732_),
    .A1(net181),
    .A2(_02730_));
 sg13g2_o21ai_1 _07999_ (.B1(_02732_),
    .Y(_02733_),
    .A1(_02727_),
    .A2(_02731_));
 sg13g2_inv_1 _08000_ (.Y(_02734_),
    .A(_01869_));
 sg13g2_o21ai_1 _08001_ (.B1(net57),
    .Y(_02735_),
    .A1(_02734_),
    .A2(_02727_));
 sg13g2_o21ai_1 _08002_ (.B1(net54),
    .Y(_02736_),
    .A1(net78),
    .A2(net181));
 sg13g2_nor2_1 _08003_ (.A(net81),
    .B(net54),
    .Y(_02737_));
 sg13g2_a21oi_1 _08004_ (.A1(net168),
    .A2(_02736_),
    .Y(_02738_),
    .B1(_02737_));
 sg13g2_nor2_1 _08005_ (.A(_02730_),
    .B(_02738_),
    .Y(_02739_));
 sg13g2_nand2b_1 _08006_ (.Y(_02740_),
    .B(net168),
    .A_N(net181));
 sg13g2_o21ai_1 _08007_ (.B1(net54),
    .Y(_02741_),
    .A1(net81),
    .A2(_02740_));
 sg13g2_a22oi_1 _08008_ (.Y(_02742_),
    .B1(_02737_),
    .B2(net168),
    .A2(_02741_),
    .A1(net57));
 sg13g2_and3_1 _08009_ (.X(_02743_),
    .A(_02742_),
    .B(_02724_),
    .C(_02723_));
 sg13g2_nor3_1 _08010_ (.A(net78),
    .B(net182),
    .C(_02720_),
    .Y(_02744_));
 sg13g2_nand2_1 _08011_ (.Y(_02745_),
    .A(_02724_),
    .B(_02721_));
 sg13g2_nand3_1 _08012_ (.B(_02744_),
    .C(_02745_),
    .A(net56),
    .Y(_02746_));
 sg13g2_a221oi_1 _08013_ (.B2(_02742_),
    .C1(_02730_),
    .B1(_02746_),
    .A1(_02743_),
    .Y(_02747_),
    .A2(_02719_));
 sg13g2_a21o_1 _08014_ (.A2(_02739_),
    .A1(_02727_),
    .B1(_02747_),
    .X(_02748_));
 sg13g2_buf_1 fanout438 (.A(net439),
    .X(net438));
 sg13g2_a221oi_1 _08016_ (.B2(_02735_),
    .C1(_02748_),
    .B1(_02733_),
    .A1(_02710_),
    .Y(_02750_),
    .A2(_02729_));
 sg13g2_buf_2 fanout437 (.A(net439),
    .X(net437));
 sg13g2_nor2_2 _08018_ (.A(net17),
    .B(_02750_),
    .Y(_02752_));
 sg13g2_buf_1 fanout436 (.A(net439),
    .X(net436));
 sg13g2_nand2_1 _08020_ (.Y(_02754_),
    .A(net29),
    .B(_02609_));
 sg13g2_and2_1 _08021_ (.A(_02522_),
    .B(_02754_),
    .X(_02755_));
 sg13g2_and2_1 _08022_ (.A(_02748_),
    .B(_02755_),
    .X(_02756_));
 sg13g2_nor2_1 _08023_ (.A(net30),
    .B(_02609_),
    .Y(_02757_));
 sg13g2_nand2_1 _08024_ (.Y(_02758_),
    .A(net23),
    .B(_02757_));
 sg13g2_a21oi_1 _08025_ (.A1(net17),
    .A2(_02750_),
    .Y(_02759_),
    .B1(_02758_));
 sg13g2_a21o_1 _08026_ (.A2(_02752_),
    .A1(_02757_),
    .B1(_02759_),
    .X(_02760_));
 sg13g2_inv_1 _08027_ (.Y(_02761_),
    .A(_02748_));
 sg13g2_nor4_1 _08028_ (.A(net23),
    .B(_02761_),
    .C(_02754_),
    .D(_02752_),
    .Y(_02762_));
 sg13g2_a221oi_1 _08029_ (.B2(_02748_),
    .C1(_02762_),
    .B1(_02760_),
    .A1(_02752_),
    .Y(_02763_),
    .A2(_02756_));
 sg13g2_a21oi_1 _08030_ (.A1(_02757_),
    .A2(_02752_),
    .Y(_02764_),
    .B1(_02759_));
 sg13g2_and2_1 _08031_ (.A(net17),
    .B(_02750_),
    .X(_02765_));
 sg13g2_nand2_1 _08032_ (.Y(_02766_),
    .A(net23),
    .B(_02604_));
 sg13g2_nor2_1 _08033_ (.A(_02522_),
    .B(_02604_),
    .Y(_02767_));
 sg13g2_a21o_1 _08034_ (.A2(_02766_),
    .A1(net30),
    .B1(_02767_),
    .X(_02768_));
 sg13g2_a22oi_1 _08035_ (.Y(_02769_),
    .B1(_02765_),
    .B2(_02768_),
    .A2(_02755_),
    .A1(_02752_));
 sg13g2_nor2_1 _08036_ (.A(net23),
    .B(_02754_),
    .Y(_02770_));
 sg13g2_o21ai_1 _08037_ (.B1(_02770_),
    .Y(_02771_),
    .A1(net17),
    .A2(_02750_));
 sg13g2_nand4_1 _08038_ (.B(_02764_),
    .C(_02769_),
    .A(_02761_),
    .Y(_02772_),
    .D(_02771_));
 sg13g2_xnor2_1 _08039_ (.Y(_02773_),
    .A(_02522_),
    .B(_02604_));
 sg13g2_xnor2_1 _08040_ (.Y(_02774_),
    .A(net30),
    .B(_02773_));
 sg13g2_xnor2_1 _08041_ (.Y(_02775_),
    .A(_02382_),
    .B(_02774_));
 sg13g2_xnor2_1 _08042_ (.Y(_02776_),
    .A(_02750_),
    .B(_02775_));
 sg13g2_nand2_1 _08043_ (.Y(_02777_),
    .A(_02146_),
    .B(_02776_));
 sg13g2_a21o_1 _08044_ (.A2(_02772_),
    .A1(_02763_),
    .B1(_02777_),
    .X(_02778_));
 sg13g2_mux2_1 _08045_ (.A0(_02773_),
    .A1(_02766_),
    .S(net30),
    .X(_02779_));
 sg13g2_nand2b_1 _08046_ (.Y(_02780_),
    .B(_02748_),
    .A_N(_02779_));
 sg13g2_a21oi_1 _08047_ (.A1(_02761_),
    .A2(_02770_),
    .Y(_02781_),
    .B1(_02750_));
 sg13g2_nand2b_1 _08048_ (.Y(_02782_),
    .B(_02770_),
    .A_N(_02382_));
 sg13g2_a221oi_1 _08049_ (.B2(_02750_),
    .C1(_02752_),
    .B1(_02782_),
    .A1(_02780_),
    .Y(_02783_),
    .A2(_02781_));
 sg13g2_a21o_1 _08050_ (.A2(_02752_),
    .A1(_02748_),
    .B1(_02765_),
    .X(_02784_));
 sg13g2_and2_1 _08051_ (.A(net30),
    .B(_02773_),
    .X(_02785_));
 sg13g2_nor2_1 _08052_ (.A(net30),
    .B(_02767_),
    .Y(_02786_));
 sg13g2_nor3_1 _08053_ (.A(_02146_),
    .B(_02785_),
    .C(_02786_),
    .Y(_02787_));
 sg13g2_a22oi_1 _08054_ (.Y(_02788_),
    .B1(_02784_),
    .B2(_02787_),
    .A2(_02783_),
    .A1(_02269_));
 sg13g2_and4_1 _08055_ (.A(_02569_),
    .B(_02684_),
    .C(_02778_),
    .D(_02788_),
    .X(_02789_));
 sg13g2_buf_2 fanout435 (.A(net439),
    .X(net435));
 sg13g2_inv_1 _08057_ (.Y(_02791_),
    .A(net19));
 sg13g2_xor2_1 _08058_ (.B(net22),
    .A(_02463_),
    .X(_02792_));
 sg13g2_xnor2_1 _08059_ (.Y(_02793_),
    .A(net25),
    .B(_02311_));
 sg13g2_xnor2_1 _08060_ (.Y(_02794_),
    .A(_02792_),
    .B(_02793_));
 sg13g2_o21ai_1 _08061_ (.B1(_01998_),
    .Y(_02795_),
    .A1(net109),
    .A2(_01999_));
 sg13g2_nor2_1 _08062_ (.A(net109),
    .B(_01999_),
    .Y(_02796_));
 sg13g2_a21o_1 _08063_ (.A2(_02796_),
    .A1(net186),
    .B1(_02053_),
    .X(_02797_));
 sg13g2_nand2_1 _08064_ (.Y(_02798_),
    .A(net81),
    .B(net55));
 sg13g2_nand2_1 _08065_ (.Y(_02799_),
    .A(net55),
    .B(net59));
 sg13g2_nor2b_1 _08066_ (.A(net129),
    .B_N(net191),
    .Y(_02800_));
 sg13g2_a21oi_1 _08067_ (.A1(_02176_),
    .A2(net194),
    .Y(_02801_),
    .B1(_02800_));
 sg13g2_nor2_1 _08068_ (.A(_02176_),
    .B(net194),
    .Y(_02802_));
 sg13g2_nor2b_1 _08069_ (.A(net197),
    .B_N(net75),
    .Y(_02803_));
 sg13g2_o21ai_1 _08070_ (.B1(net74),
    .Y(_02804_),
    .A1(_02174_),
    .A2(_02803_));
 sg13g2_a221oi_1 _08071_ (.B2(_02174_),
    .C1(_02800_),
    .B1(_02803_),
    .A1(_02176_),
    .Y(_02805_),
    .A2(net194));
 sg13g2_nand2b_1 _08072_ (.Y(_02806_),
    .B(net109),
    .A_N(net189));
 sg13g2_nand2b_1 _08073_ (.Y(_02807_),
    .B(\median_processor.input_storage[5] ),
    .A_N(net187));
 sg13g2_nand2b_1 _08074_ (.Y(_02808_),
    .B(net129),
    .A_N(net191));
 sg13g2_nand3_1 _08075_ (.B(_02807_),
    .C(_02808_),
    .A(_02806_),
    .Y(_02809_));
 sg13g2_a221oi_1 _08076_ (.B2(_02805_),
    .C1(_02809_),
    .B1(_02804_),
    .A1(_02801_),
    .Y(_02810_),
    .A2(_02802_));
 sg13g2_a221oi_1 _08077_ (.B2(_02799_),
    .C1(_02810_),
    .B1(_02798_),
    .A1(_02795_),
    .Y(_02811_),
    .A2(_02797_));
 sg13g2_buf_1 fanout434 (.A(net493),
    .X(net434));
 sg13g2_nor2_1 _08079_ (.A(net184),
    .B(_02798_),
    .Y(_02813_));
 sg13g2_nand2_1 _08080_ (.Y(_02814_),
    .A(net57),
    .B(_02708_));
 sg13g2_nor3_1 _08081_ (.A(_02811_),
    .B(_02813_),
    .C(_02814_),
    .Y(_02815_));
 sg13g2_nor2_1 _08082_ (.A(net56),
    .B(net184),
    .Y(_02816_));
 sg13g2_a221oi_1 _08083_ (.B2(_02797_),
    .C1(_02810_),
    .B1(_02795_),
    .A1(net56),
    .Y(_02817_),
    .A2(net184));
 sg13g2_nor4_1 _08084_ (.A(_02250_),
    .B(net53),
    .C(_02816_),
    .D(_02817_),
    .Y(_02818_));
 sg13g2_o21ai_1 _08085_ (.B1(_02705_),
    .Y(_02819_),
    .A1(_02815_),
    .A2(_02818_));
 sg13g2_nand2_1 _08086_ (.Y(_02820_),
    .A(net79),
    .B(net59));
 sg13g2_nand2_1 _08087_ (.Y(_02821_),
    .A(net79),
    .B(net81));
 sg13g2_a221oi_1 _08088_ (.B2(_02821_),
    .C1(_02810_),
    .B1(_02820_),
    .A1(_02795_),
    .Y(_02822_),
    .A2(_02797_));
 sg13g2_buf_2 fanout433 (.A(net434),
    .X(net433));
 sg13g2_nand2_1 _08090_ (.Y(_02824_),
    .A(net79),
    .B(net55));
 sg13g2_o21ai_1 _08091_ (.B1(_02824_),
    .Y(_02825_),
    .A1(net184),
    .A2(_02821_));
 sg13g2_or4_2 _08092_ (.A(_02811_),
    .B(_02813_),
    .C(_02822_),
    .D(_02825_),
    .X(_02826_));
 sg13g2_buf_1 fanout432 (.A(net433),
    .X(net432));
 sg13g2_nor3_1 _08094_ (.A(_02058_),
    .B(_02250_),
    .C(net165),
    .Y(_02828_));
 sg13g2_or2_1 _08095_ (.X(_02829_),
    .B(_02817_),
    .A(_02816_));
 sg13g2_buf_1 fanout431 (.A(net432),
    .X(net431));
 sg13g2_a22oi_1 _08097_ (.Y(_02831_),
    .B1(_02828_),
    .B2(_02829_),
    .A2(_02826_),
    .A1(_02730_));
 sg13g2_and2_1 _08098_ (.A(_02819_),
    .B(_02831_),
    .X(_02832_));
 sg13g2_buf_1 fanout430 (.A(net432),
    .X(net430));
 sg13g2_nor3_1 _08100_ (.A(_02791_),
    .B(_02794_),
    .C(_02832_),
    .Y(_02834_));
 sg13g2_o21ai_1 _08101_ (.B1(net165),
    .Y(_02835_),
    .A1(_02816_),
    .A2(_02817_));
 sg13g2_a21oi_1 _08102_ (.A1(net181),
    .A2(_02835_),
    .Y(_02836_),
    .B1(_02058_));
 sg13g2_a21o_1 _08103_ (.A2(_02829_),
    .A1(net55),
    .B1(_02836_),
    .X(_02837_));
 sg13g2_nand4_1 _08104_ (.B(_02705_),
    .C(_02794_),
    .A(net19),
    .Y(_02838_),
    .D(_02837_));
 sg13g2_nand2b_1 _08105_ (.Y(_02839_),
    .B(_02838_),
    .A_N(_02834_));
 sg13g2_nand2_1 _08106_ (.Y(_02840_),
    .A(_02311_),
    .B(_02463_));
 sg13g2_nand2_1 _08107_ (.Y(_02841_),
    .A(net22),
    .B(_02840_));
 sg13g2_nor3_1 _08108_ (.A(_02299_),
    .B(_02302_),
    .C(_02308_),
    .Y(_02842_));
 sg13g2_nand4_1 _08109_ (.B(_02309_),
    .C(_02438_),
    .A(_02842_),
    .Y(_02843_),
    .D(_02461_));
 sg13g2_a221oi_1 _08110_ (.B2(_02843_),
    .C1(net25),
    .B1(_02841_),
    .A1(_02819_),
    .Y(_02844_),
    .A2(_02831_));
 sg13g2_nand4_1 _08111_ (.B(_02461_),
    .C(_02641_),
    .A(_02438_),
    .Y(_02845_),
    .D(_02662_));
 sg13g2_or2_1 _08112_ (.X(_02846_),
    .B(_02845_),
    .A(_02311_));
 sg13g2_a21oi_1 _08113_ (.A1(net25),
    .A2(_02832_),
    .Y(_02847_),
    .B1(_02846_));
 sg13g2_or2_1 _08114_ (.X(_02848_),
    .B(_02847_),
    .A(_02844_));
 sg13g2_and2_1 _08115_ (.A(net25),
    .B(_02311_),
    .X(_02849_));
 sg13g2_nor2b_1 _08116_ (.A(_02463_),
    .B_N(net22),
    .Y(_02850_));
 sg13g2_a22oi_1 _08117_ (.Y(_02851_),
    .B1(_02641_),
    .B2(_02662_),
    .A2(_02461_),
    .A1(_02438_));
 sg13g2_nor2_1 _08118_ (.A(net26),
    .B(_02311_),
    .Y(_02852_));
 sg13g2_nor2_1 _08119_ (.A(_02792_),
    .B(_02793_),
    .Y(_02853_));
 sg13g2_a221oi_1 _08120_ (.B2(_02852_),
    .C1(_02853_),
    .B1(_02851_),
    .A1(_02849_),
    .Y(_02854_),
    .A2(_02850_));
 sg13g2_inv_1 _08121_ (.Y(_02855_),
    .A(_02854_));
 sg13g2_nor2_1 _08122_ (.A(_02822_),
    .B(_02825_),
    .Y(_02856_));
 sg13g2_nand2_1 _08123_ (.Y(_02857_),
    .A(_02705_),
    .B(_02708_));
 sg13g2_nand2b_1 _08124_ (.Y(_02858_),
    .B(_02857_),
    .A_N(net19));
 sg13g2_nand2_1 _08125_ (.Y(_02859_),
    .A(net165),
    .B(_02705_));
 sg13g2_nand2b_1 _08126_ (.Y(_02860_),
    .B(net19),
    .A_N(_02859_));
 sg13g2_nand3_1 _08127_ (.B(_02858_),
    .C(_02860_),
    .A(_02856_),
    .Y(_02861_));
 sg13g2_a21oi_1 _08128_ (.A1(net19),
    .A2(_02705_),
    .Y(_02862_),
    .B1(_02829_));
 sg13g2_nor2_1 _08129_ (.A(net181),
    .B(_02862_),
    .Y(_02863_));
 sg13g2_nand3_1 _08130_ (.B(_02826_),
    .C(_02857_),
    .A(_02791_),
    .Y(_02864_));
 sg13g2_o21ai_1 _08131_ (.B1(_02864_),
    .Y(_02865_),
    .A1(_02861_),
    .A2(_02863_));
 sg13g2_a21o_1 _08132_ (.A2(_02845_),
    .A1(net25),
    .B1(_02851_),
    .X(_02866_));
 sg13g2_o21ai_1 _08133_ (.B1(_02250_),
    .Y(_02867_),
    .A1(_02705_),
    .A2(_02829_));
 sg13g2_nor2b_1 _08134_ (.A(net19),
    .B_N(_02859_),
    .Y(_02868_));
 sg13g2_nand4_1 _08135_ (.B(_02866_),
    .C(_02867_),
    .A(_02856_),
    .Y(_02869_),
    .D(_02868_));
 sg13g2_nand2_1 _08136_ (.Y(_02870_),
    .A(_02819_),
    .B(_02831_));
 sg13g2_a22oi_1 _08137_ (.Y(_02871_),
    .B1(_02866_),
    .B2(_02311_),
    .A2(_02851_),
    .A1(net25));
 sg13g2_nor4_2 _08138_ (.A(_02811_),
    .B(_02813_),
    .C(_02822_),
    .Y(_02872_),
    .D(_02825_));
 sg13g2_nor3_1 _08139_ (.A(net19),
    .B(_02872_),
    .C(_02857_),
    .Y(_02873_));
 sg13g2_o21ai_1 _08140_ (.B1(_02873_),
    .Y(_02874_),
    .A1(_02870_),
    .A2(_02871_));
 sg13g2_nand2_1 _08141_ (.Y(_02875_),
    .A(net25),
    .B(_02840_));
 sg13g2_xor2_1 _08142_ (.B(net22),
    .A(net25),
    .X(_02876_));
 sg13g2_a21oi_1 _08143_ (.A1(_02843_),
    .A2(_02840_),
    .Y(_02877_),
    .B1(_02876_));
 sg13g2_o21ai_1 _08144_ (.B1(_02877_),
    .Y(_02878_),
    .A1(_02832_),
    .A2(_02875_));
 sg13g2_nand3_1 _08145_ (.B(_02840_),
    .C(_02876_),
    .A(_02843_),
    .Y(_02879_));
 sg13g2_a22oi_1 _08146_ (.Y(_02880_),
    .B1(_02878_),
    .B2(_02879_),
    .A2(_02874_),
    .A1(_02869_));
 sg13g2_a221oi_1 _08147_ (.B2(_02865_),
    .C1(_02880_),
    .B1(_02855_),
    .A1(_02839_),
    .Y(_02881_),
    .A2(_02848_));
 sg13g2_buf_1 fanout429 (.A(net432),
    .X(net429));
 sg13g2_mux2_1 _08149_ (.A0(net75),
    .A1(net197),
    .S(net8),
    .X(_02883_));
 sg13g2_inv_1 _08150_ (.Y(_02884_),
    .A(_02883_));
 sg13g2_nand2_1 _08151_ (.Y(_02885_),
    .A(_02569_),
    .B(_02684_));
 sg13g2_a21oi_2 _08152_ (.B1(_02885_),
    .Y(_02886_),
    .A2(_02788_),
    .A1(_02778_));
 sg13g2_buf_1 fanout428 (.A(net434),
    .X(net428));
 sg13g2_inv_1 _08154_ (.Y(_02888_),
    .A(net179));
 sg13g2_nand2b_2 _08155_ (.Y(_02889_),
    .B(_02683_),
    .A_N(_02666_));
 sg13g2_buf_1 fanout427 (.A(net428),
    .X(net427));
 sg13g2_nor3_1 _08157_ (.A(net163),
    .B(net10),
    .C(_02889_),
    .Y(_02891_));
 sg13g2_nor2_1 _08158_ (.A(net145),
    .B(net9),
    .Y(_02892_));
 sg13g2_or2_2 _08159_ (.X(_02893_),
    .B(net11),
    .A(net12));
 sg13g2_buf_2 fanout426 (.A(net427),
    .X(net426));
 sg13g2_or3_1 _08161_ (.A(_02891_),
    .B(_02892_),
    .C(_02893_),
    .X(_02895_));
 sg13g2_a221oi_1 _08162_ (.B2(_02888_),
    .C1(_02895_),
    .B1(_02886_),
    .A1(net6),
    .Y(_02896_),
    .A2(_02884_));
 sg13g2_nor3_1 _08163_ (.A(_02281_),
    .B(_02427_),
    .C(_02896_),
    .Y(_02897_));
 sg13g2_or2_1 _08164_ (.X(_02898_),
    .B(_02426_),
    .A(_02420_));
 sg13g2_buf_1 fanout425 (.A(net427),
    .X(net425));
 sg13g2_nor3_1 _08166_ (.A(net24),
    .B(_02486_),
    .C(_02629_),
    .Y(_02900_));
 sg13g2_nand2_1 _08167_ (.Y(_02901_),
    .A(net24),
    .B(_02826_));
 sg13g2_nand2_1 _08168_ (.Y(_02902_),
    .A(_02486_),
    .B(_02629_));
 sg13g2_nor2_1 _08169_ (.A(_02901_),
    .B(_02902_),
    .Y(_02903_));
 sg13g2_a21oi_1 _08170_ (.A1(_02872_),
    .A2(_02900_),
    .Y(_02904_),
    .B1(_02903_));
 sg13g2_xnor2_1 _08171_ (.Y(_02905_),
    .A(net24),
    .B(_02872_));
 sg13g2_nand4_1 _08172_ (.B(_02486_),
    .C(_02629_),
    .A(net20),
    .Y(_02906_),
    .D(_02905_));
 sg13g2_o21ai_1 _08173_ (.B1(_02906_),
    .Y(_02907_),
    .A1(net20),
    .A2(_02904_));
 sg13g2_a21oi_2 _08174_ (.B1(_02192_),
    .Y(_02908_),
    .A2(_02187_),
    .A1(_02184_));
 sg13g2_nor3_1 _08175_ (.A(net24),
    .B(_02908_),
    .C(_02826_),
    .Y(_02909_));
 sg13g2_a21oi_1 _08176_ (.A1(_02908_),
    .A2(_02905_),
    .Y(_02910_),
    .B1(_02909_));
 sg13g2_xnor2_1 _08177_ (.Y(_02911_),
    .A(_02486_),
    .B(_02629_));
 sg13g2_o21ai_1 _08178_ (.B1(net56),
    .Y(_02912_),
    .A1(net168),
    .A2(_02727_));
 sg13g2_a22oi_1 _08179_ (.Y(_02913_),
    .B1(_02729_),
    .B2(_02912_),
    .A2(net53),
    .A1(net78));
 sg13g2_nor2_1 _08180_ (.A(_02707_),
    .B(_02913_),
    .Y(_02914_));
 sg13g2_o21ai_1 _08181_ (.B1(_02914_),
    .Y(_02915_),
    .A1(_02910_),
    .A2(_02911_));
 sg13g2_nor2_1 _08182_ (.A(_02486_),
    .B(_02629_),
    .Y(_02916_));
 sg13g2_a21o_1 _08183_ (.A2(_02905_),
    .A1(_02908_),
    .B1(_02909_),
    .X(_02917_));
 sg13g2_nand2_1 _08184_ (.Y(_02918_),
    .A(net20),
    .B(_02905_));
 sg13g2_nand2b_1 _08185_ (.Y(_02919_),
    .B(_02908_),
    .A_N(_02901_));
 sg13g2_a21oi_1 _08186_ (.A1(_02918_),
    .A2(_02919_),
    .Y(_02920_),
    .B1(_02911_));
 sg13g2_a221oi_1 _08187_ (.B2(net20),
    .C1(_02920_),
    .B1(_02903_),
    .A1(_02916_),
    .Y(_02921_),
    .A2(_02917_));
 sg13g2_nand2b_1 _08188_ (.Y(_02922_),
    .B(_02921_),
    .A_N(_02914_));
 sg13g2_o21ai_1 _08189_ (.B1(_02922_),
    .Y(_02923_),
    .A1(_02907_),
    .A2(_02915_));
 sg13g2_or2_1 _08190_ (.X(_02924_),
    .B(_02916_),
    .A(net24));
 sg13g2_nand4_1 _08191_ (.B(_02826_),
    .C(_02902_),
    .A(net20),
    .Y(_02925_),
    .D(_02924_));
 sg13g2_xnor2_1 _08192_ (.Y(_02926_),
    .A(_02908_),
    .B(_02826_));
 sg13g2_nand3_1 _08193_ (.B(_02924_),
    .C(_02926_),
    .A(_02902_),
    .Y(_02927_));
 sg13g2_xnor2_1 _08194_ (.Y(_02928_),
    .A(net24),
    .B(_02911_));
 sg13g2_mux2_1 _08195_ (.A0(_02925_),
    .A1(_02927_),
    .S(_02928_),
    .X(_02929_));
 sg13g2_mux2_1 _08196_ (.A0(_02929_),
    .A1(_02921_),
    .S(_02914_),
    .X(_02930_));
 sg13g2_mux2_1 _08197_ (.A0(_02923_),
    .A1(_02930_),
    .S(_02331_),
    .X(_02931_));
 sg13g2_inv_1 _08198_ (.Y(_02932_),
    .A(_02881_));
 sg13g2_nor3_1 _08199_ (.A(net14),
    .B(net11),
    .C(_02932_),
    .Y(_02933_));
 sg13g2_nand4_1 _08200_ (.B(_02789_),
    .C(_02931_),
    .A(_02898_),
    .Y(_02934_),
    .D(_02933_));
 sg13g2_buf_2 fanout424 (.A(net427),
    .X(net424));
 sg13g2_buf_2 fanout423 (.A(net428),
    .X(net423));
 sg13g2_o21ai_1 _08203_ (.B1(net3),
    .Y(_02937_),
    .A1(net96),
    .A2(net5));
 sg13g2_inv_1 _08204_ (.Y(_02938_),
    .A(\median_processor.median_processor.median_out[0] ));
 sg13g2_or2_1 _08205_ (.X(_02939_),
    .B(net3),
    .A(_02938_));
 sg13g2_o21ai_1 _08206_ (.B1(_02939_),
    .Y(_00064_),
    .A1(_02897_),
    .A2(_02937_));
 sg13g2_nand2_1 _08207_ (.Y(_02940_),
    .A(\median_processor.input_storage[41] ),
    .B(net11));
 sg13g2_nand2_1 _08208_ (.Y(_02941_),
    .A(net110),
    .B(net12));
 sg13g2_o21ai_1 _08209_ (.B1(_02941_),
    .Y(_02942_),
    .A1(net12),
    .A2(_02940_));
 sg13g2_mux2_1 _08210_ (.A0(net74),
    .A1(\median_processor.input_storage[1] ),
    .S(net8),
    .X(_02943_));
 sg13g2_inv_1 _08211_ (.Y(_02944_),
    .A(_02943_));
 sg13g2_nor3_1 _08212_ (.A(net161),
    .B(net10),
    .C(_02889_),
    .Y(_02945_));
 sg13g2_nor2_1 _08213_ (.A(net142),
    .B(net9),
    .Y(_02946_));
 sg13g2_or3_1 _08214_ (.A(_02893_),
    .B(_02945_),
    .C(_02946_),
    .X(_02947_));
 sg13g2_a221oi_1 _08215_ (.B2(net6),
    .C1(_02947_),
    .B1(_02944_),
    .A1(_02503_),
    .Y(_02948_),
    .A2(_02886_));
 sg13g2_nor3_1 _08216_ (.A(_02427_),
    .B(_02942_),
    .C(_02948_),
    .Y(_02949_));
 sg13g2_o21ai_1 _08217_ (.B1(net3),
    .Y(_02950_),
    .A1(net94),
    .A2(net5));
 sg13g2_buf_2 fanout422 (.A(net423),
    .X(net422));
 sg13g2_inv_1 _08219_ (.Y(_02952_),
    .A(\median_processor.median_processor.median_out[1] ));
 sg13g2_or2_1 _08220_ (.X(_02953_),
    .B(net3),
    .A(_02952_));
 sg13g2_o21ai_1 _08221_ (.B1(_02953_),
    .Y(_00065_),
    .A1(_02949_),
    .A2(_02950_));
 sg13g2_nand2_1 _08222_ (.Y(_02954_),
    .A(net125),
    .B(net11));
 sg13g2_nand2_1 _08223_ (.Y(_02955_),
    .A(net108),
    .B(net12));
 sg13g2_o21ai_1 _08224_ (.B1(_02955_),
    .Y(_02956_),
    .A1(net12),
    .A2(_02954_));
 sg13g2_mux2_1 _08225_ (.A0(net195),
    .A1(net151),
    .S(net8),
    .X(_02957_));
 sg13g2_inv_1 _08226_ (.Y(_02958_),
    .A(_02957_));
 sg13g2_nor3_1 _08227_ (.A(net160),
    .B(net10),
    .C(_02889_),
    .Y(_02959_));
 sg13g2_nor2_1 _08228_ (.A(net141),
    .B(net9),
    .Y(_02960_));
 sg13g2_or3_1 _08229_ (.A(_02893_),
    .B(_02959_),
    .C(_02960_),
    .X(_02961_));
 sg13g2_a221oi_1 _08230_ (.B2(net6),
    .C1(_02961_),
    .B1(_02958_),
    .A1(_02579_),
    .Y(_02962_),
    .A2(_02886_));
 sg13g2_nor3_1 _08231_ (.A(_02427_),
    .B(_02956_),
    .C(_02962_),
    .Y(_02963_));
 sg13g2_o21ai_1 _08232_ (.B1(net3),
    .Y(_02964_),
    .A1(net92),
    .A2(net5));
 sg13g2_buf_2 fanout421 (.A(net428),
    .X(net421));
 sg13g2_inv_1 _08234_ (.Y(_02966_),
    .A(\median_processor.median_processor.median_out[2] ));
 sg13g2_or2_1 _08235_ (.X(_02967_),
    .B(net3),
    .A(_02966_));
 sg13g2_o21ai_1 _08236_ (.B1(_02967_),
    .Y(_00066_),
    .A1(_02963_),
    .A2(_02964_));
 sg13g2_nand2_1 _08237_ (.Y(_02968_),
    .A(net124),
    .B(net11));
 sg13g2_nand2_1 _08238_ (.Y(_02969_),
    .A(net106),
    .B(net12));
 sg13g2_o21ai_1 _08239_ (.B1(_02969_),
    .Y(_02970_),
    .A1(net13),
    .A2(_02968_));
 sg13g2_mux2_1 _08240_ (.A0(net191),
    .A1(net128),
    .S(net8),
    .X(_02971_));
 sg13g2_inv_1 _08241_ (.Y(_02972_),
    .A(_02971_));
 sg13g2_nor3_1 _08242_ (.A(net158),
    .B(net10),
    .C(_02889_),
    .Y(_02973_));
 sg13g2_nor2_1 _08243_ (.A(net139),
    .B(net9),
    .Y(_02974_));
 sg13g2_or3_1 _08244_ (.A(_02893_),
    .B(_02973_),
    .C(_02974_),
    .X(_02975_));
 sg13g2_a221oi_1 _08245_ (.B2(net6),
    .C1(_02975_),
    .B1(_02972_),
    .A1(_01895_),
    .Y(_02976_),
    .A2(_02886_));
 sg13g2_nor3_1 _08246_ (.A(_02427_),
    .B(_02970_),
    .C(_02976_),
    .Y(_02977_));
 sg13g2_o21ai_1 _08247_ (.B1(net3),
    .Y(_02978_),
    .A1(net91),
    .A2(net5));
 sg13g2_inv_1 _08248_ (.Y(_02979_),
    .A(\median_processor.median_processor.median_out[3] ));
 sg13g2_or2_1 _08249_ (.X(_02980_),
    .B(net3),
    .A(_02979_));
 sg13g2_o21ai_1 _08250_ (.B1(_02980_),
    .Y(_00067_),
    .A1(_02977_),
    .A2(_02978_));
 sg13g2_nand2_1 _08251_ (.Y(_02981_),
    .A(net122),
    .B(net11));
 sg13g2_nand2_1 _08252_ (.Y(_02982_),
    .A(net103),
    .B(net13));
 sg13g2_o21ai_1 _08253_ (.B1(_02982_),
    .Y(_02983_),
    .A1(net13),
    .A2(_02981_));
 sg13g2_mux2_1 _08254_ (.A0(net189),
    .A1(net109),
    .S(net8),
    .X(_02984_));
 sg13g2_inv_1 _08255_ (.Y(_02985_),
    .A(_02984_));
 sg13g2_nor3_1 _08256_ (.A(net156),
    .B(net10),
    .C(_02889_),
    .Y(_02986_));
 sg13g2_nor2_1 _08257_ (.A(net136),
    .B(net9),
    .Y(_02987_));
 sg13g2_or3_1 _08258_ (.A(_02893_),
    .B(_02986_),
    .C(_02987_),
    .X(_02988_));
 sg13g2_a221oi_1 _08259_ (.B2(net6),
    .C1(_02988_),
    .B1(_02985_),
    .A1(_01877_),
    .Y(_02989_),
    .A2(_02886_));
 sg13g2_nor3_1 _08260_ (.A(_02427_),
    .B(_02983_),
    .C(_02989_),
    .Y(_02990_));
 sg13g2_o21ai_1 _08261_ (.B1(net4),
    .Y(_02991_),
    .A1(net87),
    .A2(net5));
 sg13g2_buf_2 fanout420 (.A(net421),
    .X(net420));
 sg13g2_inv_1 _08263_ (.Y(_02993_),
    .A(\median_processor.median_processor.median_out[4] ));
 sg13g2_or2_1 _08264_ (.X(_02994_),
    .B(net4),
    .A(_02993_));
 sg13g2_o21ai_1 _08265_ (.B1(_02994_),
    .Y(_00068_),
    .A1(_02990_),
    .A2(_02991_));
 sg13g2_nand2_1 _08266_ (.Y(_02995_),
    .A(net118),
    .B(net11));
 sg13g2_nand2_1 _08267_ (.Y(_02996_),
    .A(net101),
    .B(net13));
 sg13g2_o21ai_1 _08268_ (.B1(_02996_),
    .Y(_02997_),
    .A1(net13),
    .A2(_02995_));
 sg13g2_mux2_1 _08269_ (.A0(net187),
    .A1(net89),
    .S(net8),
    .X(_02998_));
 sg13g2_inv_1 _08270_ (.Y(_02999_),
    .A(_02998_));
 sg13g2_nor3_1 _08271_ (.A(net154),
    .B(net10),
    .C(_02889_),
    .Y(_03000_));
 sg13g2_nor2_1 _08272_ (.A(net134),
    .B(net9),
    .Y(_03001_));
 sg13g2_or3_1 _08273_ (.A(_02893_),
    .B(_03000_),
    .C(_03001_),
    .X(_03002_));
 sg13g2_a221oi_1 _08274_ (.B2(net6),
    .C1(_03002_),
    .B1(_02999_),
    .A1(_01873_),
    .Y(_03003_),
    .A2(_02886_));
 sg13g2_nor3_1 _08275_ (.A(_02427_),
    .B(_02997_),
    .C(_03003_),
    .Y(_03004_));
 sg13g2_o21ai_1 _08276_ (.B1(net4),
    .Y(_03005_),
    .A1(net86),
    .A2(net5));
 sg13g2_inv_1 _08277_ (.Y(_03006_),
    .A(\median_processor.median_processor.median_out[5] ));
 sg13g2_or2_1 _08278_ (.X(_03007_),
    .B(_02934_),
    .A(_03006_));
 sg13g2_o21ai_1 _08279_ (.B1(_03007_),
    .Y(_00069_),
    .A1(_03004_),
    .A2(_03005_));
 sg13g2_nand2_1 _08280_ (.Y(_03008_),
    .A(net117),
    .B(_02277_));
 sg13g2_nand2_1 _08281_ (.Y(_03009_),
    .A(net99),
    .B(net14));
 sg13g2_o21ai_1 _08282_ (.B1(_03009_),
    .Y(_03010_),
    .A1(net14),
    .A2(_03008_));
 sg13g2_mux2_1 _08283_ (.A0(net184),
    .A1(net80),
    .S(net8),
    .X(_03011_));
 sg13g2_inv_1 _08284_ (.Y(_03012_),
    .A(_03011_));
 sg13g2_nor3_1 _08285_ (.A(net149),
    .B(net10),
    .C(_02889_),
    .Y(_03013_));
 sg13g2_nor2_1 _08286_ (.A(net132),
    .B(net9),
    .Y(_03014_));
 sg13g2_or3_1 _08287_ (.A(_02893_),
    .B(_03013_),
    .C(_03014_),
    .X(_03015_));
 sg13g2_a221oi_1 _08288_ (.B2(net6),
    .C1(_03015_),
    .B1(_03012_),
    .A1(_02364_),
    .Y(_03016_),
    .A2(_02886_));
 sg13g2_nor3_1 _08289_ (.A(_02427_),
    .B(_03010_),
    .C(_03016_),
    .Y(_03017_));
 sg13g2_o21ai_1 _08290_ (.B1(net4),
    .Y(_03018_),
    .A1(net84),
    .A2(net5));
 sg13g2_inv_1 _08291_ (.Y(_03019_),
    .A(\median_processor.median_processor.median_out[6] ));
 sg13g2_or2_1 _08292_ (.X(_03020_),
    .B(net4),
    .A(_03019_));
 sg13g2_o21ai_1 _08293_ (.B1(_03020_),
    .Y(_00070_),
    .A1(_03017_),
    .A2(_03018_));
 sg13g2_nand2_1 _08294_ (.Y(_03021_),
    .A(net113),
    .B(_02277_));
 sg13g2_nand2_1 _08295_ (.Y(_03022_),
    .A(net97),
    .B(net14));
 sg13g2_o21ai_1 _08296_ (.B1(_03022_),
    .Y(_03023_),
    .A1(net14),
    .A2(_03021_));
 sg13g2_mux2_1 _08297_ (.A0(net181),
    .A1(net78),
    .S(net8),
    .X(_03024_));
 sg13g2_inv_1 _08298_ (.Y(_03025_),
    .A(_03024_));
 sg13g2_nor3_1 _08299_ (.A(net146),
    .B(net10),
    .C(_02889_),
    .Y(_03026_));
 sg13g2_nor2_1 _08300_ (.A(net130),
    .B(net9),
    .Y(_03027_));
 sg13g2_or3_1 _08301_ (.A(_02893_),
    .B(_03026_),
    .C(_03027_),
    .X(_03028_));
 sg13g2_a221oi_1 _08302_ (.B2(net6),
    .C1(_03028_),
    .B1(_03025_),
    .A1(net53),
    .Y(_03029_),
    .A2(_02886_));
 sg13g2_nor3_1 _08303_ (.A(_02427_),
    .B(_03023_),
    .C(_03029_),
    .Y(_03030_));
 sg13g2_o21ai_1 _08304_ (.B1(net4),
    .Y(_03031_),
    .A1(net83),
    .A2(net5));
 sg13g2_inv_1 _08305_ (.Y(_03032_),
    .A(\median_processor.median_processor.median_out[7] ));
 sg13g2_or2_1 _08306_ (.X(_03033_),
    .B(net4),
    .A(_03032_));
 sg13g2_o21ai_1 _08307_ (.B1(_03033_),
    .Y(_00071_),
    .A1(_03030_),
    .A2(_03031_));
 sg13g2_buf_1 fanout419 (.A(net421),
    .X(net419));
 sg13g2_buf_1 fanout418 (.A(net434),
    .X(net418));
 sg13g2_buf_1 fanout417 (.A(net418),
    .X(net417));
 sg13g2_buf_1 fanout416 (.A(net417),
    .X(net416));
 sg13g2_inv_1 _08312_ (.Y(_03038_),
    .A(data_in_p2c_1));
 sg13g2_nand2b_1 _08313_ (.Y(_03039_),
    .B(\median_processor.wr_enable ),
    .A_N(reg_addr_p2c_1));
 sg13g2_nor2_1 _08314_ (.A(reg_addr_p2c_3),
    .B(reg_addr_p2c_2),
    .Y(_03040_));
 sg13g2_nand2b_1 _08315_ (.Y(_03041_),
    .B(_03040_),
    .A_N(_03039_));
 sg13g2_buf_1 fanout415 (.A(net416),
    .X(net415));
 sg13g2_buf_2 fanout414 (.A(net416),
    .X(net414));
 sg13g2_nand2_1 _08318_ (.Y(_03044_),
    .A(net197),
    .B(net51));
 sg13g2_o21ai_1 _08319_ (.B1(_03044_),
    .Y(_03045_),
    .A1(_03038_),
    .A2(net51));
 sg13g2_and2_1 _08320_ (.A(net451),
    .B(_03045_),
    .X(_00000_));
 sg13g2_nand3_1 _08321_ (.B(\median_processor.wr_enable ),
    .C(_03040_),
    .A(reg_addr_p2c_1),
    .Y(_03046_));
 sg13g2_buf_2 fanout413 (.A(net414),
    .X(net413));
 sg13g2_buf_1 fanout412 (.A(net416),
    .X(net412));
 sg13g2_buf_1 fanout411 (.A(net416),
    .X(net411));
 sg13g2_inv_2 _08325_ (.Y(_03050_),
    .A(data_in_p2c_3));
 sg13g2_nor2_1 _08326_ (.A(_03050_),
    .B(net49),
    .Y(_03051_));
 sg13g2_a21oi_1 _08327_ (.A1(net194),
    .A2(net49),
    .Y(_03052_),
    .B1(_03051_));
 sg13g2_buf_1 fanout410 (.A(net417),
    .X(net410));
 sg13g2_buf_1 fanout409 (.A(net410),
    .X(net409));
 sg13g2_nor2b_1 _08330_ (.A(_03052_),
    .B_N(net452),
    .Y(_00001_));
 sg13g2_buf_2 fanout408 (.A(net410),
    .X(net408));
 sg13g2_inv_1 _08332_ (.Y(_03056_),
    .A(net503));
 sg13g2_nor2_1 _08333_ (.A(_03056_),
    .B(net49),
    .Y(_03057_));
 sg13g2_a21oi_1 _08334_ (.A1(net193),
    .A2(net49),
    .Y(_03058_),
    .B1(_03057_));
 sg13g2_nor2b_1 _08335_ (.A(_03058_),
    .B_N(net452),
    .Y(_00002_));
 sg13g2_buf_2 fanout407 (.A(net417),
    .X(net407));
 sg13g2_buf_2 fanout406 (.A(net407),
    .X(net406));
 sg13g2_mux2_1 _08338_ (.A0(net502),
    .A1(net189),
    .S(net49),
    .X(_03061_));
 sg13g2_and2_1 _08339_ (.A(net477),
    .B(_03061_),
    .X(_00003_));
 sg13g2_buf_1 fanout405 (.A(net418),
    .X(net405));
 sg13g2_inv_1 _08341_ (.Y(_03063_),
    .A(net500));
 sg13g2_nor2_1 _08342_ (.A(_03063_),
    .B(net50),
    .Y(_03064_));
 sg13g2_a21oi_1 _08343_ (.A1(net188),
    .A2(net50),
    .Y(_03065_),
    .B1(_03064_));
 sg13g2_nor2b_1 _08344_ (.A(_03065_),
    .B_N(net476),
    .Y(_00004_));
 sg13g2_buf_2 fanout404 (.A(net405),
    .X(net404));
 sg13g2_inv_1 _08346_ (.Y(_03067_),
    .A(net498));
 sg13g2_nor2_1 _08347_ (.A(_03067_),
    .B(net50),
    .Y(_03068_));
 sg13g2_a21oi_1 _08348_ (.A1(net185),
    .A2(net50),
    .Y(_03069_),
    .B1(_03068_));
 sg13g2_nor2b_1 _08349_ (.A(_03069_),
    .B_N(net478),
    .Y(_00005_));
 sg13g2_buf_2 fanout403 (.A(net404),
    .X(net403));
 sg13g2_inv_1 _08351_ (.Y(_03071_),
    .A(data_in_p2c_8));
 sg13g2_nor2_1 _08352_ (.A(_03071_),
    .B(net50),
    .Y(_03072_));
 sg13g2_a21oi_1 _08353_ (.A1(net181),
    .A2(net50),
    .Y(_03073_),
    .B1(_03072_));
 sg13g2_nor2b_1 _08354_ (.A(_03073_),
    .B_N(net479),
    .Y(_00006_));
 sg13g2_nand2b_1 _08355_ (.Y(_03074_),
    .B(reg_addr_p2c_2),
    .A_N(reg_addr_p2c_3));
 sg13g2_nor2_1 _08356_ (.A(_03039_),
    .B(_03074_),
    .Y(_03075_));
 sg13g2_buf_2 fanout402 (.A(net405),
    .X(net402));
 sg13g2_buf_2 fanout401 (.A(net402),
    .X(net401));
 sg13g2_nand2_1 _08359_ (.Y(_03078_),
    .A(data_in_p2c_1),
    .B(net46));
 sg13g2_o21ai_1 _08360_ (.B1(_03078_),
    .Y(_03079_),
    .A1(_02888_),
    .A2(net46));
 sg13g2_and2_1 _08361_ (.A(net469),
    .B(_03079_),
    .X(_00007_));
 sg13g2_buf_2 fanout400 (.A(net418),
    .X(net400));
 sg13g2_buf_2 fanout399 (.A(net400),
    .X(net399));
 sg13g2_nand2_1 _08364_ (.Y(_03082_),
    .A(net505),
    .B(net47));
 sg13g2_o21ai_1 _08365_ (.B1(_03082_),
    .Y(_03083_),
    .A1(_02503_),
    .A2(net46));
 sg13g2_and2_1 _08366_ (.A(net467),
    .B(_03083_),
    .X(_00008_));
 sg13g2_nand2_1 _08367_ (.Y(_03084_),
    .A(data_in_p2c_3),
    .B(net47));
 sg13g2_o21ai_1 _08368_ (.B1(_03084_),
    .Y(_03085_),
    .A1(_02579_),
    .A2(net47));
 sg13g2_and2_1 _08369_ (.A(net467),
    .B(_03085_),
    .X(_00009_));
 sg13g2_nand2_1 _08370_ (.Y(_03086_),
    .A(net503),
    .B(net46));
 sg13g2_o21ai_1 _08371_ (.B1(_03086_),
    .Y(_03087_),
    .A1(_01895_),
    .A2(net46));
 sg13g2_and2_1 _08372_ (.A(net467),
    .B(_03087_),
    .X(_00010_));
 sg13g2_mux2_1 _08373_ (.A0(net505),
    .A1(\median_processor.input_storage[1] ),
    .S(net51),
    .X(_03088_));
 sg13g2_and2_1 _08374_ (.A(net469),
    .B(_03088_),
    .X(_00011_));
 sg13g2_nand2_1 _08375_ (.Y(_03089_),
    .A(net502),
    .B(net46));
 sg13g2_o21ai_1 _08376_ (.B1(_03089_),
    .Y(_03090_),
    .A1(_01877_),
    .A2(net47));
 sg13g2_and2_1 _08377_ (.A(net484),
    .B(_03090_),
    .X(_00012_));
 sg13g2_nand2_1 _08378_ (.Y(_03091_),
    .A(data_in_p2c_6),
    .B(net46));
 sg13g2_o21ai_1 _08379_ (.B1(_03091_),
    .Y(_03092_),
    .A1(_01873_),
    .A2(net46));
 sg13g2_and2_1 _08380_ (.A(net477),
    .B(_03092_),
    .X(_00013_));
 sg13g2_nand2_1 _08381_ (.Y(_03093_),
    .A(net499),
    .B(net48));
 sg13g2_o21ai_1 _08382_ (.B1(_03093_),
    .Y(_03094_),
    .A1(_02364_),
    .A2(net48));
 sg13g2_and2_1 _08383_ (.A(net487),
    .B(_03094_),
    .X(_00014_));
 sg13g2_buf_1 fanout398 (.A(net493),
    .X(net398));
 sg13g2_nand2_1 _08385_ (.Y(_03096_),
    .A(data_in_p2c_8),
    .B(net48));
 sg13g2_o21ai_1 _08386_ (.B1(_03096_),
    .Y(_03097_),
    .A1(net53),
    .A2(net48));
 sg13g2_and2_1 _08387_ (.A(net487),
    .B(_03097_),
    .X(_00015_));
 sg13g2_nand2_1 _08388_ (.Y(_03098_),
    .A(reg_addr_p2c_1),
    .B(\median_processor.wr_enable ));
 sg13g2_nor2_1 _08389_ (.A(_03098_),
    .B(_03074_),
    .Y(_03099_));
 sg13g2_buf_1 fanout397 (.A(net398),
    .X(net397));
 sg13g2_nand2_1 _08391_ (.Y(_03101_),
    .A(data_in_p2c_1),
    .B(net45));
 sg13g2_o21ai_1 _08392_ (.B1(_03101_),
    .Y(_03102_),
    .A1(_02391_),
    .A2(net45));
 sg13g2_and2_1 _08393_ (.A(net469),
    .B(_03102_),
    .X(_00016_));
 sg13g2_nand2_1 _08394_ (.Y(_03103_),
    .A(net505),
    .B(net45));
 sg13g2_o21ai_1 _08395_ (.B1(_03103_),
    .Y(_03104_),
    .A1(_01709_),
    .A2(net45));
 sg13g2_and2_1 _08396_ (.A(net467),
    .B(_03104_),
    .X(_00017_));
 sg13g2_mux2_1 _08397_ (.A0(net159),
    .A1(data_in_p2c_3),
    .S(net45),
    .X(_03105_));
 sg13g2_and2_1 _08398_ (.A(net466),
    .B(_03105_),
    .X(_00018_));
 sg13g2_nand2_1 _08399_ (.Y(_03106_),
    .A(data_in_p2c_4),
    .B(net44));
 sg13g2_o21ai_1 _08400_ (.B1(_03106_),
    .Y(_03107_),
    .A1(_01719_),
    .A2(net44));
 sg13g2_and2_1 _08401_ (.A(net468),
    .B(_03107_),
    .X(_00019_));
 sg13g2_mux2_1 _08402_ (.A0(\median_processor.input_storage[28] ),
    .A1(net502),
    .S(net44),
    .X(_03108_));
 sg13g2_and2_1 _08403_ (.A(net484),
    .B(_03108_),
    .X(_00020_));
 sg13g2_mux2_1 _08404_ (.A0(net154),
    .A1(net500),
    .S(net44),
    .X(_03109_));
 sg13g2_and2_1 _08405_ (.A(net477),
    .B(_03109_),
    .X(_00021_));
 sg13g2_nand2_1 _08406_ (.Y(_03110_),
    .A(net151),
    .B(net51));
 sg13g2_o21ai_1 _08407_ (.B1(_03110_),
    .Y(_03111_),
    .A1(_03050_),
    .A2(net51));
 sg13g2_and2_1 _08408_ (.A(net453),
    .B(_03111_),
    .X(_00022_));
 sg13g2_nand2_1 _08409_ (.Y(_03112_),
    .A(net498),
    .B(net44));
 sg13g2_o21ai_1 _08410_ (.B1(_03112_),
    .Y(_03113_),
    .A1(_02107_),
    .A2(net44));
 sg13g2_and2_1 _08411_ (.A(net479),
    .B(_03113_),
    .X(_00023_));
 sg13g2_nand2_1 _08412_ (.Y(_03114_),
    .A(data_in_p2c_8),
    .B(net44));
 sg13g2_o21ai_1 _08413_ (.B1(_03114_),
    .Y(_03115_),
    .A1(_01759_),
    .A2(net44));
 sg13g2_and2_1 _08414_ (.A(net479),
    .B(_03115_),
    .X(_00024_));
 sg13g2_buf_1 fanout396 (.A(net397),
    .X(net396));
 sg13g2_nand2b_1 _08416_ (.Y(_03117_),
    .B(reg_addr_p2c_3),
    .A_N(reg_addr_p2c_2));
 sg13g2_nor2_1 _08417_ (.A(_03039_),
    .B(_03117_),
    .Y(_03118_));
 sg13g2_buf_2 fanout395 (.A(net397),
    .X(net395));
 sg13g2_buf_2 fanout394 (.A(net396),
    .X(net394));
 sg13g2_mux2_1 _08420_ (.A0(net145),
    .A1(data_in_p2c_1),
    .S(net42),
    .X(_03121_));
 sg13g2_and2_1 _08421_ (.A(net465),
    .B(_03121_),
    .X(_00025_));
 sg13g2_mux2_1 _08422_ (.A0(net143),
    .A1(net505),
    .S(net42),
    .X(_03122_));
 sg13g2_and2_1 _08423_ (.A(net465),
    .B(_03122_),
    .X(_00026_));
 sg13g2_nand2_1 _08424_ (.Y(_03123_),
    .A(data_in_p2c_3),
    .B(net42));
 sg13g2_o21ai_1 _08425_ (.B1(_03123_),
    .Y(_03124_),
    .A1(_01918_),
    .A2(net42));
 sg13g2_and2_1 _08426_ (.A(net466),
    .B(_03124_),
    .X(_00027_));
 sg13g2_nand2_1 _08427_ (.Y(_03125_),
    .A(data_in_p2c_4),
    .B(net42));
 sg13g2_o21ai_1 _08428_ (.B1(_03125_),
    .Y(_03126_),
    .A1(_01926_),
    .A2(net42));
 sg13g2_and2_1 _08429_ (.A(net468),
    .B(_03126_),
    .X(_00028_));
 sg13g2_nand2_1 _08430_ (.Y(_03127_),
    .A(net502),
    .B(net42));
 sg13g2_o21ai_1 _08431_ (.B1(_03127_),
    .Y(_03128_),
    .A1(_01941_),
    .A2(net42));
 sg13g2_and2_1 _08432_ (.A(net484),
    .B(_03128_),
    .X(_00029_));
 sg13g2_nand2_1 _08433_ (.Y(_03129_),
    .A(net500),
    .B(net43));
 sg13g2_o21ai_1 _08434_ (.B1(_03129_),
    .Y(_03130_),
    .A1(_02154_),
    .A2(net43));
 sg13g2_and2_1 _08435_ (.A(net477),
    .B(_03130_),
    .X(_00030_));
 sg13g2_nand2_1 _08436_ (.Y(_03131_),
    .A(net498),
    .B(net43));
 sg13g2_o21ai_1 _08437_ (.B1(_03131_),
    .Y(_03132_),
    .A1(net61),
    .A2(net43));
 sg13g2_and2_1 _08438_ (.A(net479),
    .B(_03132_),
    .X(_00031_));
 sg13g2_nand2_1 _08439_ (.Y(_03133_),
    .A(data_in_p2c_8),
    .B(net43));
 sg13g2_o21ai_1 _08440_ (.B1(_03133_),
    .Y(_03134_),
    .A1(net63),
    .A2(net43));
 sg13g2_and2_1 _08441_ (.A(net485),
    .B(_03134_),
    .X(_00032_));
 sg13g2_nand2_1 _08442_ (.Y(_03135_),
    .A(net129),
    .B(net51));
 sg13g2_o21ai_1 _08443_ (.B1(_03135_),
    .Y(_03136_),
    .A1(_03056_),
    .A2(net51));
 sg13g2_and2_1 _08444_ (.A(net452),
    .B(_03136_),
    .X(_00033_));
 sg13g2_nor2_1 _08445_ (.A(_03098_),
    .B(_03117_),
    .Y(_03137_));
 sg13g2_buf_1 fanout393 (.A(net397),
    .X(net393));
 sg13g2_buf_2 fanout392 (.A(net397),
    .X(net392));
 sg13g2_mux2_1 _08448_ (.A0(net127),
    .A1(data_in_p2c_1),
    .S(net40),
    .X(_03140_));
 sg13g2_and2_1 _08449_ (.A(net469),
    .B(_03140_),
    .X(_00034_));
 sg13g2_buf_1 fanout391 (.A(net398),
    .X(net391));
 sg13g2_nand2_1 _08451_ (.Y(_03142_),
    .A(net505),
    .B(net40));
 sg13g2_o21ai_1 _08452_ (.B1(_03142_),
    .Y(_03143_),
    .A1(net70),
    .A2(net40));
 sg13g2_and2_1 _08453_ (.A(net469),
    .B(_03143_),
    .X(_00035_));
 sg13g2_nand2_1 _08454_ (.Y(_03144_),
    .A(data_in_p2c_3),
    .B(net40));
 sg13g2_o21ai_1 _08455_ (.B1(_03144_),
    .Y(_03145_),
    .A1(_01780_),
    .A2(net40));
 sg13g2_and2_1 _08456_ (.A(net469),
    .B(_03145_),
    .X(_00036_));
 sg13g2_nand2_1 _08457_ (.Y(_03146_),
    .A(net503),
    .B(net40));
 sg13g2_o21ai_1 _08458_ (.B1(_03146_),
    .Y(_03147_),
    .A1(net69),
    .A2(net40));
 sg13g2_and2_1 _08459_ (.A(net469),
    .B(_03147_),
    .X(_00037_));
 sg13g2_nand2_1 _08460_ (.Y(_03148_),
    .A(net502),
    .B(net40));
 sg13g2_o21ai_1 _08461_ (.B1(_03148_),
    .Y(_03149_),
    .A1(_02103_),
    .A2(net41));
 sg13g2_and2_1 _08462_ (.A(net477),
    .B(_03149_),
    .X(_00038_));
 sg13g2_nand2_1 _08463_ (.Y(_03150_),
    .A(net500),
    .B(net41));
 sg13g2_o21ai_1 _08464_ (.B1(_03150_),
    .Y(_03151_),
    .A1(net68),
    .A2(net41));
 sg13g2_and2_1 _08465_ (.A(net486),
    .B(_03151_),
    .X(_00039_));
 sg13g2_nand2_1 _08466_ (.Y(_03152_),
    .A(net499),
    .B(net41));
 sg13g2_o21ai_1 _08467_ (.B1(_03152_),
    .Y(_03153_),
    .A1(_02118_),
    .A2(net41));
 sg13g2_and2_1 _08468_ (.A(net486),
    .B(_03153_),
    .X(_00040_));
 sg13g2_nand2_1 _08469_ (.Y(_03154_),
    .A(data_in_p2c_8),
    .B(net41));
 sg13g2_o21ai_1 _08470_ (.B1(_03154_),
    .Y(_03155_),
    .A1(_01765_),
    .A2(net41));
 sg13g2_and2_1 _08471_ (.A(net486),
    .B(_03155_),
    .X(_00041_));
 sg13g2_nand2_1 _08472_ (.Y(_03156_),
    .A(reg_addr_p2c_3),
    .B(reg_addr_p2c_2));
 sg13g2_nor2_1 _08473_ (.A(_03039_),
    .B(_03156_),
    .Y(_03157_));
 sg13g2_buf_1 fanout390 (.A(net391),
    .X(net390));
 sg13g2_buf_1 fanout389 (.A(net391),
    .X(net389));
 sg13g2_nand2_1 _08476_ (.Y(_03160_),
    .A(data_in_p2c_1),
    .B(net38));
 sg13g2_o21ai_1 _08477_ (.B1(_03160_),
    .Y(_03161_),
    .A1(_01884_),
    .A2(net38));
 sg13g2_and2_1 _08478_ (.A(net467),
    .B(_03161_),
    .X(_00042_));
 sg13g2_nand2_1 _08479_ (.Y(_03162_),
    .A(net505),
    .B(net38));
 sg13g2_o21ai_1 _08480_ (.B1(_03162_),
    .Y(_03163_),
    .A1(_01885_),
    .A2(net38));
 sg13g2_and2_1 _08481_ (.A(net467),
    .B(_03163_),
    .X(_00043_));
 sg13g2_mux2_1 _08482_ (.A0(net501),
    .A1(net109),
    .S(net51),
    .X(_03164_));
 sg13g2_and2_1 _08483_ (.A(net452),
    .B(_03164_),
    .X(_00044_));
 sg13g2_buf_1 fanout388 (.A(net391),
    .X(net388));
 sg13g2_nand2_1 _08485_ (.Y(_03166_),
    .A(data_in_p2c_3),
    .B(net38));
 sg13g2_o21ai_1 _08486_ (.B1(_03166_),
    .Y(_03167_),
    .A1(_01931_),
    .A2(net38));
 sg13g2_and2_1 _08487_ (.A(net466),
    .B(_03167_),
    .X(_00045_));
 sg13g2_nand2_1 _08488_ (.Y(_03168_),
    .A(data_in_p2c_4),
    .B(net38));
 sg13g2_o21ai_1 _08489_ (.B1(_03168_),
    .Y(_03169_),
    .A1(_01712_),
    .A2(net38));
 sg13g2_and2_1 _08490_ (.A(net468),
    .B(_03169_),
    .X(_00046_));
 sg13g2_nand2_1 _08491_ (.Y(_03170_),
    .A(net502),
    .B(net39));
 sg13g2_o21ai_1 _08492_ (.B1(_03170_),
    .Y(_03171_),
    .A1(_01733_),
    .A2(net39));
 sg13g2_and2_1 _08493_ (.A(net484),
    .B(_03171_),
    .X(_00047_));
 sg13g2_nand2_1 _08494_ (.Y(_03172_),
    .A(data_in_p2c_6),
    .B(net39));
 sg13g2_o21ai_1 _08495_ (.B1(_03172_),
    .Y(_03173_),
    .A1(_01730_),
    .A2(net39));
 sg13g2_and2_1 _08496_ (.A(net486),
    .B(_03173_),
    .X(_00048_));
 sg13g2_nand2_1 _08497_ (.Y(_03174_),
    .A(net499),
    .B(net39));
 sg13g2_o21ai_1 _08498_ (.B1(_03174_),
    .Y(_03175_),
    .A1(_01755_),
    .A2(net39));
 sg13g2_and2_1 _08499_ (.A(net485),
    .B(_03175_),
    .X(_00049_));
 sg13g2_nand2_1 _08500_ (.Y(_03176_),
    .A(data_in_p2c_8),
    .B(net39));
 sg13g2_o21ai_1 _08501_ (.B1(_03176_),
    .Y(_03177_),
    .A1(net73),
    .A2(net39));
 sg13g2_and2_1 _08502_ (.A(net485),
    .B(_03177_),
    .X(_00050_));
 sg13g2_or2_1 _08503_ (.X(_03178_),
    .B(_03156_),
    .A(_03098_));
 sg13g2_buf_1 fanout387 (.A(net391),
    .X(net387));
 sg13g2_buf_1 fanout386 (.A(net398),
    .X(net386));
 sg13g2_nand2_1 _08506_ (.Y(_03181_),
    .A(net96),
    .B(net36));
 sg13g2_o21ai_1 _08507_ (.B1(_03181_),
    .Y(_03182_),
    .A1(_03038_),
    .A2(net36));
 sg13g2_and2_1 _08508_ (.A(net451),
    .B(_03182_),
    .X(_00051_));
 sg13g2_mux2_1 _08509_ (.A0(net504),
    .A1(net94),
    .S(net36),
    .X(_03183_));
 sg13g2_and2_1 _08510_ (.A(net453),
    .B(_03183_),
    .X(_00052_));
 sg13g2_nand2_1 _08511_ (.Y(_03184_),
    .A(net92),
    .B(net36));
 sg13g2_o21ai_1 _08512_ (.B1(_03184_),
    .Y(_03185_),
    .A1(_03050_),
    .A2(net36));
 sg13g2_and2_1 _08513_ (.A(net453),
    .B(_03185_),
    .X(_00053_));
 sg13g2_nor2_1 _08514_ (.A(_03056_),
    .B(net36),
    .Y(_03186_));
 sg13g2_a21oi_1 _08515_ (.A1(net91),
    .A2(net36),
    .Y(_03187_),
    .B1(_03186_));
 sg13g2_nor2b_1 _08516_ (.A(_03187_),
    .B_N(net452),
    .Y(_00054_));
 sg13g2_nand2_1 _08517_ (.Y(_03188_),
    .A(net89),
    .B(net52));
 sg13g2_o21ai_1 _08518_ (.B1(_03188_),
    .Y(_03189_),
    .A1(_03063_),
    .A2(net52));
 sg13g2_and2_1 _08519_ (.A(net476),
    .B(_03189_),
    .X(_00055_));
 sg13g2_buf_2 fanout385 (.A(net386),
    .X(net385));
 sg13g2_mux2_1 _08521_ (.A0(net501),
    .A1(net87),
    .S(net36),
    .X(_03191_));
 sg13g2_and2_1 _08522_ (.A(net476),
    .B(_03191_),
    .X(_00056_));
 sg13g2_nand2_1 _08523_ (.Y(_03192_),
    .A(net86),
    .B(net37));
 sg13g2_o21ai_1 _08524_ (.B1(_03192_),
    .Y(_03193_),
    .A1(_03063_),
    .A2(net37));
 sg13g2_and2_1 _08525_ (.A(net476),
    .B(_03193_),
    .X(_00057_));
 sg13g2_nand2_1 _08526_ (.Y(_03194_),
    .A(net84),
    .B(net37));
 sg13g2_o21ai_1 _08527_ (.B1(_03194_),
    .Y(_03195_),
    .A1(_03067_),
    .A2(net37));
 sg13g2_and2_1 _08528_ (.A(net478),
    .B(_03195_),
    .X(_00058_));
 sg13g2_nand2_1 _08529_ (.Y(_03196_),
    .A(net83),
    .B(net37));
 sg13g2_o21ai_1 _08530_ (.B1(_03196_),
    .Y(_03197_),
    .A1(_03071_),
    .A2(net37));
 sg13g2_and2_1 _08531_ (.A(net479),
    .B(_03197_),
    .X(_00059_));
 sg13g2_nand2_1 _08532_ (.Y(_03198_),
    .A(net81),
    .B(net52));
 sg13g2_o21ai_1 _08533_ (.B1(_03198_),
    .Y(_03199_),
    .A1(_03067_),
    .A2(net52));
 sg13g2_and2_1 _08534_ (.A(net478),
    .B(_03199_),
    .X(_00060_));
 sg13g2_nand2_1 _08535_ (.Y(_03200_),
    .A(net79),
    .B(net52));
 sg13g2_o21ai_1 _08536_ (.B1(_03200_),
    .Y(_03201_),
    .A1(_03071_),
    .A2(net52));
 sg13g2_and2_1 _08537_ (.A(net479),
    .B(_03201_),
    .X(_00061_));
 sg13g2_nor2_1 _08538_ (.A(_03038_),
    .B(net49),
    .Y(_03202_));
 sg13g2_a21oi_1 _08539_ (.A1(net75),
    .A2(net49),
    .Y(_03203_),
    .B1(_03202_));
 sg13g2_nor2b_1 _08540_ (.A(_03203_),
    .B_N(net453),
    .Y(_00062_));
 sg13g2_mux2_1 _08541_ (.A0(net504),
    .A1(net74),
    .S(net49),
    .X(_03204_));
 sg13g2_and2_1 _08542_ (.A(net451),
    .B(_03204_),
    .X(_00063_));
 sg13g2_buf_2 fanout384 (.A(net385),
    .X(net384));
 sg13g2_buf_2 fanout383 (.A(net386),
    .X(net383));
 sg13g2_and2_1 _08545_ (.A(net314),
    .B(net613),
    .X(_03207_));
 sg13g2_buf_2 fanout382 (.A(net386),
    .X(net382));
 sg13g2_buf_1 fanout381 (.A(net398),
    .X(net381));
 sg13g2_xnor2_1 _08548_ (.Y(_03210_),
    .A(\rando_generator.lfsr_reg[27] ),
    .B(\rando_generator.lfsr_reg[30] ));
 sg13g2_and2_1 _08549_ (.A(net199),
    .B(_03210_),
    .X(_00072_));
 sg13g2_and2_1 _08550_ (.A(\rando_generator.lfsr_reg[9] ),
    .B(net200),
    .X(_00073_));
 sg13g2_and2_1 _08551_ (.A(\rando_generator.lfsr_reg[10] ),
    .B(net200),
    .X(_00074_));
 sg13g2_and2_1 _08552_ (.A(\rando_generator.lfsr_reg[11] ),
    .B(net201),
    .X(_00075_));
 sg13g2_and2_1 _08553_ (.A(\rando_generator.lfsr_reg[12] ),
    .B(net201),
    .X(_00076_));
 sg13g2_and2_1 _08554_ (.A(\rando_generator.lfsr_reg[13] ),
    .B(net203),
    .X(_00077_));
 sg13g2_and2_1 _08555_ (.A(\rando_generator.lfsr_reg[14] ),
    .B(net201),
    .X(_00078_));
 sg13g2_and2_1 _08556_ (.A(\rando_generator.lfsr_reg[15] ),
    .B(net201),
    .X(_00079_));
 sg13g2_and2_1 _08557_ (.A(\rando_generator.lfsr_reg[16] ),
    .B(net201),
    .X(_00080_));
 sg13g2_and2_1 _08558_ (.A(\rando_generator.lfsr_reg[17] ),
    .B(net201),
    .X(_00081_));
 sg13g2_buf_2 fanout380 (.A(net381),
    .X(net380));
 sg13g2_and2_1 _08560_ (.A(\rando_generator.lfsr_reg[18] ),
    .B(net201),
    .X(_00082_));
 sg13g2_and2_1 _08561_ (.A(lfsr_out_c2p),
    .B(net199),
    .X(_00083_));
 sg13g2_and2_1 _08562_ (.A(\rando_generator.lfsr_reg[19] ),
    .B(net202),
    .X(_00084_));
 sg13g2_and2_1 _08563_ (.A(\rando_generator.lfsr_reg[20] ),
    .B(net202),
    .X(_00085_));
 sg13g2_and2_1 _08564_ (.A(\rando_generator.lfsr_reg[21] ),
    .B(net202),
    .X(_00086_));
 sg13g2_and2_1 _08565_ (.A(\rando_generator.lfsr_reg[22] ),
    .B(net202),
    .X(_00087_));
 sg13g2_and2_1 _08566_ (.A(\rando_generator.lfsr_reg[23] ),
    .B(net202),
    .X(_00088_));
 sg13g2_and2_1 _08567_ (.A(\rando_generator.lfsr_reg[24] ),
    .B(net202),
    .X(_00089_));
 sg13g2_and2_1 _08568_ (.A(\rando_generator.lfsr_reg[25] ),
    .B(net203),
    .X(_00090_));
 sg13g2_and2_1 _08569_ (.A(\rando_generator.lfsr_reg[26] ),
    .B(net202),
    .X(_00091_));
 sg13g2_buf_1 fanout379 (.A(net380),
    .X(net379));
 sg13g2_and2_1 _08571_ (.A(\rando_generator.lfsr_reg[27] ),
    .B(net200),
    .X(_00092_));
 sg13g2_and2_1 _08572_ (.A(\rando_generator.lfsr_reg[28] ),
    .B(net199),
    .X(_00093_));
 sg13g2_and2_1 _08573_ (.A(\rando_generator.lfsr_reg[1] ),
    .B(net199),
    .X(_00094_));
 sg13g2_and2_1 _08574_ (.A(\rando_generator.lfsr_reg[29] ),
    .B(net199),
    .X(_00095_));
 sg13g2_and2_1 _08575_ (.A(\rando_generator.lfsr_reg[2] ),
    .B(net199),
    .X(_00096_));
 sg13g2_and2_1 _08576_ (.A(\rando_generator.lfsr_reg[3] ),
    .B(net199),
    .X(_00097_));
 sg13g2_and2_1 _08577_ (.A(\rando_generator.lfsr_reg[4] ),
    .B(net199),
    .X(_00098_));
 sg13g2_and2_1 _08578_ (.A(\rando_generator.lfsr_reg[5] ),
    .B(net200),
    .X(_00099_));
 sg13g2_and2_1 _08579_ (.A(\rando_generator.lfsr_reg[6] ),
    .B(net200),
    .X(_00100_));
 sg13g2_and2_1 _08580_ (.A(\rando_generator.lfsr_reg[7] ),
    .B(net202),
    .X(_00101_));
 sg13g2_and2_1 _08581_ (.A(\rando_generator.lfsr_reg[8] ),
    .B(net201),
    .X(_00102_));
 sg13g2_buf_1 fanout378 (.A(net381),
    .X(net378));
 sg13g2_buf_2 fanout377 (.A(net378),
    .X(net377));
 sg13g2_mux2_1 _08584_ (.A0(\shift_storage.storage[0] ),
    .A1(\shift_storage.shreg_in ),
    .S(net613),
    .X(_03215_));
 sg13g2_and2_1 _08585_ (.A(net315),
    .B(_03215_),
    .X(_00103_));
 sg13g2_mux2_1 _08586_ (.A0(\shift_storage.storage[1000] ),
    .A1(\shift_storage.storage[999] ),
    .S(net709),
    .X(_03216_));
 sg13g2_and2_1 _08587_ (.A(net415),
    .B(_03216_),
    .X(_00104_));
 sg13g2_mux2_1 _08588_ (.A0(\shift_storage.storage[1001] ),
    .A1(\shift_storage.storage[1000] ),
    .S(net723),
    .X(_03217_));
 sg13g2_and2_1 _08589_ (.A(net429),
    .B(_03217_),
    .X(_00105_));
 sg13g2_buf_1 fanout376 (.A(net493),
    .X(net376));
 sg13g2_buf_1 fanout375 (.A(net376),
    .X(net375));
 sg13g2_mux2_1 _08592_ (.A0(\shift_storage.storage[1002] ),
    .A1(\shift_storage.storage[1001] ),
    .S(net723),
    .X(_03220_));
 sg13g2_and2_1 _08593_ (.A(net429),
    .B(_03220_),
    .X(_00106_));
 sg13g2_mux2_1 _08594_ (.A0(\shift_storage.storage[1003] ),
    .A1(\shift_storage.storage[1002] ),
    .S(net723),
    .X(_03221_));
 sg13g2_and2_1 _08595_ (.A(net429),
    .B(_03221_),
    .X(_00107_));
 sg13g2_mux2_1 _08596_ (.A0(\shift_storage.storage[1004] ),
    .A1(\shift_storage.storage[1003] ),
    .S(net724),
    .X(_03222_));
 sg13g2_and2_1 _08597_ (.A(net429),
    .B(_03222_),
    .X(_00108_));
 sg13g2_mux2_1 _08598_ (.A0(\shift_storage.storage[1005] ),
    .A1(\shift_storage.storage[1004] ),
    .S(net723),
    .X(_03223_));
 sg13g2_and2_1 _08599_ (.A(net429),
    .B(_03223_),
    .X(_00109_));
 sg13g2_mux2_1 _08600_ (.A0(\shift_storage.storage[1006] ),
    .A1(\shift_storage.storage[1005] ),
    .S(net723),
    .X(_03224_));
 sg13g2_and2_1 _08601_ (.A(net429),
    .B(_03224_),
    .X(_00110_));
 sg13g2_mux2_1 _08602_ (.A0(\shift_storage.storage[1007] ),
    .A1(\shift_storage.storage[1006] ),
    .S(net723),
    .X(_03225_));
 sg13g2_and2_1 _08603_ (.A(net422),
    .B(_03225_),
    .X(_00111_));
 sg13g2_mux2_1 _08604_ (.A0(\shift_storage.storage[1008] ),
    .A1(\shift_storage.storage[1007] ),
    .S(net716),
    .X(_03226_));
 sg13g2_and2_1 _08605_ (.A(net422),
    .B(_03226_),
    .X(_00112_));
 sg13g2_buf_1 fanout374 (.A(net375),
    .X(net374));
 sg13g2_mux2_1 _08607_ (.A0(\shift_storage.storage[1009] ),
    .A1(\shift_storage.storage[1008] ),
    .S(net717),
    .X(_03228_));
 sg13g2_and2_1 _08608_ (.A(net423),
    .B(_03228_),
    .X(_00113_));
 sg13g2_mux2_1 _08609_ (.A0(\shift_storage.storage[100] ),
    .A1(\shift_storage.storage[99] ),
    .S(net620),
    .X(_03229_));
 sg13g2_and2_1 _08610_ (.A(net322),
    .B(_03229_),
    .X(_00114_));
 sg13g2_mux2_1 _08611_ (.A0(\shift_storage.storage[1010] ),
    .A1(\shift_storage.storage[1009] ),
    .S(net717),
    .X(_03230_));
 sg13g2_and2_1 _08612_ (.A(net423),
    .B(_03230_),
    .X(_00115_));
 sg13g2_buf_2 fanout373 (.A(net375),
    .X(net373));
 sg13g2_mux2_1 _08614_ (.A0(\shift_storage.storage[1011] ),
    .A1(\shift_storage.storage[1010] ),
    .S(net717),
    .X(_03232_));
 sg13g2_and2_1 _08615_ (.A(net423),
    .B(_03232_),
    .X(_00116_));
 sg13g2_mux2_1 _08616_ (.A0(\shift_storage.storage[1012] ),
    .A1(\shift_storage.storage[1011] ),
    .S(net717),
    .X(_03233_));
 sg13g2_and2_1 _08617_ (.A(net423),
    .B(_03233_),
    .X(_00117_));
 sg13g2_mux2_1 _08618_ (.A0(\shift_storage.storage[1013] ),
    .A1(\shift_storage.storage[1012] ),
    .S(net717),
    .X(_03234_));
 sg13g2_and2_1 _08619_ (.A(net423),
    .B(_03234_),
    .X(_00118_));
 sg13g2_mux2_1 _08620_ (.A0(\shift_storage.storage[1014] ),
    .A1(\shift_storage.storage[1013] ),
    .S(net717),
    .X(_03235_));
 sg13g2_and2_1 _08621_ (.A(net428),
    .B(_03235_),
    .X(_00119_));
 sg13g2_mux2_1 _08622_ (.A0(\shift_storage.storage[1015] ),
    .A1(\shift_storage.storage[1014] ),
    .S(net716),
    .X(_03236_));
 sg13g2_and2_1 _08623_ (.A(net422),
    .B(_03236_),
    .X(_00120_));
 sg13g2_mux2_1 _08624_ (.A0(\shift_storage.storage[1016] ),
    .A1(\shift_storage.storage[1015] ),
    .S(net716),
    .X(_03237_));
 sg13g2_and2_1 _08625_ (.A(net422),
    .B(_03237_),
    .X(_00121_));
 sg13g2_mux2_1 _08626_ (.A0(\shift_storage.storage[1017] ),
    .A1(\shift_storage.storage[1016] ),
    .S(net716),
    .X(_03238_));
 sg13g2_and2_1 _08627_ (.A(net422),
    .B(_03238_),
    .X(_00122_));
 sg13g2_buf_2 fanout372 (.A(net375),
    .X(net372));
 sg13g2_mux2_1 _08629_ (.A0(\shift_storage.storage[1018] ),
    .A1(\shift_storage.storage[1017] ),
    .S(net716),
    .X(_03240_));
 sg13g2_and2_1 _08630_ (.A(net422),
    .B(_03240_),
    .X(_00123_));
 sg13g2_mux2_1 _08631_ (.A0(\shift_storage.storage[1019] ),
    .A1(\shift_storage.storage[1018] ),
    .S(net716),
    .X(_03241_));
 sg13g2_and2_1 _08632_ (.A(net422),
    .B(_03241_),
    .X(_00124_));
 sg13g2_mux2_1 _08633_ (.A0(\shift_storage.storage[101] ),
    .A1(\shift_storage.storage[100] ),
    .S(net619),
    .X(_03242_));
 sg13g2_and2_1 _08634_ (.A(net322),
    .B(_03242_),
    .X(_00125_));
 sg13g2_buf_2 fanout371 (.A(net372),
    .X(net371));
 sg13g2_mux2_1 _08636_ (.A0(\shift_storage.storage[1020] ),
    .A1(\shift_storage.storage[1019] ),
    .S(net715),
    .X(_03244_));
 sg13g2_and2_1 _08637_ (.A(net421),
    .B(_03244_),
    .X(_00126_));
 sg13g2_mux2_1 _08638_ (.A0(\shift_storage.storage[1021] ),
    .A1(\shift_storage.storage[1020] ),
    .S(net697),
    .X(_03245_));
 sg13g2_and2_1 _08639_ (.A(net402),
    .B(_03245_),
    .X(_00127_));
 sg13g2_mux2_1 _08640_ (.A0(\shift_storage.storage[1022] ),
    .A1(\shift_storage.storage[1021] ),
    .S(net697),
    .X(_03246_));
 sg13g2_and2_1 _08641_ (.A(net402),
    .B(_03246_),
    .X(_00128_));
 sg13g2_mux2_1 _08642_ (.A0(\shift_storage.storage[1023] ),
    .A1(\shift_storage.storage[1022] ),
    .S(net700),
    .X(_03247_));
 sg13g2_and2_1 _08643_ (.A(net405),
    .B(_03247_),
    .X(_00129_));
 sg13g2_mux2_1 _08644_ (.A0(\shift_storage.storage[1024] ),
    .A1(\shift_storage.storage[1023] ),
    .S(net700),
    .X(_03248_));
 sg13g2_and2_1 _08645_ (.A(net405),
    .B(_03248_),
    .X(_00130_));
 sg13g2_mux2_1 _08646_ (.A0(\shift_storage.storage[1025] ),
    .A1(\shift_storage.storage[1024] ),
    .S(net697),
    .X(_03249_));
 sg13g2_and2_1 _08647_ (.A(net402),
    .B(_03249_),
    .X(_00131_));
 sg13g2_mux2_1 _08648_ (.A0(\shift_storage.storage[1026] ),
    .A1(\shift_storage.storage[1025] ),
    .S(net669),
    .X(_03250_));
 sg13g2_and2_1 _08649_ (.A(net374),
    .B(_03250_),
    .X(_00132_));
 sg13g2_buf_2 fanout370 (.A(net376),
    .X(net370));
 sg13g2_mux2_1 _08651_ (.A0(\shift_storage.storage[1027] ),
    .A1(\shift_storage.storage[1026] ),
    .S(net670),
    .X(_03252_));
 sg13g2_and2_1 _08652_ (.A(net374),
    .B(_03252_),
    .X(_00133_));
 sg13g2_mux2_1 _08653_ (.A0(\shift_storage.storage[1028] ),
    .A1(\shift_storage.storage[1027] ),
    .S(net670),
    .X(_03253_));
 sg13g2_and2_1 _08654_ (.A(net374),
    .B(_03253_),
    .X(_00134_));
 sg13g2_mux2_1 _08655_ (.A0(\shift_storage.storage[1029] ),
    .A1(\shift_storage.storage[1028] ),
    .S(net670),
    .X(_03254_));
 sg13g2_and2_1 _08656_ (.A(net373),
    .B(_03254_),
    .X(_00135_));
 sg13g2_buf_2 fanout369 (.A(net370),
    .X(net369));
 sg13g2_mux2_1 _08658_ (.A0(\shift_storage.storage[102] ),
    .A1(\shift_storage.storage[101] ),
    .S(net619),
    .X(_03256_));
 sg13g2_and2_1 _08659_ (.A(net321),
    .B(_03256_),
    .X(_00136_));
 sg13g2_mux2_1 _08660_ (.A0(\shift_storage.storage[1030] ),
    .A1(\shift_storage.storage[1029] ),
    .S(net670),
    .X(_03257_));
 sg13g2_and2_1 _08661_ (.A(net374),
    .B(_03257_),
    .X(_00137_));
 sg13g2_mux2_1 _08662_ (.A0(\shift_storage.storage[1031] ),
    .A1(\shift_storage.storage[1030] ),
    .S(net670),
    .X(_03258_));
 sg13g2_and2_1 _08663_ (.A(net372),
    .B(_03258_),
    .X(_00138_));
 sg13g2_mux2_1 _08664_ (.A0(\shift_storage.storage[1032] ),
    .A1(\shift_storage.storage[1031] ),
    .S(net668),
    .X(_03259_));
 sg13g2_and2_1 _08665_ (.A(net375),
    .B(_03259_),
    .X(_00139_));
 sg13g2_mux2_1 _08666_ (.A0(\shift_storage.storage[1033] ),
    .A1(\shift_storage.storage[1032] ),
    .S(net669),
    .X(_03260_));
 sg13g2_and2_1 _08667_ (.A(net373),
    .B(_03260_),
    .X(_00140_));
 sg13g2_mux2_1 _08668_ (.A0(\shift_storage.storage[1034] ),
    .A1(\shift_storage.storage[1033] ),
    .S(net670),
    .X(_03261_));
 sg13g2_and2_1 _08669_ (.A(net389),
    .B(_03261_),
    .X(_00141_));
 sg13g2_mux2_1 _08670_ (.A0(\shift_storage.storage[1035] ),
    .A1(\shift_storage.storage[1034] ),
    .S(net684),
    .X(_03262_));
 sg13g2_and2_1 _08671_ (.A(net389),
    .B(_03262_),
    .X(_00142_));
 sg13g2_buf_1 fanout368 (.A(net376),
    .X(net368));
 sg13g2_mux2_1 _08673_ (.A0(\shift_storage.storage[1036] ),
    .A1(\shift_storage.storage[1035] ),
    .S(net684),
    .X(_03264_));
 sg13g2_and2_1 _08674_ (.A(net389),
    .B(_03264_),
    .X(_00143_));
 sg13g2_mux2_1 _08675_ (.A0(\shift_storage.storage[1037] ),
    .A1(\shift_storage.storage[1036] ),
    .S(net684),
    .X(_03265_));
 sg13g2_and2_1 _08676_ (.A(net389),
    .B(_03265_),
    .X(_00144_));
 sg13g2_mux2_1 _08677_ (.A0(\shift_storage.storage[1038] ),
    .A1(\shift_storage.storage[1037] ),
    .S(net684),
    .X(_03266_));
 sg13g2_and2_1 _08678_ (.A(net389),
    .B(_03266_),
    .X(_00145_));
 sg13g2_buf_2 fanout367 (.A(net368),
    .X(net367));
 sg13g2_mux2_1 _08680_ (.A0(\shift_storage.storage[1039] ),
    .A1(\shift_storage.storage[1038] ),
    .S(net684),
    .X(_03268_));
 sg13g2_and2_1 _08681_ (.A(net419),
    .B(_03268_),
    .X(_00146_));
 sg13g2_mux2_1 _08682_ (.A0(\shift_storage.storage[103] ),
    .A1(\shift_storage.storage[102] ),
    .S(net622),
    .X(_03269_));
 sg13g2_and2_1 _08683_ (.A(net323),
    .B(_03269_),
    .X(_00147_));
 sg13g2_mux2_1 _08684_ (.A0(\shift_storage.storage[1040] ),
    .A1(\shift_storage.storage[1039] ),
    .S(net713),
    .X(_03270_));
 sg13g2_and2_1 _08685_ (.A(net419),
    .B(_03270_),
    .X(_00148_));
 sg13g2_mux2_1 _08686_ (.A0(\shift_storage.storage[1041] ),
    .A1(\shift_storage.storage[1040] ),
    .S(net713),
    .X(_03271_));
 sg13g2_and2_1 _08687_ (.A(net419),
    .B(_03271_),
    .X(_00149_));
 sg13g2_mux2_1 _08688_ (.A0(\shift_storage.storage[1042] ),
    .A1(\shift_storage.storage[1041] ),
    .S(net713),
    .X(_03272_));
 sg13g2_and2_1 _08689_ (.A(net419),
    .B(_03272_),
    .X(_00150_));
 sg13g2_mux2_1 _08690_ (.A0(\shift_storage.storage[1043] ),
    .A1(\shift_storage.storage[1042] ),
    .S(net713),
    .X(_03273_));
 sg13g2_and2_1 _08691_ (.A(net421),
    .B(_03273_),
    .X(_00151_));
 sg13g2_mux2_1 _08692_ (.A0(\shift_storage.storage[1044] ),
    .A1(\shift_storage.storage[1043] ),
    .S(net713),
    .X(_03274_));
 sg13g2_and2_1 _08693_ (.A(net421),
    .B(_03274_),
    .X(_00152_));
 sg13g2_buf_1 fanout366 (.A(net376),
    .X(net366));
 sg13g2_mux2_1 _08695_ (.A0(\shift_storage.storage[1045] ),
    .A1(\shift_storage.storage[1044] ),
    .S(net715),
    .X(_03276_));
 sg13g2_and2_1 _08696_ (.A(net419),
    .B(_03276_),
    .X(_00153_));
 sg13g2_mux2_1 _08697_ (.A0(\shift_storage.storage[1046] ),
    .A1(\shift_storage.storage[1045] ),
    .S(net713),
    .X(_03277_));
 sg13g2_and2_1 _08698_ (.A(net419),
    .B(_03277_),
    .X(_00154_));
 sg13g2_mux2_1 _08699_ (.A0(\shift_storage.storage[1047] ),
    .A1(\shift_storage.storage[1046] ),
    .S(net715),
    .X(_03278_));
 sg13g2_and2_1 _08700_ (.A(net420),
    .B(_03278_),
    .X(_00155_));
 sg13g2_buf_1 fanout365 (.A(net366),
    .X(net365));
 sg13g2_mux2_1 _08702_ (.A0(\shift_storage.storage[1048] ),
    .A1(\shift_storage.storage[1047] ),
    .S(net714),
    .X(_03280_));
 sg13g2_and2_1 _08703_ (.A(net421),
    .B(_03280_),
    .X(_00156_));
 sg13g2_mux2_1 _08704_ (.A0(\shift_storage.storage[1049] ),
    .A1(\shift_storage.storage[1048] ),
    .S(net714),
    .X(_03281_));
 sg13g2_and2_1 _08705_ (.A(net421),
    .B(_03281_),
    .X(_00157_));
 sg13g2_mux2_1 _08706_ (.A0(\shift_storage.storage[104] ),
    .A1(\shift_storage.storage[103] ),
    .S(net622),
    .X(_03282_));
 sg13g2_and2_1 _08707_ (.A(net323),
    .B(_03282_),
    .X(_00158_));
 sg13g2_mux2_1 _08708_ (.A0(\shift_storage.storage[1050] ),
    .A1(\shift_storage.storage[1049] ),
    .S(net714),
    .X(_03283_));
 sg13g2_and2_1 _08709_ (.A(net420),
    .B(_03283_),
    .X(_00159_));
 sg13g2_mux2_1 _08710_ (.A0(\shift_storage.storage[1051] ),
    .A1(\shift_storage.storage[1050] ),
    .S(net715),
    .X(_03284_));
 sg13g2_and2_1 _08711_ (.A(net421),
    .B(_03284_),
    .X(_00160_));
 sg13g2_mux2_1 _08712_ (.A0(\shift_storage.storage[1052] ),
    .A1(\shift_storage.storage[1051] ),
    .S(net718),
    .X(_03285_));
 sg13g2_and2_1 _08713_ (.A(net424),
    .B(_03285_),
    .X(_00161_));
 sg13g2_mux2_1 _08714_ (.A0(\shift_storage.storage[1053] ),
    .A1(\shift_storage.storage[1052] ),
    .S(net718),
    .X(_03286_));
 sg13g2_and2_1 _08715_ (.A(net424),
    .B(_03286_),
    .X(_00162_));
 sg13g2_buf_2 fanout364 (.A(net366),
    .X(net364));
 sg13g2_mux2_1 _08717_ (.A0(\shift_storage.storage[1054] ),
    .A1(\shift_storage.storage[1053] ),
    .S(net720),
    .X(_03288_));
 sg13g2_and2_1 _08718_ (.A(net426),
    .B(_03288_),
    .X(_00163_));
 sg13g2_mux2_1 _08719_ (.A0(\shift_storage.storage[1055] ),
    .A1(\shift_storage.storage[1054] ),
    .S(net720),
    .X(_03289_));
 sg13g2_and2_1 _08720_ (.A(net426),
    .B(_03289_),
    .X(_00164_));
 sg13g2_mux2_1 _08721_ (.A0(\shift_storage.storage[1056] ),
    .A1(\shift_storage.storage[1055] ),
    .S(net720),
    .X(_03290_));
 sg13g2_and2_1 _08722_ (.A(net426),
    .B(_03290_),
    .X(_00165_));
 sg13g2_buf_1 fanout363 (.A(net366),
    .X(net363));
 sg13g2_mux2_1 _08724_ (.A0(\shift_storage.storage[1057] ),
    .A1(\shift_storage.storage[1056] ),
    .S(net720),
    .X(_03292_));
 sg13g2_and2_1 _08725_ (.A(net426),
    .B(_03292_),
    .X(_00166_));
 sg13g2_mux2_1 _08726_ (.A0(\shift_storage.storage[1058] ),
    .A1(\shift_storage.storage[1057] ),
    .S(net720),
    .X(_03293_));
 sg13g2_and2_1 _08727_ (.A(net426),
    .B(_03293_),
    .X(_00167_));
 sg13g2_mux2_1 _08728_ (.A0(\shift_storage.storage[1059] ),
    .A1(\shift_storage.storage[1058] ),
    .S(net720),
    .X(_03294_));
 sg13g2_and2_1 _08729_ (.A(net433),
    .B(_03294_),
    .X(_00168_));
 sg13g2_mux2_1 _08730_ (.A0(\shift_storage.storage[105] ),
    .A1(\shift_storage.storage[104] ),
    .S(net622),
    .X(_03295_));
 sg13g2_and2_1 _08731_ (.A(net322),
    .B(_03295_),
    .X(_00169_));
 sg13g2_mux2_1 _08732_ (.A0(\shift_storage.storage[1060] ),
    .A1(\shift_storage.storage[1059] ),
    .S(net717),
    .X(_03296_));
 sg13g2_and2_1 _08733_ (.A(net423),
    .B(_03296_),
    .X(_00170_));
 sg13g2_mux2_1 _08734_ (.A0(\shift_storage.storage[1061] ),
    .A1(\shift_storage.storage[1060] ),
    .S(net724),
    .X(_03297_));
 sg13g2_and2_1 _08735_ (.A(net430),
    .B(_03297_),
    .X(_00171_));
 sg13g2_mux2_1 _08736_ (.A0(\shift_storage.storage[1062] ),
    .A1(\shift_storage.storage[1061] ),
    .S(net724),
    .X(_03298_));
 sg13g2_and2_1 _08737_ (.A(net430),
    .B(_03298_),
    .X(_00172_));
 sg13g2_buf_2 fanout362 (.A(net366),
    .X(net362));
 sg13g2_buf_1 fanout361 (.A(net362),
    .X(net361));
 sg13g2_buf_1 fanout360 (.A(net376),
    .X(net360));
 sg13g2_mux2_1 _08741_ (.A0(\shift_storage.storage[1063] ),
    .A1(\shift_storage.storage[1062] ),
    .S(net724),
    .X(_03302_));
 sg13g2_and2_1 _08742_ (.A(net430),
    .B(_03302_),
    .X(_00173_));
 sg13g2_mux2_1 _08743_ (.A0(\shift_storage.storage[1064] ),
    .A1(\shift_storage.storage[1063] ),
    .S(net724),
    .X(_03303_));
 sg13g2_and2_1 _08744_ (.A(net430),
    .B(_03303_),
    .X(_00174_));
 sg13g2_mux2_1 _08745_ (.A0(\shift_storage.storage[1065] ),
    .A1(\shift_storage.storage[1064] ),
    .S(net727),
    .X(_03304_));
 sg13g2_and2_1 _08746_ (.A(net433),
    .B(_03304_),
    .X(_00175_));
 sg13g2_buf_2 fanout359 (.A(net360),
    .X(net359));
 sg13g2_buf_1 fanout358 (.A(net360),
    .X(net358));
 sg13g2_buf_2 fanout357 (.A(net360),
    .X(net357));
 sg13g2_mux2_1 _08750_ (.A0(\shift_storage.storage[1066] ),
    .A1(\shift_storage.storage[1065] ),
    .S(net727),
    .X(_03308_));
 sg13g2_and2_1 _08751_ (.A(net433),
    .B(_03308_),
    .X(_00176_));
 sg13g2_mux2_1 _08752_ (.A0(\shift_storage.storage[1067] ),
    .A1(\shift_storage.storage[1066] ),
    .S(net727),
    .X(_03309_));
 sg13g2_and2_1 _08753_ (.A(net433),
    .B(_03309_),
    .X(_00177_));
 sg13g2_mux2_1 _08754_ (.A0(\shift_storage.storage[1068] ),
    .A1(\shift_storage.storage[1067] ),
    .S(net727),
    .X(_03310_));
 sg13g2_and2_1 _08755_ (.A(net433),
    .B(_03310_),
    .X(_00178_));
 sg13g2_mux2_1 _08756_ (.A0(\shift_storage.storage[1069] ),
    .A1(\shift_storage.storage[1068] ),
    .S(net727),
    .X(_03311_));
 sg13g2_and2_1 _08757_ (.A(net433),
    .B(_03311_),
    .X(_00179_));
 sg13g2_mux2_1 _08758_ (.A0(\shift_storage.storage[106] ),
    .A1(\shift_storage.storage[105] ),
    .S(net619),
    .X(_03312_));
 sg13g2_and2_1 _08759_ (.A(net321),
    .B(_03312_),
    .X(_00180_));
 sg13g2_mux2_1 _08760_ (.A0(\shift_storage.storage[1070] ),
    .A1(\shift_storage.storage[1069] ),
    .S(net727),
    .X(_03313_));
 sg13g2_and2_1 _08761_ (.A(net433),
    .B(_03313_),
    .X(_00181_));
 sg13g2_mux2_1 _08762_ (.A0(\shift_storage.storage[1071] ),
    .A1(\shift_storage.storage[1070] ),
    .S(net727),
    .X(_03314_));
 sg13g2_and2_1 _08763_ (.A(net434),
    .B(_03314_),
    .X(_00182_));
 sg13g2_buf_1 fanout356 (.A(\median_processor.rst ),
    .X(net356));
 sg13g2_mux2_1 _08765_ (.A0(\shift_storage.storage[1072] ),
    .A1(\shift_storage.storage[1071] ),
    .S(net720),
    .X(_03316_));
 sg13g2_and2_1 _08766_ (.A(net426),
    .B(_03316_),
    .X(_00183_));
 sg13g2_mux2_1 _08767_ (.A0(\shift_storage.storage[1073] ),
    .A1(\shift_storage.storage[1072] ),
    .S(net720),
    .X(_03317_));
 sg13g2_and2_1 _08768_ (.A(net426),
    .B(_03317_),
    .X(_00184_));
 sg13g2_mux2_1 _08769_ (.A0(\shift_storage.storage[1074] ),
    .A1(\shift_storage.storage[1073] ),
    .S(net721),
    .X(_03318_));
 sg13g2_and2_1 _08770_ (.A(net427),
    .B(_03318_),
    .X(_00185_));
 sg13g2_buf_1 fanout355 (.A(net356),
    .X(net355));
 sg13g2_mux2_1 _08772_ (.A0(\shift_storage.storage[1075] ),
    .A1(\shift_storage.storage[1074] ),
    .S(net721),
    .X(_03320_));
 sg13g2_and2_1 _08773_ (.A(net426),
    .B(_03320_),
    .X(_00186_));
 sg13g2_mux2_1 _08774_ (.A0(\shift_storage.storage[1076] ),
    .A1(\shift_storage.storage[1075] ),
    .S(net721),
    .X(_03321_));
 sg13g2_and2_1 _08775_ (.A(net425),
    .B(_03321_),
    .X(_00187_));
 sg13g2_mux2_1 _08776_ (.A0(\shift_storage.storage[1077] ),
    .A1(\shift_storage.storage[1076] ),
    .S(net719),
    .X(_03322_));
 sg13g2_and2_1 _08777_ (.A(net425),
    .B(_03322_),
    .X(_00188_));
 sg13g2_mux2_1 _08778_ (.A0(\shift_storage.storage[1078] ),
    .A1(\shift_storage.storage[1077] ),
    .S(net719),
    .X(_03323_));
 sg13g2_and2_1 _08779_ (.A(net425),
    .B(_03323_),
    .X(_00189_));
 sg13g2_mux2_1 _08780_ (.A0(\shift_storage.storage[1079] ),
    .A1(\shift_storage.storage[1078] ),
    .S(net719),
    .X(_03324_));
 sg13g2_and2_1 _08781_ (.A(net425),
    .B(_03324_),
    .X(_00190_));
 sg13g2_mux2_1 _08782_ (.A0(\shift_storage.storage[107] ),
    .A1(\shift_storage.storage[106] ),
    .S(net573),
    .X(_03325_));
 sg13g2_and2_1 _08783_ (.A(net272),
    .B(_03325_),
    .X(_00191_));
 sg13g2_mux2_1 _08784_ (.A0(\shift_storage.storage[1080] ),
    .A1(\shift_storage.storage[1079] ),
    .S(net718),
    .X(_03326_));
 sg13g2_and2_1 _08785_ (.A(net424),
    .B(_03326_),
    .X(_00192_));
 sg13g2_buf_2 fanout354 (.A(net355),
    .X(net354));
 sg13g2_mux2_1 _08787_ (.A0(\shift_storage.storage[1081] ),
    .A1(\shift_storage.storage[1080] ),
    .S(net718),
    .X(_03328_));
 sg13g2_and2_1 _08788_ (.A(net424),
    .B(_03328_),
    .X(_00193_));
 sg13g2_mux2_1 _08789_ (.A0(\shift_storage.storage[1082] ),
    .A1(\shift_storage.storage[1081] ),
    .S(net718),
    .X(_03329_));
 sg13g2_and2_1 _08790_ (.A(net424),
    .B(_03329_),
    .X(_00194_));
 sg13g2_mux2_1 _08791_ (.A0(\shift_storage.storage[1083] ),
    .A1(\shift_storage.storage[1082] ),
    .S(net718),
    .X(_03330_));
 sg13g2_and2_1 _08792_ (.A(net424),
    .B(_03330_),
    .X(_00195_));
 sg13g2_buf_1 fanout353 (.A(net354),
    .X(net353));
 sg13g2_mux2_1 _08794_ (.A0(\shift_storage.storage[1084] ),
    .A1(\shift_storage.storage[1083] ),
    .S(net718),
    .X(_03332_));
 sg13g2_and2_1 _08795_ (.A(net420),
    .B(_03332_),
    .X(_00196_));
 sg13g2_mux2_1 _08796_ (.A0(\shift_storage.storage[1085] ),
    .A1(\shift_storage.storage[1084] ),
    .S(net714),
    .X(_03333_));
 sg13g2_and2_1 _08797_ (.A(net420),
    .B(_03333_),
    .X(_00197_));
 sg13g2_mux2_1 _08798_ (.A0(\shift_storage.storage[1086] ),
    .A1(\shift_storage.storage[1085] ),
    .S(net714),
    .X(_03334_));
 sg13g2_and2_1 _08799_ (.A(net420),
    .B(_03334_),
    .X(_00198_));
 sg13g2_mux2_1 _08800_ (.A0(\shift_storage.storage[1087] ),
    .A1(\shift_storage.storage[1086] ),
    .S(net714),
    .X(_03335_));
 sg13g2_and2_1 _08801_ (.A(net420),
    .B(_03335_),
    .X(_00199_));
 sg13g2_mux2_1 _08802_ (.A0(\shift_storage.storage[1088] ),
    .A1(\shift_storage.storage[1087] ),
    .S(net714),
    .X(_03336_));
 sg13g2_and2_1 _08803_ (.A(net420),
    .B(_03336_),
    .X(_00200_));
 sg13g2_mux2_1 _08804_ (.A0(\shift_storage.storage[1089] ),
    .A1(\shift_storage.storage[1088] ),
    .S(net714),
    .X(_03337_));
 sg13g2_and2_1 _08805_ (.A(net420),
    .B(_03337_),
    .X(_00201_));
 sg13g2_mux2_1 _08806_ (.A0(\shift_storage.storage[108] ),
    .A1(\shift_storage.storage[107] ),
    .S(net574),
    .X(_03338_));
 sg13g2_and2_1 _08807_ (.A(net274),
    .B(_03338_),
    .X(_00202_));
 sg13g2_buf_2 fanout352 (.A(net353),
    .X(net352));
 sg13g2_mux2_1 _08809_ (.A0(\shift_storage.storage[1090] ),
    .A1(\shift_storage.storage[1089] ),
    .S(net713),
    .X(_03340_));
 sg13g2_and2_1 _08810_ (.A(net419),
    .B(_03340_),
    .X(_00203_));
 sg13g2_mux2_1 _08811_ (.A0(\shift_storage.storage[1091] ),
    .A1(\shift_storage.storage[1090] ),
    .S(net713),
    .X(_03341_));
 sg13g2_and2_1 _08812_ (.A(net419),
    .B(_03341_),
    .X(_00204_));
 sg13g2_mux2_1 _08813_ (.A0(\shift_storage.storage[1092] ),
    .A1(\shift_storage.storage[1091] ),
    .S(net684),
    .X(_03342_));
 sg13g2_and2_1 _08814_ (.A(net389),
    .B(_03342_),
    .X(_00205_));
 sg13g2_buf_2 fanout351 (.A(net353),
    .X(net351));
 sg13g2_mux2_1 _08816_ (.A0(\shift_storage.storage[1093] ),
    .A1(\shift_storage.storage[1092] ),
    .S(net684),
    .X(_03344_));
 sg13g2_and2_1 _08817_ (.A(net389),
    .B(_03344_),
    .X(_00206_));
 sg13g2_mux2_1 _08818_ (.A0(\shift_storage.storage[1094] ),
    .A1(\shift_storage.storage[1093] ),
    .S(net684),
    .X(_03345_));
 sg13g2_and2_1 _08819_ (.A(net389),
    .B(_03345_),
    .X(_00207_));
 sg13g2_mux2_1 _08820_ (.A0(\shift_storage.storage[1095] ),
    .A1(\shift_storage.storage[1094] ),
    .S(net685),
    .X(_03346_));
 sg13g2_and2_1 _08821_ (.A(net390),
    .B(_03346_),
    .X(_00208_));
 sg13g2_mux2_1 _08822_ (.A0(\shift_storage.storage[1096] ),
    .A1(\shift_storage.storage[1095] ),
    .S(net685),
    .X(_03347_));
 sg13g2_and2_1 _08823_ (.A(net390),
    .B(_03347_),
    .X(_00209_));
 sg13g2_mux2_1 _08824_ (.A0(\shift_storage.storage[1097] ),
    .A1(\shift_storage.storage[1096] ),
    .S(net685),
    .X(_03348_));
 sg13g2_and2_1 _08825_ (.A(net390),
    .B(_03348_),
    .X(_00210_));
 sg13g2_mux2_1 _08826_ (.A0(\shift_storage.storage[1098] ),
    .A1(\shift_storage.storage[1097] ),
    .S(net685),
    .X(_03349_));
 sg13g2_and2_1 _08827_ (.A(net390),
    .B(_03349_),
    .X(_00211_));
 sg13g2_mux2_1 _08828_ (.A0(\shift_storage.storage[1099] ),
    .A1(\shift_storage.storage[1098] ),
    .S(net685),
    .X(_03350_));
 sg13g2_and2_1 _08829_ (.A(net390),
    .B(_03350_),
    .X(_00212_));
 sg13g2_buf_1 fanout350 (.A(net354),
    .X(net350));
 sg13g2_mux2_1 _08831_ (.A0(\shift_storage.storage[109] ),
    .A1(\shift_storage.storage[108] ),
    .S(net574),
    .X(_03352_));
 sg13g2_and2_1 _08832_ (.A(net274),
    .B(_03352_),
    .X(_00213_));
 sg13g2_mux2_1 _08833_ (.A0(\shift_storage.storage[10] ),
    .A1(\shift_storage.storage[9] ),
    .S(net609),
    .X(_03353_));
 sg13g2_and2_1 _08834_ (.A(net311),
    .B(_03353_),
    .X(_00214_));
 sg13g2_mux2_1 _08835_ (.A0(\shift_storage.storage[1100] ),
    .A1(\shift_storage.storage[1099] ),
    .S(net683),
    .X(_03354_));
 sg13g2_and2_1 _08836_ (.A(net388),
    .B(_03354_),
    .X(_00215_));
 sg13g2_buf_2 fanout349 (.A(net354),
    .X(net349));
 sg13g2_mux2_1 _08838_ (.A0(\shift_storage.storage[1101] ),
    .A1(\shift_storage.storage[1100] ),
    .S(net683),
    .X(_03356_));
 sg13g2_and2_1 _08839_ (.A(net388),
    .B(_03356_),
    .X(_00216_));
 sg13g2_mux2_1 _08840_ (.A0(\shift_storage.storage[1102] ),
    .A1(\shift_storage.storage[1101] ),
    .S(net682),
    .X(_03357_));
 sg13g2_and2_1 _08841_ (.A(net387),
    .B(_03357_),
    .X(_00217_));
 sg13g2_mux2_1 _08842_ (.A0(\shift_storage.storage[1103] ),
    .A1(\shift_storage.storage[1102] ),
    .S(net682),
    .X(_03358_));
 sg13g2_and2_1 _08843_ (.A(net387),
    .B(_03358_),
    .X(_00218_));
 sg13g2_mux2_1 _08844_ (.A0(\shift_storage.storage[1104] ),
    .A1(\shift_storage.storage[1103] ),
    .S(net682),
    .X(_03359_));
 sg13g2_and2_1 _08845_ (.A(net387),
    .B(_03359_),
    .X(_00219_));
 sg13g2_mux2_1 _08846_ (.A0(\shift_storage.storage[1105] ),
    .A1(\shift_storage.storage[1104] ),
    .S(net682),
    .X(_03360_));
 sg13g2_and2_1 _08847_ (.A(net387),
    .B(_03360_),
    .X(_00220_));
 sg13g2_mux2_1 _08848_ (.A0(\shift_storage.storage[1106] ),
    .A1(\shift_storage.storage[1105] ),
    .S(net675),
    .X(_03361_));
 sg13g2_and2_1 _08849_ (.A(net380),
    .B(_03361_),
    .X(_00221_));
 sg13g2_mux2_1 _08850_ (.A0(\shift_storage.storage[1107] ),
    .A1(\shift_storage.storage[1106] ),
    .S(net675),
    .X(_03362_));
 sg13g2_and2_1 _08851_ (.A(net379),
    .B(_03362_),
    .X(_00222_));
 sg13g2_buf_2 fanout348 (.A(net355),
    .X(net348));
 sg13g2_mux2_1 _08853_ (.A0(\shift_storage.storage[1108] ),
    .A1(\shift_storage.storage[1107] ),
    .S(net674),
    .X(_03364_));
 sg13g2_and2_1 _08854_ (.A(net379),
    .B(_03364_),
    .X(_00223_));
 sg13g2_mux2_1 _08855_ (.A0(\shift_storage.storage[1109] ),
    .A1(\shift_storage.storage[1108] ),
    .S(net674),
    .X(_03365_));
 sg13g2_and2_1 _08856_ (.A(net379),
    .B(_03365_),
    .X(_00224_));
 sg13g2_mux2_1 _08857_ (.A0(\shift_storage.storage[110] ),
    .A1(\shift_storage.storage[109] ),
    .S(net574),
    .X(_03366_));
 sg13g2_and2_1 _08858_ (.A(net274),
    .B(_03366_),
    .X(_00225_));
 sg13g2_buf_1 fanout347 (.A(net355),
    .X(net347));
 sg13g2_mux2_1 _08860_ (.A0(\shift_storage.storage[1110] ),
    .A1(\shift_storage.storage[1109] ),
    .S(net681),
    .X(_03368_));
 sg13g2_and2_1 _08861_ (.A(net381),
    .B(_03368_),
    .X(_00226_));
 sg13g2_mux2_1 _08862_ (.A0(\shift_storage.storage[1111] ),
    .A1(\shift_storage.storage[1110] ),
    .S(net675),
    .X(_03369_));
 sg13g2_and2_1 _08863_ (.A(net380),
    .B(_03369_),
    .X(_00227_));
 sg13g2_mux2_1 _08864_ (.A0(\shift_storage.storage[1112] ),
    .A1(\shift_storage.storage[1111] ),
    .S(net675),
    .X(_03370_));
 sg13g2_and2_1 _08865_ (.A(net380),
    .B(_03370_),
    .X(_00228_));
 sg13g2_mux2_1 _08866_ (.A0(\shift_storage.storage[1113] ),
    .A1(\shift_storage.storage[1112] ),
    .S(net673),
    .X(_03371_));
 sg13g2_and2_1 _08867_ (.A(net378),
    .B(_03371_),
    .X(_00229_));
 sg13g2_mux2_1 _08868_ (.A0(\shift_storage.storage[1114] ),
    .A1(\shift_storage.storage[1113] ),
    .S(net673),
    .X(_03372_));
 sg13g2_and2_1 _08869_ (.A(net378),
    .B(_03372_),
    .X(_00230_));
 sg13g2_mux2_1 _08870_ (.A0(\shift_storage.storage[1115] ),
    .A1(\shift_storage.storage[1114] ),
    .S(net673),
    .X(_03373_));
 sg13g2_and2_1 _08871_ (.A(net378),
    .B(_03373_),
    .X(_00231_));
 sg13g2_mux2_1 _08872_ (.A0(\shift_storage.storage[1116] ),
    .A1(\shift_storage.storage[1115] ),
    .S(net673),
    .X(_03374_));
 sg13g2_and2_1 _08873_ (.A(net378),
    .B(_03374_),
    .X(_00232_));
 sg13g2_buf_1 fanout346 (.A(net347),
    .X(net346));
 sg13g2_mux2_1 _08875_ (.A0(\shift_storage.storage[1117] ),
    .A1(\shift_storage.storage[1116] ),
    .S(net673),
    .X(_03376_));
 sg13g2_and2_1 _08876_ (.A(net383),
    .B(_03376_),
    .X(_00233_));
 sg13g2_mux2_1 _08877_ (.A0(\shift_storage.storage[1118] ),
    .A1(\shift_storage.storage[1117] ),
    .S(net677),
    .X(_03377_));
 sg13g2_and2_1 _08878_ (.A(net383),
    .B(_03377_),
    .X(_00234_));
 sg13g2_mux2_1 _08879_ (.A0(\shift_storage.storage[1119] ),
    .A1(\shift_storage.storage[1118] ),
    .S(net678),
    .X(_03378_));
 sg13g2_and2_1 _08880_ (.A(net384),
    .B(_03378_),
    .X(_00235_));
 sg13g2_buf_1 fanout345 (.A(net347),
    .X(net345));
 sg13g2_mux2_1 _08882_ (.A0(\shift_storage.storage[111] ),
    .A1(\shift_storage.storage[110] ),
    .S(net574),
    .X(_03380_));
 sg13g2_and2_1 _08883_ (.A(net323),
    .B(_03380_),
    .X(_00236_));
 sg13g2_mux2_1 _08884_ (.A0(\shift_storage.storage[1120] ),
    .A1(\shift_storage.storage[1119] ),
    .S(net678),
    .X(_03381_));
 sg13g2_and2_1 _08885_ (.A(net384),
    .B(_03381_),
    .X(_00237_));
 sg13g2_mux2_1 _08886_ (.A0(\shift_storage.storage[1121] ),
    .A1(\shift_storage.storage[1120] ),
    .S(net675),
    .X(_03382_));
 sg13g2_and2_1 _08887_ (.A(net380),
    .B(_03382_),
    .X(_00238_));
 sg13g2_mux2_1 _08888_ (.A0(\shift_storage.storage[1122] ),
    .A1(\shift_storage.storage[1121] ),
    .S(net675),
    .X(_03383_));
 sg13g2_and2_1 _08889_ (.A(net380),
    .B(_03383_),
    .X(_00239_));
 sg13g2_mux2_1 _08890_ (.A0(\shift_storage.storage[1123] ),
    .A1(\shift_storage.storage[1122] ),
    .S(net675),
    .X(_03384_));
 sg13g2_and2_1 _08891_ (.A(net381),
    .B(_03384_),
    .X(_00240_));
 sg13g2_mux2_1 _08892_ (.A0(\shift_storage.storage[1124] ),
    .A1(\shift_storage.storage[1123] ),
    .S(net683),
    .X(_03385_));
 sg13g2_and2_1 _08893_ (.A(net388),
    .B(_03385_),
    .X(_00241_));
 sg13g2_mux2_1 _08894_ (.A0(\shift_storage.storage[1125] ),
    .A1(\shift_storage.storage[1124] ),
    .S(net683),
    .X(_03386_));
 sg13g2_and2_1 _08895_ (.A(net388),
    .B(_03386_),
    .X(_00242_));
 sg13g2_buf_1 fanout344 (.A(net347),
    .X(net344));
 sg13g2_buf_2 fanout343 (.A(net347),
    .X(net343));
 sg13g2_mux2_1 _08898_ (.A0(\shift_storage.storage[1126] ),
    .A1(\shift_storage.storage[1125] ),
    .S(net683),
    .X(_03389_));
 sg13g2_and2_1 _08899_ (.A(net388),
    .B(_03389_),
    .X(_00243_));
 sg13g2_mux2_1 _08900_ (.A0(\shift_storage.storage[1127] ),
    .A1(\shift_storage.storage[1126] ),
    .S(net683),
    .X(_03390_));
 sg13g2_and2_1 _08901_ (.A(net388),
    .B(_03390_),
    .X(_00244_));
 sg13g2_mux2_1 _08902_ (.A0(\shift_storage.storage[1128] ),
    .A1(\shift_storage.storage[1127] ),
    .S(net683),
    .X(_03391_));
 sg13g2_and2_1 _08903_ (.A(net388),
    .B(_03391_),
    .X(_00245_));
 sg13g2_buf_1 fanout342 (.A(net356),
    .X(net342));
 sg13g2_buf_2 fanout341 (.A(net342),
    .X(net341));
 sg13g2_mux2_1 _08906_ (.A0(\shift_storage.storage[1129] ),
    .A1(\shift_storage.storage[1128] ),
    .S(net688),
    .X(_03394_));
 sg13g2_and2_1 _08907_ (.A(net392),
    .B(_03394_),
    .X(_00246_));
 sg13g2_mux2_1 _08908_ (.A0(\shift_storage.storage[112] ),
    .A1(\shift_storage.storage[111] ),
    .S(net622),
    .X(_03395_));
 sg13g2_and2_1 _08909_ (.A(net323),
    .B(_03395_),
    .X(_00247_));
 sg13g2_mux2_1 _08910_ (.A0(\shift_storage.storage[1130] ),
    .A1(\shift_storage.storage[1129] ),
    .S(net689),
    .X(_03396_));
 sg13g2_and2_1 _08911_ (.A(net395),
    .B(_03396_),
    .X(_00248_));
 sg13g2_mux2_1 _08912_ (.A0(\shift_storage.storage[1131] ),
    .A1(\shift_storage.storage[1130] ),
    .S(net689),
    .X(_03397_));
 sg13g2_and2_1 _08913_ (.A(net395),
    .B(_03397_),
    .X(_00249_));
 sg13g2_mux2_1 _08914_ (.A0(\shift_storage.storage[1132] ),
    .A1(\shift_storage.storage[1131] ),
    .S(net689),
    .X(_03398_));
 sg13g2_and2_1 _08915_ (.A(net390),
    .B(_03398_),
    .X(_00250_));
 sg13g2_mux2_1 _08916_ (.A0(\shift_storage.storage[1133] ),
    .A1(\shift_storage.storage[1132] ),
    .S(net685),
    .X(_03399_));
 sg13g2_and2_1 _08917_ (.A(net390),
    .B(_03399_),
    .X(_00251_));
 sg13g2_mux2_1 _08918_ (.A0(\shift_storage.storage[1134] ),
    .A1(\shift_storage.storage[1133] ),
    .S(net685),
    .X(_03400_));
 sg13g2_and2_1 _08919_ (.A(net390),
    .B(_03400_),
    .X(_00252_));
 sg13g2_buf_2 fanout340 (.A(net341),
    .X(net340));
 sg13g2_mux2_1 _08921_ (.A0(\shift_storage.storage[1135] ),
    .A1(\shift_storage.storage[1134] ),
    .S(net689),
    .X(_03402_));
 sg13g2_and2_1 _08922_ (.A(net395),
    .B(_03402_),
    .X(_00253_));
 sg13g2_mux2_1 _08923_ (.A0(\shift_storage.storage[1136] ),
    .A1(\shift_storage.storage[1135] ),
    .S(net691),
    .X(_03403_));
 sg13g2_and2_1 _08924_ (.A(net395),
    .B(_03403_),
    .X(_00254_));
 sg13g2_mux2_1 _08925_ (.A0(\shift_storage.storage[1137] ),
    .A1(\shift_storage.storage[1136] ),
    .S(net689),
    .X(_03404_));
 sg13g2_and2_1 _08926_ (.A(net395),
    .B(_03404_),
    .X(_00255_));
 sg13g2_buf_1 fanout339 (.A(net342),
    .X(net339));
 sg13g2_mux2_1 _08928_ (.A0(\shift_storage.storage[1138] ),
    .A1(\shift_storage.storage[1137] ),
    .S(net689),
    .X(_03406_));
 sg13g2_and2_1 _08929_ (.A(net395),
    .B(_03406_),
    .X(_00256_));
 sg13g2_mux2_1 _08930_ (.A0(\shift_storage.storage[1139] ),
    .A1(\shift_storage.storage[1138] ),
    .S(net691),
    .X(_03407_));
 sg13g2_and2_1 _08931_ (.A(net395),
    .B(_03407_),
    .X(_00257_));
 sg13g2_mux2_1 _08932_ (.A0(\shift_storage.storage[113] ),
    .A1(\shift_storage.storage[112] ),
    .S(net622),
    .X(_03408_));
 sg13g2_and2_1 _08933_ (.A(net325),
    .B(_03408_),
    .X(_00258_));
 sg13g2_mux2_1 _08934_ (.A0(\shift_storage.storage[1140] ),
    .A1(\shift_storage.storage[1139] ),
    .S(net690),
    .X(_03409_));
 sg13g2_and2_1 _08935_ (.A(net396),
    .B(_03409_),
    .X(_00259_));
 sg13g2_mux2_1 _08936_ (.A0(\shift_storage.storage[1141] ),
    .A1(\shift_storage.storage[1140] ),
    .S(net690),
    .X(_03410_));
 sg13g2_and2_1 _08937_ (.A(net394),
    .B(_03410_),
    .X(_00260_));
 sg13g2_mux2_1 _08938_ (.A0(\shift_storage.storage[1142] ),
    .A1(\shift_storage.storage[1141] ),
    .S(net719),
    .X(_03411_));
 sg13g2_and2_1 _08939_ (.A(net424),
    .B(_03411_),
    .X(_00261_));
 sg13g2_mux2_1 _08940_ (.A0(\shift_storage.storage[1143] ),
    .A1(\shift_storage.storage[1142] ),
    .S(net718),
    .X(_03412_));
 sg13g2_and2_1 _08941_ (.A(net424),
    .B(_03412_),
    .X(_00262_));
 sg13g2_buf_1 fanout338 (.A(net339),
    .X(net338));
 sg13g2_mux2_1 _08943_ (.A0(\shift_storage.storage[1144] ),
    .A1(\shift_storage.storage[1143] ),
    .S(net719),
    .X(_03414_));
 sg13g2_and2_1 _08944_ (.A(net425),
    .B(_03414_),
    .X(_00263_));
 sg13g2_mux2_1 _08945_ (.A0(\shift_storage.storage[1145] ),
    .A1(\shift_storage.storage[1144] ),
    .S(net719),
    .X(_03415_));
 sg13g2_and2_1 _08946_ (.A(net394),
    .B(_03415_),
    .X(_00264_));
 sg13g2_mux2_1 _08947_ (.A0(\shift_storage.storage[1146] ),
    .A1(\shift_storage.storage[1145] ),
    .S(net719),
    .X(_03416_));
 sg13g2_and2_1 _08948_ (.A(net394),
    .B(_03416_),
    .X(_00265_));
 sg13g2_buf_1 fanout337 (.A(net339),
    .X(net337));
 sg13g2_mux2_1 _08950_ (.A0(\shift_storage.storage[1147] ),
    .A1(\shift_storage.storage[1146] ),
    .S(net758),
    .X(_03418_));
 sg13g2_and2_1 _08951_ (.A(net471),
    .B(_03418_),
    .X(_00266_));
 sg13g2_mux2_1 _08952_ (.A0(\shift_storage.storage[1148] ),
    .A1(\shift_storage.storage[1147] ),
    .S(net758),
    .X(_03419_));
 sg13g2_and2_1 _08953_ (.A(net471),
    .B(_03419_),
    .X(_00267_));
 sg13g2_mux2_1 _08954_ (.A0(\shift_storage.storage[1149] ),
    .A1(\shift_storage.storage[1148] ),
    .S(net758),
    .X(_03420_));
 sg13g2_and2_1 _08955_ (.A(net471),
    .B(_03420_),
    .X(_00268_));
 sg13g2_mux2_1 _08956_ (.A0(\shift_storage.storage[114] ),
    .A1(\shift_storage.storage[113] ),
    .S(net630),
    .X(_03421_));
 sg13g2_and2_1 _08957_ (.A(net332),
    .B(_03421_),
    .X(_00269_));
 sg13g2_mux2_1 _08958_ (.A0(\shift_storage.storage[1150] ),
    .A1(\shift_storage.storage[1149] ),
    .S(net759),
    .X(_03422_));
 sg13g2_and2_1 _08959_ (.A(net472),
    .B(_03422_),
    .X(_00270_));
 sg13g2_mux2_1 _08960_ (.A0(\shift_storage.storage[1151] ),
    .A1(\shift_storage.storage[1150] ),
    .S(net758),
    .X(_03423_));
 sg13g2_and2_1 _08961_ (.A(net472),
    .B(_03423_),
    .X(_00271_));
 sg13g2_mux2_1 _08962_ (.A0(\shift_storage.storage[1152] ),
    .A1(\shift_storage.storage[1151] ),
    .S(net760),
    .X(_03424_));
 sg13g2_and2_1 _08963_ (.A(net473),
    .B(_03424_),
    .X(_00272_));
 sg13g2_buf_1 fanout336 (.A(net342),
    .X(net336));
 sg13g2_mux2_1 _08965_ (.A0(\shift_storage.storage[1153] ),
    .A1(\shift_storage.storage[1152] ),
    .S(net760),
    .X(_03426_));
 sg13g2_and2_1 _08966_ (.A(net473),
    .B(_03426_),
    .X(_00273_));
 sg13g2_mux2_1 _08967_ (.A0(\shift_storage.storage[1154] ),
    .A1(\shift_storage.storage[1153] ),
    .S(net760),
    .X(_03427_));
 sg13g2_and2_1 _08968_ (.A(net473),
    .B(_03427_),
    .X(_00274_));
 sg13g2_mux2_1 _08969_ (.A0(\shift_storage.storage[1155] ),
    .A1(\shift_storage.storage[1154] ),
    .S(net760),
    .X(_03428_));
 sg13g2_and2_1 _08970_ (.A(net473),
    .B(_03428_),
    .X(_00275_));
 sg13g2_buf_2 fanout335 (.A(net336),
    .X(net335));
 sg13g2_mux2_1 _08972_ (.A0(\shift_storage.storage[1156] ),
    .A1(\shift_storage.storage[1155] ),
    .S(net760),
    .X(_03430_));
 sg13g2_and2_1 _08973_ (.A(net473),
    .B(_03430_),
    .X(_00276_));
 sg13g2_mux2_1 _08974_ (.A0(\shift_storage.storage[1157] ),
    .A1(\shift_storage.storage[1156] ),
    .S(net760),
    .X(_03431_));
 sg13g2_and2_1 _08975_ (.A(net473),
    .B(_03431_),
    .X(_00277_));
 sg13g2_mux2_1 _08976_ (.A0(\shift_storage.storage[1158] ),
    .A1(\shift_storage.storage[1157] ),
    .S(net761),
    .X(_03432_));
 sg13g2_and2_1 _08977_ (.A(net474),
    .B(_03432_),
    .X(_00278_));
 sg13g2_mux2_1 _08978_ (.A0(\shift_storage.storage[1159] ),
    .A1(\shift_storage.storage[1158] ),
    .S(net761),
    .X(_03433_));
 sg13g2_and2_1 _08979_ (.A(net474),
    .B(_03433_),
    .X(_00279_));
 sg13g2_mux2_1 _08980_ (.A0(\shift_storage.storage[115] ),
    .A1(\shift_storage.storage[114] ),
    .S(net583),
    .X(_03434_));
 sg13g2_and2_1 _08981_ (.A(net283),
    .B(_03434_),
    .X(_00280_));
 sg13g2_mux2_1 _08982_ (.A0(\shift_storage.storage[1160] ),
    .A1(\shift_storage.storage[1159] ),
    .S(net765),
    .X(_03435_));
 sg13g2_and2_1 _08983_ (.A(net481),
    .B(_03435_),
    .X(_00281_));
 sg13g2_mux2_1 _08984_ (.A0(\shift_storage.storage[1161] ),
    .A1(\shift_storage.storage[1160] ),
    .S(net765),
    .X(_03436_));
 sg13g2_and2_1 _08985_ (.A(net481),
    .B(_03436_),
    .X(_00282_));
 sg13g2_buf_2 fanout334 (.A(net335),
    .X(net334));
 sg13g2_mux2_1 _08987_ (.A0(\shift_storage.storage[1162] ),
    .A1(\shift_storage.storage[1161] ),
    .S(net767),
    .X(_03438_));
 sg13g2_and2_1 _08988_ (.A(net483),
    .B(_03438_),
    .X(_00283_));
 sg13g2_mux2_1 _08989_ (.A0(\shift_storage.storage[1163] ),
    .A1(\shift_storage.storage[1162] ),
    .S(net765),
    .X(_03439_));
 sg13g2_and2_1 _08990_ (.A(net481),
    .B(_03439_),
    .X(_00284_));
 sg13g2_mux2_1 _08991_ (.A0(\shift_storage.storage[1164] ),
    .A1(\shift_storage.storage[1163] ),
    .S(net765),
    .X(_03440_));
 sg13g2_and2_1 _08992_ (.A(net481),
    .B(_03440_),
    .X(_00285_));
 sg13g2_buf_1 fanout333 (.A(net336),
    .X(net333));
 sg13g2_mux2_1 _08994_ (.A0(\shift_storage.storage[1165] ),
    .A1(\shift_storage.storage[1164] ),
    .S(net765),
    .X(_03442_));
 sg13g2_and2_1 _08995_ (.A(net481),
    .B(_03442_),
    .X(_00286_));
 sg13g2_mux2_1 _08996_ (.A0(\shift_storage.storage[1166] ),
    .A1(\shift_storage.storage[1165] ),
    .S(net765),
    .X(_03443_));
 sg13g2_and2_1 _08997_ (.A(net481),
    .B(_03443_),
    .X(_00287_));
 sg13g2_mux2_1 _08998_ (.A0(\shift_storage.storage[1167] ),
    .A1(\shift_storage.storage[1166] ),
    .S(net765),
    .X(_03444_));
 sg13g2_and2_1 _08999_ (.A(net481),
    .B(_03444_),
    .X(_00288_));
 sg13g2_mux2_1 _09000_ (.A0(\shift_storage.storage[1168] ),
    .A1(\shift_storage.storage[1167] ),
    .S(net765),
    .X(_03445_));
 sg13g2_and2_1 _09001_ (.A(net481),
    .B(_03445_),
    .X(_00289_));
 sg13g2_mux2_1 _09002_ (.A0(\shift_storage.storage[1169] ),
    .A1(\shift_storage.storage[1168] ),
    .S(net761),
    .X(_03446_));
 sg13g2_and2_1 _09003_ (.A(net474),
    .B(_03446_),
    .X(_00290_));
 sg13g2_mux2_1 _09004_ (.A0(\shift_storage.storage[116] ),
    .A1(\shift_storage.storage[115] ),
    .S(net583),
    .X(_03447_));
 sg13g2_and2_1 _09005_ (.A(net283),
    .B(_03447_),
    .X(_00291_));
 sg13g2_mux2_1 _09006_ (.A0(\shift_storage.storage[1170] ),
    .A1(\shift_storage.storage[1169] ),
    .S(net761),
    .X(_03448_));
 sg13g2_and2_1 _09007_ (.A(net474),
    .B(_03448_),
    .X(_00292_));
 sg13g2_buf_2 fanout332 (.A(net336),
    .X(net332));
 sg13g2_mux2_1 _09009_ (.A0(\shift_storage.storage[1171] ),
    .A1(\shift_storage.storage[1170] ),
    .S(net761),
    .X(_03450_));
 sg13g2_and2_1 _09010_ (.A(net474),
    .B(_03450_),
    .X(_00293_));
 sg13g2_mux2_1 _09011_ (.A0(\shift_storage.storage[1172] ),
    .A1(\shift_storage.storage[1171] ),
    .S(net761),
    .X(_03451_));
 sg13g2_and2_1 _09012_ (.A(net474),
    .B(_03451_),
    .X(_00294_));
 sg13g2_mux2_1 _09013_ (.A0(\shift_storage.storage[1173] ),
    .A1(\shift_storage.storage[1172] ),
    .S(net761),
    .X(_03452_));
 sg13g2_and2_1 _09014_ (.A(net475),
    .B(_03452_),
    .X(_00295_));
 sg13g2_buf_1 fanout331 (.A(net342),
    .X(net331));
 sg13g2_mux2_1 _09016_ (.A0(\shift_storage.storage[1174] ),
    .A1(\shift_storage.storage[1173] ),
    .S(net759),
    .X(_03454_));
 sg13g2_and2_1 _09017_ (.A(net472),
    .B(_03454_),
    .X(_00296_));
 sg13g2_mux2_1 _09018_ (.A0(\shift_storage.storage[1175] ),
    .A1(\shift_storage.storage[1174] ),
    .S(net759),
    .X(_03455_));
 sg13g2_and2_1 _09019_ (.A(net472),
    .B(_03455_),
    .X(_00297_));
 sg13g2_mux2_1 _09020_ (.A0(\shift_storage.storage[1176] ),
    .A1(\shift_storage.storage[1175] ),
    .S(net759),
    .X(_03456_));
 sg13g2_and2_1 _09021_ (.A(net472),
    .B(_03456_),
    .X(_00298_));
 sg13g2_mux2_1 _09022_ (.A0(\shift_storage.storage[1177] ),
    .A1(\shift_storage.storage[1176] ),
    .S(net759),
    .X(_03457_));
 sg13g2_and2_1 _09023_ (.A(net474),
    .B(_03457_),
    .X(_00299_));
 sg13g2_mux2_1 _09024_ (.A0(\shift_storage.storage[1178] ),
    .A1(\shift_storage.storage[1177] ),
    .S(net760),
    .X(_03458_));
 sg13g2_and2_1 _09025_ (.A(net473),
    .B(_03458_),
    .X(_00300_));
 sg13g2_mux2_1 _09026_ (.A0(\shift_storage.storage[1179] ),
    .A1(\shift_storage.storage[1178] ),
    .S(net760),
    .X(_03459_));
 sg13g2_and2_1 _09027_ (.A(net473),
    .B(_03459_),
    .X(_00301_));
 sg13g2_mux2_1 _09028_ (.A0(\shift_storage.storage[117] ),
    .A1(\shift_storage.storage[116] ),
    .S(net583),
    .X(_03460_));
 sg13g2_and2_1 _09029_ (.A(net283),
    .B(_03460_),
    .X(_00302_));
 sg13g2_buf_1 fanout330 (.A(net331),
    .X(net330));
 sg13g2_mux2_1 _09031_ (.A0(\shift_storage.storage[1180] ),
    .A1(\shift_storage.storage[1179] ),
    .S(net758),
    .X(_03462_));
 sg13g2_and2_1 _09032_ (.A(net471),
    .B(_03462_),
    .X(_00303_));
 sg13g2_mux2_1 _09033_ (.A0(\shift_storage.storage[1181] ),
    .A1(\shift_storage.storage[1180] ),
    .S(net759),
    .X(_03463_));
 sg13g2_and2_1 _09034_ (.A(net471),
    .B(_03463_),
    .X(_00304_));
 sg13g2_mux2_1 _09035_ (.A0(\shift_storage.storage[1182] ),
    .A1(\shift_storage.storage[1181] ),
    .S(net758),
    .X(_03464_));
 sg13g2_and2_1 _09036_ (.A(net471),
    .B(_03464_),
    .X(_00305_));
 sg13g2_buf_1 fanout329 (.A(net331),
    .X(net329));
 sg13g2_mux2_1 _09038_ (.A0(\shift_storage.storage[1183] ),
    .A1(\shift_storage.storage[1182] ),
    .S(net762),
    .X(_03466_));
 sg13g2_and2_1 _09039_ (.A(net472),
    .B(_03466_),
    .X(_00306_));
 sg13g2_mux2_1 _09040_ (.A0(\shift_storage.storage[1184] ),
    .A1(\shift_storage.storage[1183] ),
    .S(net758),
    .X(_03467_));
 sg13g2_and2_1 _09041_ (.A(net471),
    .B(_03467_),
    .X(_00307_));
 sg13g2_mux2_1 _09042_ (.A0(\shift_storage.storage[1185] ),
    .A1(\shift_storage.storage[1184] ),
    .S(net758),
    .X(_03468_));
 sg13g2_and2_1 _09043_ (.A(net471),
    .B(_03468_),
    .X(_00308_));
 sg13g2_mux2_1 _09044_ (.A0(\shift_storage.storage[1186] ),
    .A1(\shift_storage.storage[1185] ),
    .S(net742),
    .X(_03469_));
 sg13g2_and2_1 _09045_ (.A(net449),
    .B(_03469_),
    .X(_00309_));
 sg13g2_mux2_1 _09046_ (.A0(\shift_storage.storage[1187] ),
    .A1(\shift_storage.storage[1186] ),
    .S(net742),
    .X(_03470_));
 sg13g2_and2_1 _09047_ (.A(net449),
    .B(_03470_),
    .X(_00310_));
 sg13g2_mux2_1 _09048_ (.A0(\shift_storage.storage[1188] ),
    .A1(\shift_storage.storage[1187] ),
    .S(net742),
    .X(_03471_));
 sg13g2_and2_1 _09049_ (.A(net449),
    .B(_03471_),
    .X(_00311_));
 sg13g2_mux2_1 _09050_ (.A0(\shift_storage.storage[1189] ),
    .A1(\shift_storage.storage[1188] ),
    .S(net743),
    .X(_03472_));
 sg13g2_and2_1 _09051_ (.A(net449),
    .B(_03472_),
    .X(_00312_));
 sg13g2_buf_2 fanout328 (.A(net331),
    .X(net328));
 sg13g2_buf_1 fanout327 (.A(net328),
    .X(net327));
 sg13g2_mux2_1 _09054_ (.A0(\shift_storage.storage[118] ),
    .A1(\shift_storage.storage[117] ),
    .S(net585),
    .X(_03475_));
 sg13g2_and2_1 _09055_ (.A(net285),
    .B(_03475_),
    .X(_00313_));
 sg13g2_mux2_1 _09056_ (.A0(\shift_storage.storage[1190] ),
    .A1(\shift_storage.storage[1189] ),
    .S(net690),
    .X(_03476_));
 sg13g2_and2_1 _09057_ (.A(net396),
    .B(_03476_),
    .X(_00314_));
 sg13g2_mux2_1 _09058_ (.A0(\shift_storage.storage[1191] ),
    .A1(\shift_storage.storage[1190] ),
    .S(net691),
    .X(_03477_));
 sg13g2_and2_1 _09059_ (.A(net396),
    .B(_03477_),
    .X(_00315_));
 sg13g2_buf_1 fanout326 (.A(net342),
    .X(net326));
 sg13g2_buf_1 fanout325 (.A(net326),
    .X(net325));
 sg13g2_mux2_1 _09062_ (.A0(\shift_storage.storage[1192] ),
    .A1(\shift_storage.storage[1191] ),
    .S(net690),
    .X(_03480_));
 sg13g2_and2_1 _09063_ (.A(net394),
    .B(_03480_),
    .X(_00316_));
 sg13g2_mux2_1 _09064_ (.A0(\shift_storage.storage[1193] ),
    .A1(\shift_storage.storage[1192] ),
    .S(net690),
    .X(_03481_));
 sg13g2_and2_1 _09065_ (.A(net394),
    .B(_03481_),
    .X(_00317_));
 sg13g2_mux2_1 _09066_ (.A0(\shift_storage.storage[1194] ),
    .A1(\shift_storage.storage[1193] ),
    .S(net690),
    .X(_03482_));
 sg13g2_and2_1 _09067_ (.A(net394),
    .B(_03482_),
    .X(_00318_));
 sg13g2_mux2_1 _09068_ (.A0(\shift_storage.storage[1195] ),
    .A1(\shift_storage.storage[1194] ),
    .S(net689),
    .X(_03483_));
 sg13g2_and2_1 _09069_ (.A(net395),
    .B(_03483_),
    .X(_00319_));
 sg13g2_mux2_1 _09070_ (.A0(\shift_storage.storage[1196] ),
    .A1(\shift_storage.storage[1195] ),
    .S(net689),
    .X(_03484_));
 sg13g2_and2_1 _09071_ (.A(net392),
    .B(_03484_),
    .X(_00320_));
 sg13g2_mux2_1 _09072_ (.A0(\shift_storage.storage[1197] ),
    .A1(\shift_storage.storage[1196] ),
    .S(net688),
    .X(_03485_));
 sg13g2_and2_1 _09073_ (.A(net392),
    .B(_03485_),
    .X(_00321_));
 sg13g2_mux2_1 _09074_ (.A0(\shift_storage.storage[1198] ),
    .A1(\shift_storage.storage[1197] ),
    .S(net688),
    .X(_03486_));
 sg13g2_and2_1 _09075_ (.A(net392),
    .B(_03486_),
    .X(_00322_));
 sg13g2_buf_2 fanout324 (.A(net325),
    .X(net324));
 sg13g2_mux2_1 _09077_ (.A0(\shift_storage.storage[1199] ),
    .A1(\shift_storage.storage[1198] ),
    .S(net688),
    .X(_03488_));
 sg13g2_and2_1 _09078_ (.A(net392),
    .B(_03488_),
    .X(_00323_));
 sg13g2_mux2_1 _09079_ (.A0(\shift_storage.storage[119] ),
    .A1(\shift_storage.storage[118] ),
    .S(net585),
    .X(_03489_));
 sg13g2_and2_1 _09080_ (.A(net285),
    .B(_03489_),
    .X(_00324_));
 sg13g2_mux2_1 _09081_ (.A0(\shift_storage.storage[11] ),
    .A1(\shift_storage.storage[10] ),
    .S(net609),
    .X(_03490_));
 sg13g2_and2_1 _09082_ (.A(net311),
    .B(_03490_),
    .X(_00325_));
 sg13g2_buf_2 fanout323 (.A(net325),
    .X(net323));
 sg13g2_mux2_1 _09084_ (.A0(\shift_storage.storage[1200] ),
    .A1(\shift_storage.storage[1199] ),
    .S(net688),
    .X(_03492_));
 sg13g2_and2_1 _09085_ (.A(net392),
    .B(_03492_),
    .X(_00326_));
 sg13g2_mux2_1 _09086_ (.A0(\shift_storage.storage[1201] ),
    .A1(\shift_storage.storage[1200] ),
    .S(net688),
    .X(_03493_));
 sg13g2_and2_1 _09087_ (.A(net392),
    .B(_03493_),
    .X(_00327_));
 sg13g2_mux2_1 _09088_ (.A0(\shift_storage.storage[1202] ),
    .A1(\shift_storage.storage[1201] ),
    .S(net688),
    .X(_03494_));
 sg13g2_and2_1 _09089_ (.A(net380),
    .B(_03494_),
    .X(_00328_));
 sg13g2_mux2_1 _09090_ (.A0(\shift_storage.storage[1203] ),
    .A1(\shift_storage.storage[1202] ),
    .S(net679),
    .X(_03495_));
 sg13g2_and2_1 _09091_ (.A(net385),
    .B(_03495_),
    .X(_00329_));
 sg13g2_mux2_1 _09092_ (.A0(\shift_storage.storage[1204] ),
    .A1(\shift_storage.storage[1203] ),
    .S(net679),
    .X(_03496_));
 sg13g2_and2_1 _09093_ (.A(net384),
    .B(_03496_),
    .X(_00330_));
 sg13g2_mux2_1 _09094_ (.A0(\shift_storage.storage[1205] ),
    .A1(\shift_storage.storage[1204] ),
    .S(net678),
    .X(_03497_));
 sg13g2_and2_1 _09095_ (.A(net385),
    .B(_03497_),
    .X(_00331_));
 sg13g2_mux2_1 _09096_ (.A0(\shift_storage.storage[1206] ),
    .A1(\shift_storage.storage[1205] ),
    .S(net678),
    .X(_03498_));
 sg13g2_and2_1 _09097_ (.A(net384),
    .B(_03498_),
    .X(_00332_));
 sg13g2_buf_2 fanout322 (.A(net326),
    .X(net322));
 sg13g2_mux2_1 _09099_ (.A0(\shift_storage.storage[1207] ),
    .A1(\shift_storage.storage[1206] ),
    .S(net679),
    .X(_03500_));
 sg13g2_and2_1 _09100_ (.A(net386),
    .B(_03500_),
    .X(_00333_));
 sg13g2_mux2_1 _09101_ (.A0(\shift_storage.storage[1208] ),
    .A1(\shift_storage.storage[1207] ),
    .S(net679),
    .X(_03501_));
 sg13g2_and2_1 _09102_ (.A(net385),
    .B(_03501_),
    .X(_00334_));
 sg13g2_mux2_1 _09103_ (.A0(\shift_storage.storage[1209] ),
    .A1(\shift_storage.storage[1208] ),
    .S(net679),
    .X(_03502_));
 sg13g2_and2_1 _09104_ (.A(net385),
    .B(_03502_),
    .X(_00335_));
 sg13g2_buf_2 fanout321 (.A(net322),
    .X(net321));
 sg13g2_mux2_1 _09106_ (.A0(\shift_storage.storage[120] ),
    .A1(\shift_storage.storage[119] ),
    .S(net585),
    .X(_03504_));
 sg13g2_and2_1 _09107_ (.A(net285),
    .B(_03504_),
    .X(_00336_));
 sg13g2_mux2_1 _09108_ (.A0(\shift_storage.storage[1210] ),
    .A1(\shift_storage.storage[1209] ),
    .S(net680),
    .X(_03505_));
 sg13g2_and2_1 _09109_ (.A(net386),
    .B(_03505_),
    .X(_00337_));
 sg13g2_mux2_1 _09110_ (.A0(\shift_storage.storage[1211] ),
    .A1(\shift_storage.storage[1210] ),
    .S(net680),
    .X(_03506_));
 sg13g2_and2_1 _09111_ (.A(net385),
    .B(_03506_),
    .X(_00338_));
 sg13g2_mux2_1 _09112_ (.A0(\shift_storage.storage[1212] ),
    .A1(\shift_storage.storage[1211] ),
    .S(net679),
    .X(_03507_));
 sg13g2_and2_1 _09113_ (.A(net437),
    .B(_03507_),
    .X(_00339_));
 sg13g2_mux2_1 _09114_ (.A0(\shift_storage.storage[1213] ),
    .A1(\shift_storage.storage[1212] ),
    .S(net679),
    .X(_03508_));
 sg13g2_and2_1 _09115_ (.A(net385),
    .B(_03508_),
    .X(_00340_));
 sg13g2_mux2_1 _09116_ (.A0(\shift_storage.storage[1214] ),
    .A1(\shift_storage.storage[1213] ),
    .S(net687),
    .X(_03509_));
 sg13g2_and2_1 _09117_ (.A(net385),
    .B(_03509_),
    .X(_00341_));
 sg13g2_mux2_1 _09118_ (.A0(\shift_storage.storage[1215] ),
    .A1(\shift_storage.storage[1214] ),
    .S(net687),
    .X(_03510_));
 sg13g2_and2_1 _09119_ (.A(net393),
    .B(_03510_),
    .X(_00342_));
 sg13g2_buf_1 fanout320 (.A(net356),
    .X(net320));
 sg13g2_mux2_1 _09121_ (.A0(\shift_storage.storage[1216] ),
    .A1(\shift_storage.storage[1215] ),
    .S(net687),
    .X(_03512_));
 sg13g2_and2_1 _09122_ (.A(net392),
    .B(_03512_),
    .X(_00343_));
 sg13g2_mux2_1 _09123_ (.A0(\shift_storage.storage[1217] ),
    .A1(\shift_storage.storage[1216] ),
    .S(net741),
    .X(_03513_));
 sg13g2_and2_1 _09124_ (.A(net448),
    .B(_03513_),
    .X(_00344_));
 sg13g2_mux2_1 _09125_ (.A0(\shift_storage.storage[1218] ),
    .A1(\shift_storage.storage[1217] ),
    .S(net741),
    .X(_03514_));
 sg13g2_and2_1 _09126_ (.A(net446),
    .B(_03514_),
    .X(_00345_));
 sg13g2_buf_1 fanout319 (.A(net320),
    .X(net319));
 sg13g2_mux2_1 _09128_ (.A0(\shift_storage.storage[1219] ),
    .A1(\shift_storage.storage[1218] ),
    .S(net741),
    .X(_03516_));
 sg13g2_and2_1 _09129_ (.A(net446),
    .B(_03516_),
    .X(_00346_));
 sg13g2_mux2_1 _09130_ (.A0(\shift_storage.storage[121] ),
    .A1(\shift_storage.storage[120] ),
    .S(net585),
    .X(_03517_));
 sg13g2_and2_1 _09131_ (.A(net286),
    .B(_03517_),
    .X(_00347_));
 sg13g2_mux2_1 _09132_ (.A0(\shift_storage.storage[1220] ),
    .A1(\shift_storage.storage[1219] ),
    .S(net741),
    .X(_03518_));
 sg13g2_and2_1 _09133_ (.A(net446),
    .B(_03518_),
    .X(_00348_));
 sg13g2_mux2_1 _09134_ (.A0(\shift_storage.storage[1221] ),
    .A1(\shift_storage.storage[1220] ),
    .S(net741),
    .X(_03519_));
 sg13g2_and2_1 _09135_ (.A(net446),
    .B(_03519_),
    .X(_00349_));
 sg13g2_mux2_1 _09136_ (.A0(\shift_storage.storage[1222] ),
    .A1(\shift_storage.storage[1221] ),
    .S(net741),
    .X(_03520_));
 sg13g2_and2_1 _09137_ (.A(net446),
    .B(_03520_),
    .X(_00350_));
 sg13g2_mux2_1 _09138_ (.A0(\shift_storage.storage[1223] ),
    .A1(\shift_storage.storage[1222] ),
    .S(net744),
    .X(_03521_));
 sg13g2_and2_1 _09139_ (.A(net450),
    .B(_03521_),
    .X(_00351_));
 sg13g2_mux2_1 _09140_ (.A0(\shift_storage.storage[1224] ),
    .A1(\shift_storage.storage[1223] ),
    .S(net744),
    .X(_03522_));
 sg13g2_and2_1 _09141_ (.A(net450),
    .B(_03522_),
    .X(_00352_));
 sg13g2_buf_1 fanout318 (.A(net319),
    .X(net318));
 sg13g2_mux2_1 _09143_ (.A0(\shift_storage.storage[1225] ),
    .A1(\shift_storage.storage[1224] ),
    .S(net740),
    .X(_03524_));
 sg13g2_and2_1 _09144_ (.A(net447),
    .B(_03524_),
    .X(_00353_));
 sg13g2_mux2_1 _09145_ (.A0(\shift_storage.storage[1226] ),
    .A1(\shift_storage.storage[1225] ),
    .S(net740),
    .X(_03525_));
 sg13g2_and2_1 _09146_ (.A(net448),
    .B(_03525_),
    .X(_00354_));
 sg13g2_mux2_1 _09147_ (.A0(\shift_storage.storage[1227] ),
    .A1(\shift_storage.storage[1226] ),
    .S(net740),
    .X(_03526_));
 sg13g2_and2_1 _09148_ (.A(net447),
    .B(_03526_),
    .X(_00355_));
 sg13g2_buf_2 fanout317 (.A(net318),
    .X(net317));
 sg13g2_mux2_1 _09150_ (.A0(\shift_storage.storage[1228] ),
    .A1(\shift_storage.storage[1227] ),
    .S(net740),
    .X(_03528_));
 sg13g2_and2_1 _09151_ (.A(net447),
    .B(_03528_),
    .X(_00356_));
 sg13g2_mux2_1 _09152_ (.A0(\shift_storage.storage[1229] ),
    .A1(\shift_storage.storage[1228] ),
    .S(net740),
    .X(_03529_));
 sg13g2_and2_1 _09153_ (.A(net447),
    .B(_03529_),
    .X(_00357_));
 sg13g2_mux2_1 _09154_ (.A0(\shift_storage.storage[122] ),
    .A1(\shift_storage.storage[121] ),
    .S(net585),
    .X(_03530_));
 sg13g2_and2_1 _09155_ (.A(net285),
    .B(_03530_),
    .X(_00358_));
 sg13g2_mux2_1 _09156_ (.A0(\shift_storage.storage[1230] ),
    .A1(\shift_storage.storage[1229] ),
    .S(net741),
    .X(_03531_));
 sg13g2_and2_1 _09157_ (.A(net446),
    .B(_03531_),
    .X(_00359_));
 sg13g2_mux2_1 _09158_ (.A0(\shift_storage.storage[1231] ),
    .A1(\shift_storage.storage[1230] ),
    .S(net741),
    .X(_03532_));
 sg13g2_and2_1 _09159_ (.A(net446),
    .B(_03532_),
    .X(_00360_));
 sg13g2_mux2_1 _09160_ (.A0(\shift_storage.storage[1232] ),
    .A1(\shift_storage.storage[1231] ),
    .S(net731),
    .X(_03533_));
 sg13g2_and2_1 _09161_ (.A(net437),
    .B(_03533_),
    .X(_00361_));
 sg13g2_mux2_1 _09162_ (.A0(\shift_storage.storage[1233] ),
    .A1(\shift_storage.storage[1232] ),
    .S(net731),
    .X(_03534_));
 sg13g2_and2_1 _09163_ (.A(net437),
    .B(_03534_),
    .X(_00362_));
 sg13g2_buf_2 fanout316 (.A(net317),
    .X(net316));
 sg13g2_mux2_1 _09165_ (.A0(\shift_storage.storage[1234] ),
    .A1(\shift_storage.storage[1233] ),
    .S(net731),
    .X(_03536_));
 sg13g2_and2_1 _09166_ (.A(net437),
    .B(_03536_),
    .X(_00363_));
 sg13g2_mux2_1 _09167_ (.A0(\shift_storage.storage[1235] ),
    .A1(\shift_storage.storage[1234] ),
    .S(net731),
    .X(_03537_));
 sg13g2_and2_1 _09168_ (.A(net437),
    .B(_03537_),
    .X(_00364_));
 sg13g2_mux2_1 _09169_ (.A0(\shift_storage.storage[1236] ),
    .A1(\shift_storage.storage[1235] ),
    .S(net731),
    .X(_03538_));
 sg13g2_and2_1 _09170_ (.A(net435),
    .B(_03538_),
    .X(_00365_));
 sg13g2_buf_1 fanout315 (.A(net320),
    .X(net315));
 sg13g2_mux2_1 _09172_ (.A0(\shift_storage.storage[1237] ),
    .A1(\shift_storage.storage[1236] ),
    .S(net730),
    .X(_03540_));
 sg13g2_and2_1 _09173_ (.A(net435),
    .B(_03540_),
    .X(_00366_));
 sg13g2_mux2_1 _09174_ (.A0(\shift_storage.storage[1238] ),
    .A1(\shift_storage.storage[1237] ),
    .S(net730),
    .X(_03541_));
 sg13g2_and2_1 _09175_ (.A(net435),
    .B(_03541_),
    .X(_00367_));
 sg13g2_mux2_1 _09176_ (.A0(\shift_storage.storage[1239] ),
    .A1(\shift_storage.storage[1238] ),
    .S(net730),
    .X(_03542_));
 sg13g2_and2_1 _09177_ (.A(net435),
    .B(_03542_),
    .X(_00368_));
 sg13g2_mux2_1 _09178_ (.A0(\shift_storage.storage[123] ),
    .A1(\shift_storage.storage[122] ),
    .S(net585),
    .X(_03543_));
 sg13g2_and2_1 _09179_ (.A(net285),
    .B(_03543_),
    .X(_00369_));
 sg13g2_mux2_1 _09180_ (.A0(\shift_storage.storage[1240] ),
    .A1(\shift_storage.storage[1239] ),
    .S(net729),
    .X(_03544_));
 sg13g2_and2_1 _09181_ (.A(net436),
    .B(_03544_),
    .X(_00370_));
 sg13g2_mux2_1 _09182_ (.A0(\shift_storage.storage[1241] ),
    .A1(\shift_storage.storage[1240] ),
    .S(net733),
    .X(_03545_));
 sg13g2_and2_1 _09183_ (.A(net436),
    .B(_03545_),
    .X(_00371_));
 sg13g2_mux2_1 _09184_ (.A0(\shift_storage.storage[1242] ),
    .A1(\shift_storage.storage[1241] ),
    .S(net729),
    .X(_03546_));
 sg13g2_and2_1 _09185_ (.A(net436),
    .B(_03546_),
    .X(_00372_));
 sg13g2_buf_2 fanout314 (.A(net315),
    .X(net314));
 sg13g2_mux2_1 _09187_ (.A0(\shift_storage.storage[1243] ),
    .A1(\shift_storage.storage[1242] ),
    .S(net729),
    .X(_03548_));
 sg13g2_and2_1 _09188_ (.A(net436),
    .B(_03548_),
    .X(_00373_));
 sg13g2_mux2_1 _09189_ (.A0(\shift_storage.storage[1244] ),
    .A1(\shift_storage.storage[1243] ),
    .S(net729),
    .X(_03549_));
 sg13g2_and2_1 _09190_ (.A(net442),
    .B(_03549_),
    .X(_00374_));
 sg13g2_mux2_1 _09191_ (.A0(\shift_storage.storage[1245] ),
    .A1(\shift_storage.storage[1244] ),
    .S(net734),
    .X(_03550_));
 sg13g2_and2_1 _09192_ (.A(net440),
    .B(_03550_),
    .X(_00375_));
 sg13g2_buf_1 fanout313 (.A(net320),
    .X(net313));
 sg13g2_mux2_1 _09194_ (.A0(\shift_storage.storage[1246] ),
    .A1(\shift_storage.storage[1245] ),
    .S(net734),
    .X(_03552_));
 sg13g2_and2_1 _09195_ (.A(net440),
    .B(_03552_),
    .X(_00376_));
 sg13g2_mux2_1 _09196_ (.A0(\shift_storage.storage[1247] ),
    .A1(\shift_storage.storage[1246] ),
    .S(net734),
    .X(_03553_));
 sg13g2_and2_1 _09197_ (.A(net440),
    .B(_03553_),
    .X(_00377_));
 sg13g2_mux2_1 _09198_ (.A0(\shift_storage.storage[1248] ),
    .A1(\shift_storage.storage[1247] ),
    .S(net734),
    .X(_03554_));
 sg13g2_and2_1 _09199_ (.A(net440),
    .B(_03554_),
    .X(_00378_));
 sg13g2_mux2_1 _09200_ (.A0(\shift_storage.storage[1249] ),
    .A1(\shift_storage.storage[1248] ),
    .S(net734),
    .X(_03555_));
 sg13g2_and2_1 _09201_ (.A(net340),
    .B(_03555_),
    .X(_00379_));
 sg13g2_mux2_1 _09202_ (.A0(\shift_storage.storage[124] ),
    .A1(\shift_storage.storage[123] ),
    .S(net585),
    .X(_03556_));
 sg13g2_and2_1 _09203_ (.A(net283),
    .B(_03556_),
    .X(_00380_));
 sg13g2_mux2_1 _09204_ (.A0(\shift_storage.storage[1250] ),
    .A1(\shift_storage.storage[1249] ),
    .S(net734),
    .X(_03557_));
 sg13g2_and2_1 _09205_ (.A(net440),
    .B(_03557_),
    .X(_00381_));
 sg13g2_mux2_1 _09206_ (.A0(\shift_storage.storage[1251] ),
    .A1(\shift_storage.storage[1250] ),
    .S(net735),
    .X(_03558_));
 sg13g2_and2_1 _09207_ (.A(net441),
    .B(_03558_),
    .X(_00382_));
 sg13g2_buf_1 fanout312 (.A(net313),
    .X(net312));
 sg13g2_buf_1 fanout311 (.A(net312),
    .X(net311));
 sg13g2_mux2_1 _09210_ (.A0(\shift_storage.storage[1252] ),
    .A1(\shift_storage.storage[1251] ),
    .S(net735),
    .X(_03561_));
 sg13g2_and2_1 _09211_ (.A(net441),
    .B(_03561_),
    .X(_00383_));
 sg13g2_mux2_1 _09212_ (.A0(\shift_storage.storage[1253] ),
    .A1(\shift_storage.storage[1252] ),
    .S(net735),
    .X(_03562_));
 sg13g2_and2_1 _09213_ (.A(net441),
    .B(_03562_),
    .X(_00384_));
 sg13g2_mux2_1 _09214_ (.A0(\shift_storage.storage[1254] ),
    .A1(\shift_storage.storage[1253] ),
    .S(net735),
    .X(_03563_));
 sg13g2_and2_1 _09215_ (.A(net441),
    .B(_03563_),
    .X(_00385_));
 sg13g2_buf_2 fanout310 (.A(net313),
    .X(net310));
 sg13g2_buf_1 fanout309 (.A(net320),
    .X(net309));
 sg13g2_mux2_1 _09218_ (.A0(\shift_storage.storage[1255] ),
    .A1(\shift_storage.storage[1254] ),
    .S(net735),
    .X(_03566_));
 sg13g2_and2_1 _09219_ (.A(net441),
    .B(_03566_),
    .X(_00386_));
 sg13g2_mux2_1 _09220_ (.A0(\shift_storage.storage[1256] ),
    .A1(\shift_storage.storage[1255] ),
    .S(net746),
    .X(_03567_));
 sg13g2_and2_1 _09221_ (.A(net455),
    .B(_03567_),
    .X(_00387_));
 sg13g2_mux2_1 _09222_ (.A0(\shift_storage.storage[1257] ),
    .A1(\shift_storage.storage[1256] ),
    .S(net649),
    .X(_03568_));
 sg13g2_and2_1 _09223_ (.A(net351),
    .B(_03568_),
    .X(_00388_));
 sg13g2_mux2_1 _09224_ (.A0(\shift_storage.storage[1258] ),
    .A1(\shift_storage.storage[1257] ),
    .S(net651),
    .X(_03569_));
 sg13g2_and2_1 _09225_ (.A(net353),
    .B(_03569_),
    .X(_00389_));
 sg13g2_mux2_1 _09226_ (.A0(\shift_storage.storage[1259] ),
    .A1(\shift_storage.storage[1258] ),
    .S(net649),
    .X(_03570_));
 sg13g2_and2_1 _09227_ (.A(net351),
    .B(_03570_),
    .X(_00390_));
 sg13g2_mux2_1 _09228_ (.A0(\shift_storage.storage[125] ),
    .A1(\shift_storage.storage[124] ),
    .S(net583),
    .X(_03571_));
 sg13g2_and2_1 _09229_ (.A(net287),
    .B(_03571_),
    .X(_00391_));
 sg13g2_mux2_1 _09230_ (.A0(\shift_storage.storage[1260] ),
    .A1(\shift_storage.storage[1259] ),
    .S(net649),
    .X(_03572_));
 sg13g2_and2_1 _09231_ (.A(net351),
    .B(_03572_),
    .X(_00392_));
 sg13g2_buf_2 fanout308 (.A(net309),
    .X(net308));
 sg13g2_mux2_1 _09233_ (.A0(\shift_storage.storage[1261] ),
    .A1(\shift_storage.storage[1260] ),
    .S(net649),
    .X(_03574_));
 sg13g2_and2_1 _09234_ (.A(net351),
    .B(_03574_),
    .X(_00393_));
 sg13g2_mux2_1 _09235_ (.A0(\shift_storage.storage[1262] ),
    .A1(\shift_storage.storage[1261] ),
    .S(net649),
    .X(_03575_));
 sg13g2_and2_1 _09236_ (.A(net351),
    .B(_03575_),
    .X(_00394_));
 sg13g2_mux2_1 _09237_ (.A0(\shift_storage.storage[1263] ),
    .A1(\shift_storage.storage[1262] ),
    .S(net650),
    .X(_03576_));
 sg13g2_and2_1 _09238_ (.A(net352),
    .B(_03576_),
    .X(_00395_));
 sg13g2_buf_1 fanout307 (.A(net308),
    .X(net307));
 sg13g2_mux2_1 _09240_ (.A0(\shift_storage.storage[1264] ),
    .A1(\shift_storage.storage[1263] ),
    .S(net650),
    .X(_03578_));
 sg13g2_and2_1 _09241_ (.A(net352),
    .B(_03578_),
    .X(_00396_));
 sg13g2_mux2_1 _09242_ (.A0(\shift_storage.storage[1265] ),
    .A1(\shift_storage.storage[1264] ),
    .S(net650),
    .X(_03579_));
 sg13g2_and2_1 _09243_ (.A(net352),
    .B(_03579_),
    .X(_00397_));
 sg13g2_mux2_1 _09244_ (.A0(\shift_storage.storage[1266] ),
    .A1(\shift_storage.storage[1265] ),
    .S(net650),
    .X(_03580_));
 sg13g2_and2_1 _09245_ (.A(net352),
    .B(_03580_),
    .X(_00398_));
 sg13g2_mux2_1 _09246_ (.A0(\shift_storage.storage[1267] ),
    .A1(\shift_storage.storage[1266] ),
    .S(net650),
    .X(_03581_));
 sg13g2_and2_1 _09247_ (.A(net352),
    .B(_03581_),
    .X(_00399_));
 sg13g2_mux2_1 _09248_ (.A0(\shift_storage.storage[1268] ),
    .A1(\shift_storage.storage[1267] ),
    .S(net650),
    .X(_03582_));
 sg13g2_and2_1 _09249_ (.A(net352),
    .B(_03582_),
    .X(_00400_));
 sg13g2_mux2_1 _09250_ (.A0(\shift_storage.storage[1269] ),
    .A1(\shift_storage.storage[1268] ),
    .S(net650),
    .X(_03583_));
 sg13g2_and2_1 _09251_ (.A(net352),
    .B(_03583_),
    .X(_00401_));
 sg13g2_mux2_1 _09252_ (.A0(\shift_storage.storage[126] ),
    .A1(\shift_storage.storage[125] ),
    .S(net587),
    .X(_03584_));
 sg13g2_and2_1 _09253_ (.A(net287),
    .B(_03584_),
    .X(_00402_));
 sg13g2_buf_1 fanout306 (.A(net307),
    .X(net306));
 sg13g2_mux2_1 _09255_ (.A0(\shift_storage.storage[1270] ),
    .A1(\shift_storage.storage[1269] ),
    .S(net650),
    .X(_03586_));
 sg13g2_and2_1 _09256_ (.A(net352),
    .B(_03586_),
    .X(_00403_));
 sg13g2_mux2_1 _09257_ (.A0(\shift_storage.storage[1271] ),
    .A1(\shift_storage.storage[1270] ),
    .S(net651),
    .X(_03587_));
 sg13g2_and2_1 _09258_ (.A(net353),
    .B(_03587_),
    .X(_00404_));
 sg13g2_mux2_1 _09259_ (.A0(\shift_storage.storage[1272] ),
    .A1(\shift_storage.storage[1271] ),
    .S(net749),
    .X(_03588_));
 sg13g2_and2_1 _09260_ (.A(net459),
    .B(_03588_),
    .X(_00405_));
 sg13g2_buf_1 fanout305 (.A(net309),
    .X(net305));
 sg13g2_mux2_1 _09262_ (.A0(\shift_storage.storage[1273] ),
    .A1(\shift_storage.storage[1272] ),
    .S(net746),
    .X(_03590_));
 sg13g2_and2_1 _09263_ (.A(net455),
    .B(_03590_),
    .X(_00406_));
 sg13g2_mux2_1 _09264_ (.A0(\shift_storage.storage[1274] ),
    .A1(\shift_storage.storage[1273] ),
    .S(net746),
    .X(_03591_));
 sg13g2_and2_1 _09265_ (.A(net455),
    .B(_03591_),
    .X(_00407_));
 sg13g2_mux2_1 _09266_ (.A0(\shift_storage.storage[1275] ),
    .A1(\shift_storage.storage[1274] ),
    .S(net746),
    .X(_03592_));
 sg13g2_and2_1 _09267_ (.A(net455),
    .B(_03592_),
    .X(_00408_));
 sg13g2_mux2_1 _09268_ (.A0(\shift_storage.storage[1276] ),
    .A1(\shift_storage.storage[1275] ),
    .S(net746),
    .X(_03593_));
 sg13g2_and2_1 _09269_ (.A(net455),
    .B(_03593_),
    .X(_00409_));
 sg13g2_mux2_1 _09270_ (.A0(\shift_storage.storage[1277] ),
    .A1(\shift_storage.storage[1276] ),
    .S(net746),
    .X(_03594_));
 sg13g2_and2_1 _09271_ (.A(net455),
    .B(_03594_),
    .X(_00410_));
 sg13g2_mux2_1 _09272_ (.A0(\shift_storage.storage[1278] ),
    .A1(\shift_storage.storage[1277] ),
    .S(net746),
    .X(_03595_));
 sg13g2_and2_1 _09273_ (.A(net455),
    .B(_03595_),
    .X(_00411_));
 sg13g2_mux2_1 _09274_ (.A0(\shift_storage.storage[1279] ),
    .A1(\shift_storage.storage[1278] ),
    .S(net735),
    .X(_03596_));
 sg13g2_and2_1 _09275_ (.A(net442),
    .B(_03596_),
    .X(_00412_));
 sg13g2_buf_1 fanout304 (.A(net305),
    .X(net304));
 sg13g2_mux2_1 _09277_ (.A0(\shift_storage.storage[127] ),
    .A1(\shift_storage.storage[126] ),
    .S(net583),
    .X(_03598_));
 sg13g2_and2_1 _09278_ (.A(net283),
    .B(_03598_),
    .X(_00413_));
 sg13g2_mux2_1 _09279_ (.A0(\shift_storage.storage[1280] ),
    .A1(\shift_storage.storage[1279] ),
    .S(net736),
    .X(_03599_));
 sg13g2_and2_1 _09280_ (.A(net442),
    .B(_03599_),
    .X(_00414_));
 sg13g2_mux2_1 _09281_ (.A0(\shift_storage.storage[1281] ),
    .A1(\shift_storage.storage[1280] ),
    .S(net738),
    .X(_03600_));
 sg13g2_and2_1 _09282_ (.A(net445),
    .B(_03600_),
    .X(_00415_));
 sg13g2_buf_1 fanout303 (.A(net305),
    .X(net303));
 sg13g2_mux2_1 _09284_ (.A0(\shift_storage.storage[1282] ),
    .A1(\shift_storage.storage[1281] ),
    .S(net747),
    .X(_03602_));
 sg13g2_and2_1 _09285_ (.A(net456),
    .B(_03602_),
    .X(_00416_));
 sg13g2_mux2_1 _09286_ (.A0(\shift_storage.storage[1283] ),
    .A1(\shift_storage.storage[1282] ),
    .S(net747),
    .X(_03603_));
 sg13g2_and2_1 _09287_ (.A(net456),
    .B(_03603_),
    .X(_00417_));
 sg13g2_mux2_1 _09288_ (.A0(\shift_storage.storage[1284] ),
    .A1(\shift_storage.storage[1283] ),
    .S(net747),
    .X(_03604_));
 sg13g2_and2_1 _09289_ (.A(net456),
    .B(_03604_),
    .X(_00418_));
 sg13g2_mux2_1 _09290_ (.A0(\shift_storage.storage[1285] ),
    .A1(\shift_storage.storage[1284] ),
    .S(net747),
    .X(_03605_));
 sg13g2_and2_1 _09291_ (.A(net456),
    .B(_03605_),
    .X(_00419_));
 sg13g2_mux2_1 _09292_ (.A0(\shift_storage.storage[1286] ),
    .A1(\shift_storage.storage[1285] ),
    .S(net747),
    .X(_03606_));
 sg13g2_and2_1 _09293_ (.A(net457),
    .B(_03606_),
    .X(_00420_));
 sg13g2_mux2_1 _09294_ (.A0(\shift_storage.storage[1287] ),
    .A1(\shift_storage.storage[1286] ),
    .S(net749),
    .X(_03607_));
 sg13g2_and2_1 _09295_ (.A(net459),
    .B(_03607_),
    .X(_00421_));
 sg13g2_mux2_1 _09296_ (.A0(\shift_storage.storage[1288] ),
    .A1(\shift_storage.storage[1287] ),
    .S(net746),
    .X(_03608_));
 sg13g2_and2_1 _09297_ (.A(net459),
    .B(_03608_),
    .X(_00422_));
 sg13g2_buf_1 fanout302 (.A(net304),
    .X(net302));
 sg13g2_mux2_1 _09299_ (.A0(\shift_storage.storage[1289] ),
    .A1(\shift_storage.storage[1288] ),
    .S(net749),
    .X(_03610_));
 sg13g2_and2_1 _09300_ (.A(net455),
    .B(_03610_),
    .X(_00423_));
 sg13g2_mux2_1 _09301_ (.A0(\shift_storage.storage[128] ),
    .A1(\shift_storage.storage[127] ),
    .S(net583),
    .X(_03611_));
 sg13g2_and2_1 _09302_ (.A(net287),
    .B(_03611_),
    .X(_00424_));
 sg13g2_mux2_1 _09303_ (.A0(\shift_storage.storage[1290] ),
    .A1(\shift_storage.storage[1289] ),
    .S(net749),
    .X(_03612_));
 sg13g2_and2_1 _09304_ (.A(net457),
    .B(_03612_),
    .X(_00425_));
 sg13g2_buf_2 fanout301 (.A(net305),
    .X(net301));
 sg13g2_mux2_1 _09306_ (.A0(\shift_storage.storage[1291] ),
    .A1(\shift_storage.storage[1290] ),
    .S(net749),
    .X(_03614_));
 sg13g2_and2_1 _09307_ (.A(net457),
    .B(_03614_),
    .X(_00426_));
 sg13g2_mux2_1 _09308_ (.A0(\shift_storage.storage[1292] ),
    .A1(\shift_storage.storage[1291] ),
    .S(net749),
    .X(_03615_));
 sg13g2_and2_1 _09309_ (.A(net457),
    .B(_03615_),
    .X(_00427_));
 sg13g2_mux2_1 _09310_ (.A0(\shift_storage.storage[1293] ),
    .A1(\shift_storage.storage[1292] ),
    .S(net752),
    .X(_03616_));
 sg13g2_and2_1 _09311_ (.A(net462),
    .B(_03616_),
    .X(_00428_));
 sg13g2_mux2_1 _09312_ (.A0(\shift_storage.storage[1294] ),
    .A1(\shift_storage.storage[1293] ),
    .S(net752),
    .X(_03617_));
 sg13g2_and2_1 _09313_ (.A(net462),
    .B(_03617_),
    .X(_00429_));
 sg13g2_mux2_1 _09314_ (.A0(\shift_storage.storage[1295] ),
    .A1(\shift_storage.storage[1294] ),
    .S(net752),
    .X(_03618_));
 sg13g2_and2_1 _09315_ (.A(net462),
    .B(_03618_),
    .X(_00430_));
 sg13g2_mux2_1 _09316_ (.A0(\shift_storage.storage[1296] ),
    .A1(\shift_storage.storage[1295] ),
    .S(net752),
    .X(_03619_));
 sg13g2_and2_1 _09317_ (.A(net462),
    .B(_03619_),
    .X(_00431_));
 sg13g2_mux2_1 _09318_ (.A0(\shift_storage.storage[1297] ),
    .A1(\shift_storage.storage[1296] ),
    .S(net752),
    .X(_03620_));
 sg13g2_and2_1 _09319_ (.A(net460),
    .B(_03620_),
    .X(_00432_));
 sg13g2_buf_2 fanout300 (.A(net301),
    .X(net300));
 sg13g2_mux2_1 _09321_ (.A0(\shift_storage.storage[1298] ),
    .A1(\shift_storage.storage[1297] ),
    .S(net750),
    .X(_03622_));
 sg13g2_and2_1 _09322_ (.A(net460),
    .B(_03622_),
    .X(_00433_));
 sg13g2_mux2_1 _09323_ (.A0(\shift_storage.storage[1299] ),
    .A1(\shift_storage.storage[1298] ),
    .S(net750),
    .X(_03623_));
 sg13g2_and2_1 _09324_ (.A(net460),
    .B(_03623_),
    .X(_00434_));
 sg13g2_mux2_1 _09325_ (.A0(\shift_storage.storage[129] ),
    .A1(\shift_storage.storage[128] ),
    .S(net582),
    .X(_03624_));
 sg13g2_and2_1 _09326_ (.A(net282),
    .B(_03624_),
    .X(_00435_));
 sg13g2_buf_1 fanout299 (.A(net309),
    .X(net299));
 sg13g2_mux2_1 _09328_ (.A0(\shift_storage.storage[12] ),
    .A1(\shift_storage.storage[11] ),
    .S(net610),
    .X(_03626_));
 sg13g2_and2_1 _09329_ (.A(net311),
    .B(_03626_),
    .X(_00436_));
 sg13g2_mux2_1 _09330_ (.A0(\shift_storage.storage[1300] ),
    .A1(\shift_storage.storage[1299] ),
    .S(net750),
    .X(_03627_));
 sg13g2_and2_1 _09331_ (.A(net460),
    .B(_03627_),
    .X(_00437_));
 sg13g2_mux2_1 _09332_ (.A0(\shift_storage.storage[1301] ),
    .A1(\shift_storage.storage[1300] ),
    .S(net750),
    .X(_03628_));
 sg13g2_and2_1 _09333_ (.A(net460),
    .B(_03628_),
    .X(_00438_));
 sg13g2_mux2_1 _09334_ (.A0(\shift_storage.storage[1302] ),
    .A1(\shift_storage.storage[1301] ),
    .S(net750),
    .X(_03629_));
 sg13g2_and2_1 _09335_ (.A(net460),
    .B(_03629_),
    .X(_00439_));
 sg13g2_mux2_1 _09336_ (.A0(\shift_storage.storage[1303] ),
    .A1(\shift_storage.storage[1302] ),
    .S(net750),
    .X(_03630_));
 sg13g2_and2_1 _09337_ (.A(net460),
    .B(_03630_),
    .X(_00440_));
 sg13g2_mux2_1 _09338_ (.A0(\shift_storage.storage[1304] ),
    .A1(\shift_storage.storage[1303] ),
    .S(net750),
    .X(_03631_));
 sg13g2_and2_1 _09339_ (.A(net460),
    .B(_03631_),
    .X(_00441_));
 sg13g2_mux2_1 _09340_ (.A0(\shift_storage.storage[1305] ),
    .A1(\shift_storage.storage[1304] ),
    .S(net751),
    .X(_03632_));
 sg13g2_and2_1 _09341_ (.A(net461),
    .B(_03632_),
    .X(_00442_));
 sg13g2_buf_1 fanout298 (.A(net299),
    .X(net298));
 sg13g2_mux2_1 _09343_ (.A0(\shift_storage.storage[1306] ),
    .A1(\shift_storage.storage[1305] ),
    .S(net750),
    .X(_03634_));
 sg13g2_and2_1 _09344_ (.A(net461),
    .B(_03634_),
    .X(_00443_));
 sg13g2_mux2_1 _09345_ (.A0(\shift_storage.storage[1307] ),
    .A1(\shift_storage.storage[1306] ),
    .S(net751),
    .X(_03635_));
 sg13g2_and2_1 _09346_ (.A(net461),
    .B(_03635_),
    .X(_00444_));
 sg13g2_mux2_1 _09347_ (.A0(\shift_storage.storage[1308] ),
    .A1(\shift_storage.storage[1307] ),
    .S(net751),
    .X(_03636_));
 sg13g2_and2_1 _09348_ (.A(net461),
    .B(_03636_),
    .X(_00445_));
 sg13g2_buf_2 fanout297 (.A(net298),
    .X(net297));
 sg13g2_mux2_1 _09350_ (.A0(\shift_storage.storage[1309] ),
    .A1(\shift_storage.storage[1308] ),
    .S(net753),
    .X(_03638_));
 sg13g2_and2_1 _09351_ (.A(net463),
    .B(_03638_),
    .X(_00446_));
 sg13g2_mux2_1 _09352_ (.A0(\shift_storage.storage[130] ),
    .A1(\shift_storage.storage[129] ),
    .S(net582),
    .X(_03639_));
 sg13g2_and2_1 _09353_ (.A(net282),
    .B(_03639_),
    .X(_00447_));
 sg13g2_mux2_1 _09354_ (.A0(\shift_storage.storage[1310] ),
    .A1(\shift_storage.storage[1309] ),
    .S(net753),
    .X(_03640_));
 sg13g2_and2_1 _09355_ (.A(net463),
    .B(_03640_),
    .X(_00448_));
 sg13g2_mux2_1 _09356_ (.A0(\shift_storage.storage[1311] ),
    .A1(\shift_storage.storage[1310] ),
    .S(net753),
    .X(_03641_));
 sg13g2_and2_1 _09357_ (.A(net464),
    .B(_03641_),
    .X(_00449_));
 sg13g2_mux2_1 _09358_ (.A0(\shift_storage.storage[1312] ),
    .A1(\shift_storage.storage[1311] ),
    .S(net753),
    .X(_03642_));
 sg13g2_and2_1 _09359_ (.A(net463),
    .B(_03642_),
    .X(_00450_));
 sg13g2_mux2_1 _09360_ (.A0(\shift_storage.storage[1313] ),
    .A1(\shift_storage.storage[1312] ),
    .S(net753),
    .X(_03643_));
 sg13g2_and2_1 _09361_ (.A(net463),
    .B(_03643_),
    .X(_00451_));
 sg13g2_mux2_1 _09362_ (.A0(\shift_storage.storage[1314] ),
    .A1(\shift_storage.storage[1313] ),
    .S(net755),
    .X(_03644_));
 sg13g2_and2_1 _09363_ (.A(net465),
    .B(_03644_),
    .X(_00452_));
 sg13g2_buf_1 fanout296 (.A(net299),
    .X(net296));
 sg13g2_buf_1 fanout295 (.A(net299),
    .X(net295));
 sg13g2_mux2_1 _09366_ (.A0(\shift_storage.storage[1315] ),
    .A1(\shift_storage.storage[1314] ),
    .S(net755),
    .X(_03647_));
 sg13g2_and2_1 _09367_ (.A(net465),
    .B(_03647_),
    .X(_00453_));
 sg13g2_mux2_1 _09368_ (.A0(\shift_storage.storage[1316] ),
    .A1(\shift_storage.storage[1315] ),
    .S(net755),
    .X(_03648_));
 sg13g2_and2_1 _09369_ (.A(net465),
    .B(_03648_),
    .X(_00454_));
 sg13g2_mux2_1 _09370_ (.A0(\shift_storage.storage[1317] ),
    .A1(\shift_storage.storage[1316] ),
    .S(net756),
    .X(_03649_));
 sg13g2_and2_1 _09371_ (.A(net468),
    .B(_03649_),
    .X(_00455_));
 sg13g2_buf_1 fanout294 (.A(net299),
    .X(net294));
 sg13g2_buf_1 fanout293 (.A(net294),
    .X(net293));
 sg13g2_mux2_1 _09374_ (.A0(\shift_storage.storage[1318] ),
    .A1(\shift_storage.storage[1317] ),
    .S(net756),
    .X(_03652_));
 sg13g2_and2_1 _09375_ (.A(net468),
    .B(_03652_),
    .X(_00456_));
 sg13g2_mux2_1 _09376_ (.A0(\shift_storage.storage[1319] ),
    .A1(\shift_storage.storage[1318] ),
    .S(net756),
    .X(_03653_));
 sg13g2_and2_1 _09377_ (.A(net468),
    .B(_03653_),
    .X(_00457_));
 sg13g2_mux2_1 _09378_ (.A0(\shift_storage.storage[131] ),
    .A1(\shift_storage.storage[130] ),
    .S(net575),
    .X(_03654_));
 sg13g2_and2_1 _09379_ (.A(net275),
    .B(_03654_),
    .X(_00458_));
 sg13g2_mux2_1 _09380_ (.A0(\shift_storage.storage[1320] ),
    .A1(\shift_storage.storage[1319] ),
    .S(net768),
    .X(_03655_));
 sg13g2_and2_1 _09381_ (.A(net485),
    .B(_03655_),
    .X(_00459_));
 sg13g2_mux2_1 _09382_ (.A0(\shift_storage.storage[1321] ),
    .A1(\shift_storage.storage[1320] ),
    .S(net768),
    .X(_03656_));
 sg13g2_and2_1 _09383_ (.A(net484),
    .B(_03656_),
    .X(_00460_));
 sg13g2_mux2_1 _09384_ (.A0(\shift_storage.storage[1322] ),
    .A1(\shift_storage.storage[1321] ),
    .S(net768),
    .X(_03657_));
 sg13g2_and2_1 _09385_ (.A(net484),
    .B(_03657_),
    .X(_00461_));
 sg13g2_mux2_1 _09386_ (.A0(\shift_storage.storage[1323] ),
    .A1(\shift_storage.storage[1322] ),
    .S(net768),
    .X(_03658_));
 sg13g2_and2_1 _09387_ (.A(net484),
    .B(_03658_),
    .X(_00462_));
 sg13g2_buf_2 fanout292 (.A(net294),
    .X(net292));
 sg13g2_mux2_1 _09389_ (.A0(\shift_storage.storage[1324] ),
    .A1(\shift_storage.storage[1323] ),
    .S(net768),
    .X(_03660_));
 sg13g2_and2_1 _09390_ (.A(net485),
    .B(_03660_),
    .X(_00463_));
 sg13g2_mux2_1 _09391_ (.A0(\shift_storage.storage[1325] ),
    .A1(\shift_storage.storage[1324] ),
    .S(net768),
    .X(_03661_));
 sg13g2_and2_1 _09392_ (.A(net485),
    .B(_03661_),
    .X(_00464_));
 sg13g2_mux2_1 _09393_ (.A0(\shift_storage.storage[1326] ),
    .A1(\shift_storage.storage[1325] ),
    .S(net773),
    .X(_03662_));
 sg13g2_and2_1 _09394_ (.A(net485),
    .B(_03662_),
    .X(_00465_));
 sg13g2_buf_1 fanout291 (.A(net294),
    .X(net291));
 sg13g2_mux2_1 _09396_ (.A0(\shift_storage.storage[1327] ),
    .A1(\shift_storage.storage[1326] ),
    .S(net771),
    .X(_03664_));
 sg13g2_and2_1 _09397_ (.A(net490),
    .B(_03664_),
    .X(_00466_));
 sg13g2_mux2_1 _09398_ (.A0(\shift_storage.storage[1328] ),
    .A1(\shift_storage.storage[1327] ),
    .S(net771),
    .X(_03665_));
 sg13g2_and2_1 _09399_ (.A(net490),
    .B(_03665_),
    .X(_00467_));
 sg13g2_mux2_1 _09400_ (.A0(\shift_storage.storage[1329] ),
    .A1(\shift_storage.storage[1328] ),
    .S(net771),
    .X(_03666_));
 sg13g2_and2_1 _09401_ (.A(net490),
    .B(_03666_),
    .X(_00468_));
 sg13g2_mux2_1 _09402_ (.A0(\shift_storage.storage[132] ),
    .A1(\shift_storage.storage[131] ),
    .S(net574),
    .X(_03667_));
 sg13g2_and2_1 _09403_ (.A(net274),
    .B(_03667_),
    .X(_00469_));
 sg13g2_mux2_1 _09404_ (.A0(\shift_storage.storage[1330] ),
    .A1(\shift_storage.storage[1329] ),
    .S(net771),
    .X(_03668_));
 sg13g2_and2_1 _09405_ (.A(net490),
    .B(_03668_),
    .X(_00470_));
 sg13g2_mux2_1 _09406_ (.A0(\shift_storage.storage[1331] ),
    .A1(\shift_storage.storage[1330] ),
    .S(net769),
    .X(_03669_));
 sg13g2_and2_1 _09407_ (.A(net488),
    .B(_03669_),
    .X(_00471_));
 sg13g2_mux2_1 _09408_ (.A0(\shift_storage.storage[1332] ),
    .A1(\shift_storage.storage[1331] ),
    .S(net769),
    .X(_03670_));
 sg13g2_and2_1 _09409_ (.A(net488),
    .B(_03670_),
    .X(_00472_));
 sg13g2_buf_2 fanout290 (.A(net294),
    .X(net290));
 sg13g2_mux2_1 _09411_ (.A0(\shift_storage.storage[1333] ),
    .A1(\shift_storage.storage[1332] ),
    .S(net769),
    .X(_03672_));
 sg13g2_and2_1 _09412_ (.A(net488),
    .B(_03672_),
    .X(_00473_));
 sg13g2_mux2_1 _09413_ (.A0(\shift_storage.storage[1334] ),
    .A1(\shift_storage.storage[1333] ),
    .S(net770),
    .X(_03673_));
 sg13g2_and2_1 _09414_ (.A(net489),
    .B(_03673_),
    .X(_00474_));
 sg13g2_mux2_1 _09415_ (.A0(\shift_storage.storage[1335] ),
    .A1(\shift_storage.storage[1334] ),
    .S(net770),
    .X(_03674_));
 sg13g2_and2_1 _09416_ (.A(net489),
    .B(_03674_),
    .X(_00475_));
 sg13g2_buf_1 fanout289 (.A(net356),
    .X(net289));
 sg13g2_mux2_1 _09418_ (.A0(\shift_storage.storage[1336] ),
    .A1(\shift_storage.storage[1335] ),
    .S(net770),
    .X(_03676_));
 sg13g2_and2_1 _09419_ (.A(net489),
    .B(_03676_),
    .X(_00476_));
 sg13g2_mux2_1 _09420_ (.A0(\shift_storage.storage[1337] ),
    .A1(\shift_storage.storage[1336] ),
    .S(net769),
    .X(_03677_));
 sg13g2_and2_1 _09421_ (.A(net488),
    .B(_03677_),
    .X(_00477_));
 sg13g2_mux2_1 _09422_ (.A0(\shift_storage.storage[1338] ),
    .A1(\shift_storage.storage[1337] ),
    .S(net769),
    .X(_03678_));
 sg13g2_and2_1 _09423_ (.A(net488),
    .B(_03678_),
    .X(_00478_));
 sg13g2_mux2_1 _09424_ (.A0(\shift_storage.storage[1339] ),
    .A1(\shift_storage.storage[1338] ),
    .S(net769),
    .X(_03679_));
 sg13g2_and2_1 _09425_ (.A(net488),
    .B(_03679_),
    .X(_00479_));
 sg13g2_mux2_1 _09426_ (.A0(\shift_storage.storage[133] ),
    .A1(\shift_storage.storage[132] ),
    .S(net576),
    .X(_03680_));
 sg13g2_and2_1 _09427_ (.A(net276),
    .B(_03680_),
    .X(_00480_));
 sg13g2_mux2_1 _09428_ (.A0(\shift_storage.storage[1340] ),
    .A1(\shift_storage.storage[1339] ),
    .S(net769),
    .X(_03681_));
 sg13g2_and2_1 _09429_ (.A(net488),
    .B(_03681_),
    .X(_00481_));
 sg13g2_mux2_1 _09430_ (.A0(\shift_storage.storage[1341] ),
    .A1(\shift_storage.storage[1340] ),
    .S(net771),
    .X(_03682_));
 sg13g2_and2_1 _09431_ (.A(net490),
    .B(_03682_),
    .X(_00482_));
 sg13g2_buf_1 fanout288 (.A(net289),
    .X(net288));
 sg13g2_mux2_1 _09433_ (.A0(\shift_storage.storage[1342] ),
    .A1(\shift_storage.storage[1341] ),
    .S(net771),
    .X(_03684_));
 sg13g2_and2_1 _09434_ (.A(net490),
    .B(_03684_),
    .X(_00483_));
 sg13g2_mux2_1 _09435_ (.A0(\shift_storage.storage[1343] ),
    .A1(\shift_storage.storage[1342] ),
    .S(net771),
    .X(_03685_));
 sg13g2_and2_1 _09436_ (.A(net490),
    .B(_03685_),
    .X(_00484_));
 sg13g2_mux2_1 _09437_ (.A0(\shift_storage.storage[1344] ),
    .A1(\shift_storage.storage[1343] ),
    .S(net771),
    .X(_03686_));
 sg13g2_and2_1 _09438_ (.A(net490),
    .B(_03686_),
    .X(_00485_));
 sg13g2_buf_1 fanout287 (.A(net288),
    .X(net287));
 sg13g2_mux2_1 _09440_ (.A0(\shift_storage.storage[1345] ),
    .A1(\shift_storage.storage[1344] ),
    .S(net768),
    .X(_03688_));
 sg13g2_and2_1 _09441_ (.A(net486),
    .B(_03688_),
    .X(_00486_));
 sg13g2_mux2_1 _09442_ (.A0(\shift_storage.storage[1346] ),
    .A1(\shift_storage.storage[1345] ),
    .S(net768),
    .X(_03689_));
 sg13g2_and2_1 _09443_ (.A(net484),
    .B(_03689_),
    .X(_00487_));
 sg13g2_mux2_1 _09444_ (.A0(\shift_storage.storage[1347] ),
    .A1(\shift_storage.storage[1346] ),
    .S(net755),
    .X(_03690_));
 sg13g2_and2_1 _09445_ (.A(net468),
    .B(_03690_),
    .X(_00488_));
 sg13g2_mux2_1 _09446_ (.A0(\shift_storage.storage[1348] ),
    .A1(\shift_storage.storage[1347] ),
    .S(net755),
    .X(_03691_));
 sg13g2_and2_1 _09447_ (.A(net466),
    .B(_03691_),
    .X(_00489_));
 sg13g2_mux2_1 _09448_ (.A0(\shift_storage.storage[1349] ),
    .A1(\shift_storage.storage[1348] ),
    .S(net755),
    .X(_03692_));
 sg13g2_and2_1 _09449_ (.A(net465),
    .B(_03692_),
    .X(_00490_));
 sg13g2_mux2_1 _09450_ (.A0(\shift_storage.storage[134] ),
    .A1(\shift_storage.storage[133] ),
    .S(net576),
    .X(_03693_));
 sg13g2_and2_1 _09451_ (.A(net274),
    .B(_03693_),
    .X(_00491_));
 sg13g2_mux2_1 _09452_ (.A0(\shift_storage.storage[1350] ),
    .A1(\shift_storage.storage[1349] ),
    .S(net755),
    .X(_03694_));
 sg13g2_and2_1 _09453_ (.A(net465),
    .B(_03694_),
    .X(_00492_));
 sg13g2_buf_1 fanout286 (.A(net287),
    .X(net286));
 sg13g2_mux2_1 _09455_ (.A0(\shift_storage.storage[1351] ),
    .A1(\shift_storage.storage[1350] ),
    .S(net755),
    .X(_03696_));
 sg13g2_and2_1 _09456_ (.A(net465),
    .B(_03696_),
    .X(_00493_));
 sg13g2_mux2_1 _09457_ (.A0(\shift_storage.storage[1352] ),
    .A1(\shift_storage.storage[1351] ),
    .S(net753),
    .X(_03697_));
 sg13g2_and2_1 _09458_ (.A(net463),
    .B(_03697_),
    .X(_00494_));
 sg13g2_mux2_1 _09459_ (.A0(\shift_storage.storage[1353] ),
    .A1(\shift_storage.storage[1352] ),
    .S(net753),
    .X(_03698_));
 sg13g2_and2_1 _09460_ (.A(net463),
    .B(_03698_),
    .X(_00495_));
 sg13g2_buf_2 fanout285 (.A(net286),
    .X(net285));
 sg13g2_mux2_1 _09462_ (.A0(\shift_storage.storage[1354] ),
    .A1(\shift_storage.storage[1353] ),
    .S(net754),
    .X(_03700_));
 sg13g2_and2_1 _09463_ (.A(net464),
    .B(_03700_),
    .X(_00496_));
 sg13g2_mux2_1 _09464_ (.A0(\shift_storage.storage[1355] ),
    .A1(\shift_storage.storage[1354] ),
    .S(net753),
    .X(_03701_));
 sg13g2_and2_1 _09465_ (.A(net462),
    .B(_03701_),
    .X(_00497_));
 sg13g2_mux2_1 _09466_ (.A0(\shift_storage.storage[1356] ),
    .A1(\shift_storage.storage[1355] ),
    .S(net752),
    .X(_03702_));
 sg13g2_and2_1 _09467_ (.A(net463),
    .B(_03702_),
    .X(_00498_));
 sg13g2_mux2_1 _09468_ (.A0(\shift_storage.storage[1357] ),
    .A1(\shift_storage.storage[1356] ),
    .S(net754),
    .X(_03703_));
 sg13g2_and2_1 _09469_ (.A(net462),
    .B(_03703_),
    .X(_00499_));
 sg13g2_mux2_1 _09470_ (.A0(\shift_storage.storage[1358] ),
    .A1(\shift_storage.storage[1357] ),
    .S(net752),
    .X(_03704_));
 sg13g2_and2_1 _09471_ (.A(net462),
    .B(_03704_),
    .X(_00500_));
 sg13g2_mux2_1 _09472_ (.A0(\shift_storage.storage[1359] ),
    .A1(\shift_storage.storage[1358] ),
    .S(net752),
    .X(_03705_));
 sg13g2_and2_1 _09473_ (.A(net462),
    .B(_03705_),
    .X(_00501_));
 sg13g2_mux2_1 _09474_ (.A0(\shift_storage.storage[135] ),
    .A1(\shift_storage.storage[134] ),
    .S(net574),
    .X(_03706_));
 sg13g2_and2_1 _09475_ (.A(net274),
    .B(_03706_),
    .X(_00502_));
 sg13g2_buf_2 fanout284 (.A(net286),
    .X(net284));
 sg13g2_mux2_1 _09477_ (.A0(\shift_storage.storage[1360] ),
    .A1(\shift_storage.storage[1359] ),
    .S(net748),
    .X(_03708_));
 sg13g2_and2_1 _09478_ (.A(net458),
    .B(_03708_),
    .X(_00503_));
 sg13g2_mux2_1 _09479_ (.A0(\shift_storage.storage[1361] ),
    .A1(\shift_storage.storage[1360] ),
    .S(net748),
    .X(_03709_));
 sg13g2_and2_1 _09480_ (.A(net457),
    .B(_03709_),
    .X(_00504_));
 sg13g2_mux2_1 _09481_ (.A0(\shift_storage.storage[1362] ),
    .A1(\shift_storage.storage[1361] ),
    .S(net748),
    .X(_03710_));
 sg13g2_and2_1 _09482_ (.A(net457),
    .B(_03710_),
    .X(_00505_));
 sg13g2_buf_2 fanout283 (.A(net287),
    .X(net283));
 sg13g2_mux2_1 _09484_ (.A0(\shift_storage.storage[1363] ),
    .A1(\shift_storage.storage[1362] ),
    .S(net748),
    .X(_03712_));
 sg13g2_and2_1 _09485_ (.A(net457),
    .B(_03712_),
    .X(_00506_));
 sg13g2_mux2_1 _09486_ (.A0(\shift_storage.storage[1364] ),
    .A1(\shift_storage.storage[1363] ),
    .S(net748),
    .X(_03713_));
 sg13g2_and2_1 _09487_ (.A(net457),
    .B(_03713_),
    .X(_00507_));
 sg13g2_mux2_1 _09488_ (.A0(\shift_storage.storage[1365] ),
    .A1(\shift_storage.storage[1364] ),
    .S(net748),
    .X(_03714_));
 sg13g2_and2_1 _09489_ (.A(net456),
    .B(_03714_),
    .X(_00508_));
 sg13g2_mux2_1 _09490_ (.A0(\shift_storage.storage[1366] ),
    .A1(\shift_storage.storage[1365] ),
    .S(net748),
    .X(_03715_));
 sg13g2_and2_1 _09491_ (.A(net456),
    .B(_03715_),
    .X(_00509_));
 sg13g2_mux2_1 _09492_ (.A0(\shift_storage.storage[1367] ),
    .A1(\shift_storage.storage[1366] ),
    .S(net747),
    .X(_03716_));
 sg13g2_and2_1 _09493_ (.A(net456),
    .B(_03716_),
    .X(_00510_));
 sg13g2_mux2_1 _09494_ (.A0(\shift_storage.storage[1368] ),
    .A1(\shift_storage.storage[1367] ),
    .S(net747),
    .X(_03717_));
 sg13g2_and2_1 _09495_ (.A(net456),
    .B(_03717_),
    .X(_00511_));
 sg13g2_mux2_1 _09496_ (.A0(\shift_storage.storage[1369] ),
    .A1(\shift_storage.storage[1368] ),
    .S(net747),
    .X(_03718_));
 sg13g2_and2_1 _09497_ (.A(net458),
    .B(_03718_),
    .X(_00512_));
 sg13g2_buf_2 fanout282 (.A(net283),
    .X(net282));
 sg13g2_mux2_1 _09499_ (.A0(\shift_storage.storage[136] ),
    .A1(\shift_storage.storage[135] ),
    .S(net574),
    .X(_03720_));
 sg13g2_and2_1 _09500_ (.A(net274),
    .B(_03720_),
    .X(_00513_));
 sg13g2_mux2_1 _09501_ (.A0(\shift_storage.storage[1370] ),
    .A1(\shift_storage.storage[1369] ),
    .S(net738),
    .X(_03721_));
 sg13g2_and2_1 _09502_ (.A(net444),
    .B(_03721_),
    .X(_00514_));
 sg13g2_mux2_1 _09503_ (.A0(\shift_storage.storage[1371] ),
    .A1(\shift_storage.storage[1370] ),
    .S(net738),
    .X(_03722_));
 sg13g2_and2_1 _09504_ (.A(net444),
    .B(_03722_),
    .X(_00515_));
 sg13g2_buf_1 fanout281 (.A(net288),
    .X(net281));
 sg13g2_mux2_1 _09506_ (.A0(\shift_storage.storage[1372] ),
    .A1(\shift_storage.storage[1371] ),
    .S(net738),
    .X(_03724_));
 sg13g2_and2_1 _09507_ (.A(net445),
    .B(_03724_),
    .X(_00516_));
 sg13g2_mux2_1 _09508_ (.A0(\shift_storage.storage[1373] ),
    .A1(\shift_storage.storage[1372] ),
    .S(net738),
    .X(_03725_));
 sg13g2_and2_1 _09509_ (.A(net444),
    .B(_03725_),
    .X(_00517_));
 sg13g2_mux2_1 _09510_ (.A0(\shift_storage.storage[1374] ),
    .A1(\shift_storage.storage[1373] ),
    .S(net738),
    .X(_03726_));
 sg13g2_and2_1 _09511_ (.A(net444),
    .B(_03726_),
    .X(_00518_));
 sg13g2_mux2_1 _09512_ (.A0(\shift_storage.storage[1375] ),
    .A1(\shift_storage.storage[1374] ),
    .S(net737),
    .X(_03727_));
 sg13g2_and2_1 _09513_ (.A(net443),
    .B(_03727_),
    .X(_00519_));
 sg13g2_mux2_1 _09514_ (.A0(\shift_storage.storage[1376] ),
    .A1(\shift_storage.storage[1375] ),
    .S(net745),
    .X(_03728_));
 sg13g2_and2_1 _09515_ (.A(net451),
    .B(_03728_),
    .X(_00520_));
 sg13g2_mux2_1 _09516_ (.A0(\shift_storage.storage[1377] ),
    .A1(\shift_storage.storage[1376] ),
    .S(net745),
    .X(_03729_));
 sg13g2_and2_1 _09517_ (.A(net451),
    .B(_03729_),
    .X(_00521_));
 sg13g2_mux2_1 _09518_ (.A0(\shift_storage.storage[1378] ),
    .A1(\shift_storage.storage[1377] ),
    .S(net745),
    .X(_03730_));
 sg13g2_and2_1 _09519_ (.A(net451),
    .B(_03730_),
    .X(_00522_));
 sg13g2_buf_1 fanout280 (.A(net281),
    .X(net280));
 sg13g2_buf_1 fanout279 (.A(net280),
    .X(net279));
 sg13g2_mux2_1 _09522_ (.A0(\shift_storage.storage[1379] ),
    .A1(\shift_storage.storage[1378] ),
    .S(net745),
    .X(_03733_));
 sg13g2_and2_1 _09523_ (.A(net451),
    .B(_03733_),
    .X(_00523_));
 sg13g2_mux2_1 _09524_ (.A0(\shift_storage.storage[137] ),
    .A1(\shift_storage.storage[136] ),
    .S(net574),
    .X(_03734_));
 sg13g2_and2_1 _09525_ (.A(net274),
    .B(_03734_),
    .X(_00524_));
 sg13g2_mux2_1 _09526_ (.A0(\shift_storage.storage[1380] ),
    .A1(\shift_storage.storage[1379] ),
    .S(net745),
    .X(_03735_));
 sg13g2_and2_1 _09527_ (.A(net451),
    .B(_03735_),
    .X(_00525_));
 sg13g2_buf_1 fanout278 (.A(net281),
    .X(net278));
 sg13g2_buf_2 fanout277 (.A(net281),
    .X(net277));
 sg13g2_mux2_1 _09530_ (.A0(\shift_storage.storage[1381] ),
    .A1(\shift_storage.storage[1380] ),
    .S(net745),
    .X(_03738_));
 sg13g2_and2_1 _09531_ (.A(net452),
    .B(_03738_),
    .X(_00526_));
 sg13g2_mux2_1 _09532_ (.A0(\shift_storage.storage[1382] ),
    .A1(\shift_storage.storage[1381] ),
    .S(net745),
    .X(_03739_));
 sg13g2_and2_1 _09533_ (.A(net452),
    .B(_03739_),
    .X(_00527_));
 sg13g2_mux2_1 _09534_ (.A0(\shift_storage.storage[1383] ),
    .A1(\shift_storage.storage[1382] ),
    .S(net743),
    .X(_03740_));
 sg13g2_and2_1 _09535_ (.A(net450),
    .B(_03740_),
    .X(_00528_));
 sg13g2_mux2_1 _09536_ (.A0(\shift_storage.storage[1384] ),
    .A1(\shift_storage.storage[1383] ),
    .S(net743),
    .X(_03741_));
 sg13g2_and2_1 _09537_ (.A(net450),
    .B(_03741_),
    .X(_00529_));
 sg13g2_mux2_1 _09538_ (.A0(\shift_storage.storage[1385] ),
    .A1(\shift_storage.storage[1384] ),
    .S(net744),
    .X(_03742_));
 sg13g2_and2_1 _09539_ (.A(net447),
    .B(_03742_),
    .X(_00530_));
 sg13g2_mux2_1 _09540_ (.A0(\shift_storage.storage[1386] ),
    .A1(\shift_storage.storage[1385] ),
    .S(net740),
    .X(_03743_));
 sg13g2_and2_1 _09541_ (.A(net447),
    .B(_03743_),
    .X(_00531_));
 sg13g2_mux2_1 _09542_ (.A0(\shift_storage.storage[1387] ),
    .A1(\shift_storage.storage[1386] ),
    .S(net740),
    .X(_03744_));
 sg13g2_and2_1 _09543_ (.A(net447),
    .B(_03744_),
    .X(_00532_));
 sg13g2_buf_1 fanout276 (.A(net288),
    .X(net276));
 sg13g2_mux2_1 _09545_ (.A0(\shift_storage.storage[1388] ),
    .A1(\shift_storage.storage[1387] ),
    .S(net740),
    .X(_03746_));
 sg13g2_and2_1 _09546_ (.A(net447),
    .B(_03746_),
    .X(_00533_));
 sg13g2_mux2_1 _09547_ (.A0(\shift_storage.storage[1389] ),
    .A1(\shift_storage.storage[1388] ),
    .S(net731),
    .X(_03747_));
 sg13g2_and2_1 _09548_ (.A(net437),
    .B(_03747_),
    .X(_00534_));
 sg13g2_mux2_1 _09549_ (.A0(\shift_storage.storage[138] ),
    .A1(\shift_storage.storage[137] ),
    .S(net575),
    .X(_03748_));
 sg13g2_and2_1 _09550_ (.A(net275),
    .B(_03748_),
    .X(_00535_));
 sg13g2_buf_2 fanout275 (.A(net276),
    .X(net275));
 sg13g2_mux2_1 _09552_ (.A0(\shift_storage.storage[1390] ),
    .A1(\shift_storage.storage[1389] ),
    .S(net731),
    .X(_03750_));
 sg13g2_and2_1 _09553_ (.A(net443),
    .B(_03750_),
    .X(_00536_));
 sg13g2_mux2_1 _09554_ (.A0(\shift_storage.storage[1391] ),
    .A1(\shift_storage.storage[1390] ),
    .S(net737),
    .X(_03751_));
 sg13g2_and2_1 _09555_ (.A(net443),
    .B(_03751_),
    .X(_00537_));
 sg13g2_mux2_1 _09556_ (.A0(\shift_storage.storage[1392] ),
    .A1(\shift_storage.storage[1391] ),
    .S(net737),
    .X(_03752_));
 sg13g2_and2_1 _09557_ (.A(net443),
    .B(_03752_),
    .X(_00538_));
 sg13g2_mux2_1 _09558_ (.A0(\shift_storage.storage[1393] ),
    .A1(\shift_storage.storage[1392] ),
    .S(net737),
    .X(_03753_));
 sg13g2_and2_1 _09559_ (.A(net444),
    .B(_03753_),
    .X(_00539_));
 sg13g2_mux2_1 _09560_ (.A0(\shift_storage.storage[1394] ),
    .A1(\shift_storage.storage[1393] ),
    .S(net737),
    .X(_03754_));
 sg13g2_and2_1 _09561_ (.A(net443),
    .B(_03754_),
    .X(_00540_));
 sg13g2_mux2_1 _09562_ (.A0(\shift_storage.storage[1395] ),
    .A1(\shift_storage.storage[1394] ),
    .S(net737),
    .X(_03755_));
 sg13g2_and2_1 _09563_ (.A(net443),
    .B(_03755_),
    .X(_00541_));
 sg13g2_mux2_1 _09564_ (.A0(\shift_storage.storage[1396] ),
    .A1(\shift_storage.storage[1395] ),
    .S(net738),
    .X(_03756_));
 sg13g2_and2_1 _09565_ (.A(net444),
    .B(_03756_),
    .X(_00542_));
 sg13g2_buf_1 fanout274 (.A(net276),
    .X(net274));
 sg13g2_mux2_1 _09567_ (.A0(\shift_storage.storage[1397] ),
    .A1(\shift_storage.storage[1396] ),
    .S(net738),
    .X(_03758_));
 sg13g2_and2_1 _09568_ (.A(net444),
    .B(_03758_),
    .X(_00543_));
 sg13g2_mux2_1 _09569_ (.A0(\shift_storage.storage[1398] ),
    .A1(\shift_storage.storage[1397] ),
    .S(net735),
    .X(_03759_));
 sg13g2_and2_1 _09570_ (.A(net441),
    .B(_03759_),
    .X(_00544_));
 sg13g2_mux2_1 _09571_ (.A0(\shift_storage.storage[1399] ),
    .A1(\shift_storage.storage[1398] ),
    .S(net736),
    .X(_03760_));
 sg13g2_and2_1 _09572_ (.A(net441),
    .B(_03760_),
    .X(_00545_));
 sg13g2_buf_1 fanout273 (.A(net276),
    .X(net273));
 sg13g2_mux2_1 _09574_ (.A0(\shift_storage.storage[139] ),
    .A1(\shift_storage.storage[138] ),
    .S(net575),
    .X(_03762_));
 sg13g2_and2_1 _09575_ (.A(net275),
    .B(_03762_),
    .X(_00546_));
 sg13g2_mux2_1 _09576_ (.A0(\shift_storage.storage[13] ),
    .A1(\shift_storage.storage[12] ),
    .S(net610),
    .X(_03763_));
 sg13g2_and2_1 _09577_ (.A(net311),
    .B(_03763_),
    .X(_00547_));
 sg13g2_mux2_1 _09578_ (.A0(\shift_storage.storage[1400] ),
    .A1(\shift_storage.storage[1399] ),
    .S(net735),
    .X(_03764_));
 sg13g2_and2_1 _09579_ (.A(net441),
    .B(_03764_),
    .X(_00548_));
 sg13g2_mux2_1 _09580_ (.A0(\shift_storage.storage[1401] ),
    .A1(\shift_storage.storage[1400] ),
    .S(net736),
    .X(_03765_));
 sg13g2_and2_1 _09581_ (.A(net440),
    .B(_03765_),
    .X(_00549_));
 sg13g2_mux2_1 _09582_ (.A0(\shift_storage.storage[1402] ),
    .A1(\shift_storage.storage[1401] ),
    .S(net736),
    .X(_03766_));
 sg13g2_and2_1 _09583_ (.A(net442),
    .B(_03766_),
    .X(_00550_));
 sg13g2_mux2_1 _09584_ (.A0(\shift_storage.storage[1403] ),
    .A1(\shift_storage.storage[1402] ),
    .S(net734),
    .X(_03767_));
 sg13g2_and2_1 _09585_ (.A(net440),
    .B(_03767_),
    .X(_00551_));
 sg13g2_mux2_1 _09586_ (.A0(\shift_storage.storage[1404] ),
    .A1(\shift_storage.storage[1403] ),
    .S(net734),
    .X(_03768_));
 sg13g2_and2_1 _09587_ (.A(net440),
    .B(_03768_),
    .X(_00552_));
 sg13g2_buf_2 fanout272 (.A(net276),
    .X(net272));
 sg13g2_mux2_1 _09589_ (.A0(\shift_storage.storage[1405] ),
    .A1(\shift_storage.storage[1404] ),
    .S(net737),
    .X(_03770_));
 sg13g2_and2_1 _09590_ (.A(net443),
    .B(_03770_),
    .X(_00553_));
 sg13g2_mux2_1 _09591_ (.A0(\shift_storage.storage[1406] ),
    .A1(\shift_storage.storage[1405] ),
    .S(net737),
    .X(_03771_));
 sg13g2_and2_1 _09592_ (.A(net443),
    .B(_03771_),
    .X(_00554_));
 sg13g2_mux2_1 _09593_ (.A0(\shift_storage.storage[1407] ),
    .A1(\shift_storage.storage[1406] ),
    .S(net732),
    .X(_03772_));
 sg13g2_and2_1 _09594_ (.A(net438),
    .B(_03772_),
    .X(_00555_));
 sg13g2_buf_1 fanout271 (.A(net288),
    .X(net271));
 sg13g2_mux2_1 _09596_ (.A0(\shift_storage.storage[1408] ),
    .A1(\shift_storage.storage[1407] ),
    .S(net732),
    .X(_03774_));
 sg13g2_and2_1 _09597_ (.A(net438),
    .B(_03774_),
    .X(_00556_));
 sg13g2_mux2_1 _09598_ (.A0(\shift_storage.storage[1409] ),
    .A1(\shift_storage.storage[1408] ),
    .S(net732),
    .X(_03775_));
 sg13g2_and2_1 _09599_ (.A(net438),
    .B(_03775_),
    .X(_00557_));
 sg13g2_mux2_1 _09600_ (.A0(\shift_storage.storage[140] ),
    .A1(\shift_storage.storage[139] ),
    .S(net572),
    .X(_03776_));
 sg13g2_and2_1 _09601_ (.A(net272),
    .B(_03776_),
    .X(_00558_));
 sg13g2_mux2_1 _09602_ (.A0(\shift_storage.storage[1410] ),
    .A1(\shift_storage.storage[1409] ),
    .S(net732),
    .X(_03777_));
 sg13g2_and2_1 _09603_ (.A(net438),
    .B(_03777_),
    .X(_00559_));
 sg13g2_mux2_1 _09604_ (.A0(\shift_storage.storage[1411] ),
    .A1(\shift_storage.storage[1410] ),
    .S(net732),
    .X(_03778_));
 sg13g2_and2_1 _09605_ (.A(net438),
    .B(_03778_),
    .X(_00560_));
 sg13g2_mux2_1 _09606_ (.A0(\shift_storage.storage[1412] ),
    .A1(\shift_storage.storage[1411] ),
    .S(net732),
    .X(_03779_));
 sg13g2_and2_1 _09607_ (.A(net437),
    .B(_03779_),
    .X(_00561_));
 sg13g2_mux2_1 _09608_ (.A0(\shift_storage.storage[1413] ),
    .A1(\shift_storage.storage[1412] ),
    .S(net731),
    .X(_03780_));
 sg13g2_and2_1 _09609_ (.A(net437),
    .B(_03780_),
    .X(_00562_));
 sg13g2_buf_1 fanout270 (.A(net271),
    .X(net270));
 sg13g2_mux2_1 _09611_ (.A0(\shift_storage.storage[1414] ),
    .A1(\shift_storage.storage[1413] ),
    .S(net730),
    .X(_03782_));
 sg13g2_and2_1 _09612_ (.A(net435),
    .B(_03782_),
    .X(_00563_));
 sg13g2_mux2_1 _09613_ (.A0(\shift_storage.storage[1415] ),
    .A1(\shift_storage.storage[1414] ),
    .S(net730),
    .X(_03783_));
 sg13g2_and2_1 _09614_ (.A(net435),
    .B(_03783_),
    .X(_00564_));
 sg13g2_mux2_1 _09615_ (.A0(\shift_storage.storage[1416] ),
    .A1(\shift_storage.storage[1415] ),
    .S(net730),
    .X(_03784_));
 sg13g2_and2_1 _09616_ (.A(net435),
    .B(_03784_),
    .X(_00565_));
 sg13g2_buf_1 fanout269 (.A(net271),
    .X(net269));
 sg13g2_mux2_1 _09618_ (.A0(\shift_storage.storage[1417] ),
    .A1(\shift_storage.storage[1416] ),
    .S(net730),
    .X(_03786_));
 sg13g2_and2_1 _09619_ (.A(net435),
    .B(_03786_),
    .X(_00566_));
 sg13g2_mux2_1 _09620_ (.A0(\shift_storage.storage[1418] ),
    .A1(\shift_storage.storage[1417] ),
    .S(net633),
    .X(_03787_));
 sg13g2_and2_1 _09621_ (.A(net335),
    .B(_03787_),
    .X(_00567_));
 sg13g2_mux2_1 _09622_ (.A0(\shift_storage.storage[1419] ),
    .A1(\shift_storage.storage[1418] ),
    .S(net633),
    .X(_03788_));
 sg13g2_and2_1 _09623_ (.A(net335),
    .B(_03788_),
    .X(_00568_));
 sg13g2_mux2_1 _09624_ (.A0(\shift_storage.storage[141] ),
    .A1(\shift_storage.storage[140] ),
    .S(net572),
    .X(_03789_));
 sg13g2_and2_1 _09625_ (.A(net272),
    .B(_03789_),
    .X(_00569_));
 sg13g2_mux2_1 _09626_ (.A0(\shift_storage.storage[1420] ),
    .A1(\shift_storage.storage[1419] ),
    .S(net633),
    .X(_03790_));
 sg13g2_and2_1 _09627_ (.A(net335),
    .B(_03790_),
    .X(_00570_));
 sg13g2_mux2_1 _09628_ (.A0(\shift_storage.storage[1421] ),
    .A1(\shift_storage.storage[1420] ),
    .S(net632),
    .X(_03791_));
 sg13g2_and2_1 _09629_ (.A(net334),
    .B(_03791_),
    .X(_00571_));
 sg13g2_mux2_1 _09630_ (.A0(\shift_storage.storage[1422] ),
    .A1(\shift_storage.storage[1421] ),
    .S(net729),
    .X(_03792_));
 sg13g2_and2_1 _09631_ (.A(net436),
    .B(_03792_),
    .X(_00572_));
 sg13g2_buf_2 fanout268 (.A(net271),
    .X(net268));
 sg13g2_mux2_1 _09633_ (.A0(\shift_storage.storage[1423] ),
    .A1(\shift_storage.storage[1422] ),
    .S(net729),
    .X(_03794_));
 sg13g2_and2_1 _09634_ (.A(net436),
    .B(_03794_),
    .X(_00573_));
 sg13g2_mux2_1 _09635_ (.A0(\shift_storage.storage[1424] ),
    .A1(\shift_storage.storage[1423] ),
    .S(net729),
    .X(_03795_));
 sg13g2_and2_1 _09636_ (.A(net436),
    .B(_03795_),
    .X(_00574_));
 sg13g2_mux2_1 _09637_ (.A0(\shift_storage.storage[1425] ),
    .A1(\shift_storage.storage[1424] ),
    .S(net729),
    .X(_03796_));
 sg13g2_and2_1 _09638_ (.A(net436),
    .B(_03796_),
    .X(_00575_));
 sg13g2_buf_1 fanout267 (.A(net289),
    .X(net267));
 sg13g2_mux2_1 _09640_ (.A0(\shift_storage.storage[1426] ),
    .A1(\shift_storage.storage[1425] ),
    .S(net634),
    .X(_03798_));
 sg13g2_and2_1 _09641_ (.A(net336),
    .B(_03798_),
    .X(_00576_));
 sg13g2_mux2_1 _09642_ (.A0(\shift_storage.storage[1427] ),
    .A1(\shift_storage.storage[1426] ),
    .S(net632),
    .X(_03799_));
 sg13g2_and2_1 _09643_ (.A(net334),
    .B(_03799_),
    .X(_00577_));
 sg13g2_mux2_1 _09644_ (.A0(\shift_storage.storage[1428] ),
    .A1(\shift_storage.storage[1427] ),
    .S(net637),
    .X(_03800_));
 sg13g2_and2_1 _09645_ (.A(net340),
    .B(_03800_),
    .X(_00578_));
 sg13g2_mux2_1 _09646_ (.A0(\shift_storage.storage[1429] ),
    .A1(\shift_storage.storage[1428] ),
    .S(net637),
    .X(_03801_));
 sg13g2_and2_1 _09647_ (.A(net341),
    .B(_03801_),
    .X(_00579_));
 sg13g2_mux2_1 _09648_ (.A0(\shift_storage.storage[142] ),
    .A1(\shift_storage.storage[141] ),
    .S(net572),
    .X(_03802_));
 sg13g2_and2_1 _09649_ (.A(net272),
    .B(_03802_),
    .X(_00580_));
 sg13g2_mux2_1 _09650_ (.A0(\shift_storage.storage[1430] ),
    .A1(\shift_storage.storage[1429] ),
    .S(net637),
    .X(_03803_));
 sg13g2_and2_1 _09651_ (.A(net340),
    .B(_03803_),
    .X(_00581_));
 sg13g2_mux2_1 _09652_ (.A0(\shift_storage.storage[1431] ),
    .A1(\shift_storage.storage[1430] ),
    .S(net637),
    .X(_03804_));
 sg13g2_and2_1 _09653_ (.A(net340),
    .B(_03804_),
    .X(_00582_));
 sg13g2_buf_1 fanout266 (.A(net267),
    .X(net266));
 sg13g2_mux2_1 _09655_ (.A0(\shift_storage.storage[1432] ),
    .A1(\shift_storage.storage[1431] ),
    .S(net637),
    .X(_03806_));
 sg13g2_and2_1 _09656_ (.A(net340),
    .B(_03806_),
    .X(_00583_));
 sg13g2_mux2_1 _09657_ (.A0(\shift_storage.storage[1433] ),
    .A1(\shift_storage.storage[1432] ),
    .S(net637),
    .X(_03807_));
 sg13g2_and2_1 _09658_ (.A(net340),
    .B(_03807_),
    .X(_00584_));
 sg13g2_mux2_1 _09659_ (.A0(\shift_storage.storage[1434] ),
    .A1(\shift_storage.storage[1433] ),
    .S(net637),
    .X(_03808_));
 sg13g2_and2_1 _09660_ (.A(net340),
    .B(_03808_),
    .X(_00585_));
 sg13g2_buf_2 fanout265 (.A(net266),
    .X(net265));
 sg13g2_mux2_1 _09662_ (.A0(\shift_storage.storage[1435] ),
    .A1(\shift_storage.storage[1434] ),
    .S(net637),
    .X(_03810_));
 sg13g2_and2_1 _09663_ (.A(net340),
    .B(_03810_),
    .X(_00586_));
 sg13g2_mux2_1 _09664_ (.A0(\shift_storage.storage[1436] ),
    .A1(\shift_storage.storage[1435] ),
    .S(net638),
    .X(_03811_));
 sg13g2_and2_1 _09665_ (.A(net341),
    .B(_03811_),
    .X(_00587_));
 sg13g2_mux2_1 _09666_ (.A0(\shift_storage.storage[1437] ),
    .A1(\shift_storage.storage[1436] ),
    .S(net638),
    .X(_03812_));
 sg13g2_and2_1 _09667_ (.A(net341),
    .B(_03812_),
    .X(_00588_));
 sg13g2_mux2_1 _09668_ (.A0(\shift_storage.storage[1438] ),
    .A1(\shift_storage.storage[1437] ),
    .S(net638),
    .X(_03813_));
 sg13g2_and2_1 _09669_ (.A(net341),
    .B(_03813_),
    .X(_00589_));
 sg13g2_mux2_1 _09670_ (.A0(\shift_storage.storage[1439] ),
    .A1(\shift_storage.storage[1438] ),
    .S(net638),
    .X(_03814_));
 sg13g2_and2_1 _09671_ (.A(net341),
    .B(_03814_),
    .X(_00590_));
 sg13g2_mux2_1 _09672_ (.A0(\shift_storage.storage[143] ),
    .A1(\shift_storage.storage[142] ),
    .S(net572),
    .X(_03815_));
 sg13g2_and2_1 _09673_ (.A(net273),
    .B(_03815_),
    .X(_00591_));
 sg13g2_mux2_1 _09674_ (.A0(\shift_storage.storage[1440] ),
    .A1(\shift_storage.storage[1439] ),
    .S(net638),
    .X(_03816_));
 sg13g2_and2_1 _09675_ (.A(net341),
    .B(_03816_),
    .X(_00592_));
 sg13g2_buf_1 fanout264 (.A(net265),
    .X(net264));
 sg13g2_buf_2 fanout263 (.A(net266),
    .X(net263));
 sg13g2_mux2_1 _09678_ (.A0(\shift_storage.storage[1441] ),
    .A1(\shift_storage.storage[1440] ),
    .S(net638),
    .X(_03819_));
 sg13g2_and2_1 _09679_ (.A(net341),
    .B(_03819_),
    .X(_00593_));
 sg13g2_mux2_1 _09680_ (.A0(\shift_storage.storage[1442] ),
    .A1(\shift_storage.storage[1441] ),
    .S(net638),
    .X(_03820_));
 sg13g2_and2_1 _09681_ (.A(net351),
    .B(_03820_),
    .X(_00594_));
 sg13g2_mux2_1 _09682_ (.A0(\shift_storage.storage[1443] ),
    .A1(\shift_storage.storage[1442] ),
    .S(net649),
    .X(_03821_));
 sg13g2_and2_1 _09683_ (.A(net351),
    .B(_03821_),
    .X(_00595_));
 sg13g2_buf_2 fanout262 (.A(net263),
    .X(net262));
 sg13g2_buf_1 fanout261 (.A(net267),
    .X(net261));
 sg13g2_mux2_1 _09686_ (.A0(\shift_storage.storage[1444] ),
    .A1(\shift_storage.storage[1443] ),
    .S(net649),
    .X(_03824_));
 sg13g2_and2_1 _09687_ (.A(net351),
    .B(_03824_),
    .X(_00596_));
 sg13g2_mux2_1 _09688_ (.A0(\shift_storage.storage[1445] ),
    .A1(\shift_storage.storage[1444] ),
    .S(net649),
    .X(_03825_));
 sg13g2_and2_1 _09689_ (.A(net349),
    .B(_03825_),
    .X(_00597_));
 sg13g2_mux2_1 _09690_ (.A0(\shift_storage.storage[1446] ),
    .A1(\shift_storage.storage[1445] ),
    .S(net647),
    .X(_03826_));
 sg13g2_and2_1 _09691_ (.A(net349),
    .B(_03826_),
    .X(_00598_));
 sg13g2_mux2_1 _09692_ (.A0(\shift_storage.storage[1447] ),
    .A1(\shift_storage.storage[1446] ),
    .S(net647),
    .X(_03827_));
 sg13g2_and2_1 _09693_ (.A(net349),
    .B(_03827_),
    .X(_00599_));
 sg13g2_mux2_1 _09694_ (.A0(\shift_storage.storage[1448] ),
    .A1(\shift_storage.storage[1447] ),
    .S(net648),
    .X(_03828_));
 sg13g2_and2_1 _09695_ (.A(net350),
    .B(_03828_),
    .X(_00600_));
 sg13g2_mux2_1 _09696_ (.A0(\shift_storage.storage[1449] ),
    .A1(\shift_storage.storage[1448] ),
    .S(net652),
    .X(_03829_));
 sg13g2_and2_1 _09697_ (.A(net350),
    .B(_03829_),
    .X(_00601_));
 sg13g2_mux2_1 _09698_ (.A0(\shift_storage.storage[144] ),
    .A1(\shift_storage.storage[143] ),
    .S(net573),
    .X(_03830_));
 sg13g2_and2_1 _09699_ (.A(net273),
    .B(_03830_),
    .X(_00602_));
 sg13g2_buf_2 fanout260 (.A(net261),
    .X(net260));
 sg13g2_mux2_1 _09701_ (.A0(\shift_storage.storage[1450] ),
    .A1(\shift_storage.storage[1449] ),
    .S(net648),
    .X(_03832_));
 sg13g2_and2_1 _09702_ (.A(net350),
    .B(_03832_),
    .X(_00603_));
 sg13g2_mux2_1 _09703_ (.A0(\shift_storage.storage[1451] ),
    .A1(\shift_storage.storage[1450] ),
    .S(net648),
    .X(_03833_));
 sg13g2_and2_1 _09704_ (.A(net350),
    .B(_03833_),
    .X(_00604_));
 sg13g2_mux2_1 _09705_ (.A0(\shift_storage.storage[1452] ),
    .A1(\shift_storage.storage[1451] ),
    .S(net648),
    .X(_03834_));
 sg13g2_and2_1 _09706_ (.A(net350),
    .B(_03834_),
    .X(_00605_));
 sg13g2_buf_2 fanout259 (.A(net261),
    .X(net259));
 sg13g2_mux2_1 _09708_ (.A0(\shift_storage.storage[1453] ),
    .A1(\shift_storage.storage[1452] ),
    .S(net652),
    .X(_03836_));
 sg13g2_and2_1 _09709_ (.A(net354),
    .B(_03836_),
    .X(_00606_));
 sg13g2_mux2_1 _09710_ (.A0(\shift_storage.storage[1454] ),
    .A1(\shift_storage.storage[1453] ),
    .S(net652),
    .X(_03837_));
 sg13g2_and2_1 _09711_ (.A(net354),
    .B(_03837_),
    .X(_00607_));
 sg13g2_mux2_1 _09712_ (.A0(\shift_storage.storage[1455] ),
    .A1(\shift_storage.storage[1454] ),
    .S(net652),
    .X(_03838_));
 sg13g2_and2_1 _09713_ (.A(net354),
    .B(_03838_),
    .X(_00608_));
 sg13g2_mux2_1 _09714_ (.A0(\shift_storage.storage[1456] ),
    .A1(\shift_storage.storage[1455] ),
    .S(net652),
    .X(_03839_));
 sg13g2_and2_1 _09715_ (.A(net354),
    .B(_03839_),
    .X(_00609_));
 sg13g2_mux2_1 _09716_ (.A0(\shift_storage.storage[1457] ),
    .A1(\shift_storage.storage[1456] ),
    .S(net652),
    .X(_03840_));
 sg13g2_and2_1 _09717_ (.A(net354),
    .B(_03840_),
    .X(_00610_));
 sg13g2_mux2_1 _09718_ (.A0(\shift_storage.storage[1458] ),
    .A1(\shift_storage.storage[1457] ),
    .S(net648),
    .X(_03841_));
 sg13g2_and2_1 _09719_ (.A(net350),
    .B(_03841_),
    .X(_00611_));
 sg13g2_mux2_1 _09720_ (.A0(\shift_storage.storage[1459] ),
    .A1(\shift_storage.storage[1458] ),
    .S(net648),
    .X(_03842_));
 sg13g2_and2_1 _09721_ (.A(net350),
    .B(_03842_),
    .X(_00612_));
 sg13g2_buf_1 fanout258 (.A(net267),
    .X(net258));
 sg13g2_mux2_1 _09723_ (.A0(\shift_storage.storage[145] ),
    .A1(\shift_storage.storage[144] ),
    .S(net573),
    .X(_03844_));
 sg13g2_and2_1 _09724_ (.A(net273),
    .B(_03844_),
    .X(_00613_));
 sg13g2_mux2_1 _09725_ (.A0(\shift_storage.storage[1460] ),
    .A1(\shift_storage.storage[1459] ),
    .S(net643),
    .X(_03845_));
 sg13g2_and2_1 _09726_ (.A(net346),
    .B(_03845_),
    .X(_00614_));
 sg13g2_mux2_1 _09727_ (.A0(\shift_storage.storage[1461] ),
    .A1(\shift_storage.storage[1460] ),
    .S(net643),
    .X(_03846_));
 sg13g2_and2_1 _09728_ (.A(net346),
    .B(_03846_),
    .X(_00615_));
 sg13g2_buf_2 fanout257 (.A(net267),
    .X(net257));
 sg13g2_mux2_1 _09730_ (.A0(\shift_storage.storage[1462] ),
    .A1(\shift_storage.storage[1461] ),
    .S(net643),
    .X(_03848_));
 sg13g2_and2_1 _09731_ (.A(net346),
    .B(_03848_),
    .X(_00616_));
 sg13g2_mux2_1 _09732_ (.A0(\shift_storage.storage[1463] ),
    .A1(\shift_storage.storage[1462] ),
    .S(net644),
    .X(_03849_));
 sg13g2_and2_1 _09733_ (.A(net346),
    .B(_03849_),
    .X(_00617_));
 sg13g2_mux2_1 _09734_ (.A0(\shift_storage.storage[1464] ),
    .A1(\shift_storage.storage[1463] ),
    .S(net643),
    .X(_03850_));
 sg13g2_and2_1 _09735_ (.A(net346),
    .B(_03850_),
    .X(_00618_));
 sg13g2_mux2_1 _09736_ (.A0(\shift_storage.storage[1465] ),
    .A1(\shift_storage.storage[1464] ),
    .S(net643),
    .X(_03851_));
 sg13g2_and2_1 _09737_ (.A(net346),
    .B(_03851_),
    .X(_00619_));
 sg13g2_mux2_1 _09738_ (.A0(\shift_storage.storage[1466] ),
    .A1(\shift_storage.storage[1465] ),
    .S(net643),
    .X(_03852_));
 sg13g2_and2_1 _09739_ (.A(net346),
    .B(_03852_),
    .X(_00620_));
 sg13g2_mux2_1 _09740_ (.A0(\shift_storage.storage[1467] ),
    .A1(\shift_storage.storage[1466] ),
    .S(net646),
    .X(_03853_));
 sg13g2_and2_1 _09741_ (.A(net348),
    .B(_03853_),
    .X(_00621_));
 sg13g2_mux2_1 _09742_ (.A0(\shift_storage.storage[1468] ),
    .A1(\shift_storage.storage[1467] ),
    .S(net645),
    .X(_03854_));
 sg13g2_and2_1 _09743_ (.A(net355),
    .B(_03854_),
    .X(_00622_));
 sg13g2_buf_1 fanout256 (.A(net289),
    .X(net256));
 sg13g2_mux2_1 _09745_ (.A0(\shift_storage.storage[1469] ),
    .A1(\shift_storage.storage[1468] ),
    .S(net646),
    .X(_03856_));
 sg13g2_and2_1 _09746_ (.A(net348),
    .B(_03856_),
    .X(_00623_));
 sg13g2_mux2_1 _09747_ (.A0(\shift_storage.storage[146] ),
    .A1(\shift_storage.storage[145] ),
    .S(net573),
    .X(_03857_));
 sg13g2_and2_1 _09748_ (.A(net273),
    .B(_03857_),
    .X(_00624_));
 sg13g2_mux2_1 _09749_ (.A0(\shift_storage.storage[1470] ),
    .A1(\shift_storage.storage[1469] ),
    .S(net645),
    .X(_03858_));
 sg13g2_and2_1 _09750_ (.A(net348),
    .B(_03858_),
    .X(_00625_));
 sg13g2_buf_1 fanout255 (.A(net256),
    .X(net255));
 sg13g2_mux2_1 _09752_ (.A0(\shift_storage.storage[1471] ),
    .A1(\shift_storage.storage[1470] ),
    .S(net645),
    .X(_03860_));
 sg13g2_and2_1 _09753_ (.A(net348),
    .B(_03860_),
    .X(_00626_));
 sg13g2_mux2_1 _09754_ (.A0(\shift_storage.storage[1472] ),
    .A1(\shift_storage.storage[1471] ),
    .S(net645),
    .X(_03861_));
 sg13g2_and2_1 _09755_ (.A(net348),
    .B(_03861_),
    .X(_00627_));
 sg13g2_mux2_1 _09756_ (.A0(\shift_storage.storage[1473] ),
    .A1(\shift_storage.storage[1472] ),
    .S(net645),
    .X(_03862_));
 sg13g2_and2_1 _09757_ (.A(net348),
    .B(_03862_),
    .X(_00628_));
 sg13g2_mux2_1 _09758_ (.A0(\shift_storage.storage[1474] ),
    .A1(\shift_storage.storage[1473] ),
    .S(net645),
    .X(_03863_));
 sg13g2_and2_1 _09759_ (.A(net348),
    .B(_03863_),
    .X(_00629_));
 sg13g2_mux2_1 _09760_ (.A0(\shift_storage.storage[1475] ),
    .A1(\shift_storage.storage[1474] ),
    .S(net645),
    .X(_03864_));
 sg13g2_and2_1 _09761_ (.A(net348),
    .B(_03864_),
    .X(_00630_));
 sg13g2_mux2_1 _09762_ (.A0(\shift_storage.storage[1476] ),
    .A1(\shift_storage.storage[1475] ),
    .S(net645),
    .X(_03865_));
 sg13g2_and2_1 _09763_ (.A(net344),
    .B(_03865_),
    .X(_00631_));
 sg13g2_mux2_1 _09764_ (.A0(\shift_storage.storage[1477] ),
    .A1(\shift_storage.storage[1476] ),
    .S(net641),
    .X(_03866_));
 sg13g2_and2_1 _09765_ (.A(net344),
    .B(_03866_),
    .X(_00632_));
 sg13g2_buf_2 fanout254 (.A(net255),
    .X(net254));
 sg13g2_mux2_1 _09767_ (.A0(\shift_storage.storage[1478] ),
    .A1(\shift_storage.storage[1477] ),
    .S(net641),
    .X(_03868_));
 sg13g2_and2_1 _09768_ (.A(net344),
    .B(_03868_),
    .X(_00633_));
 sg13g2_mux2_1 _09769_ (.A0(\shift_storage.storage[1479] ),
    .A1(\shift_storage.storage[1478] ),
    .S(net644),
    .X(_03869_));
 sg13g2_and2_1 _09770_ (.A(net343),
    .B(_03869_),
    .X(_00634_));
 sg13g2_mux2_1 _09771_ (.A0(\shift_storage.storage[147] ),
    .A1(\shift_storage.storage[146] ),
    .S(net573),
    .X(_03870_));
 sg13g2_and2_1 _09772_ (.A(net273),
    .B(_03870_),
    .X(_00635_));
 sg13g2_buf_1 fanout253 (.A(net255),
    .X(net253));
 sg13g2_mux2_1 _09774_ (.A0(\shift_storage.storage[1480] ),
    .A1(\shift_storage.storage[1479] ),
    .S(net641),
    .X(_03872_));
 sg13g2_and2_1 _09775_ (.A(net343),
    .B(_03872_),
    .X(_00636_));
 sg13g2_mux2_1 _09776_ (.A0(\shift_storage.storage[1481] ),
    .A1(\shift_storage.storage[1480] ),
    .S(net641),
    .X(_03873_));
 sg13g2_and2_1 _09777_ (.A(net344),
    .B(_03873_),
    .X(_00637_));
 sg13g2_mux2_1 _09778_ (.A0(\shift_storage.storage[1482] ),
    .A1(\shift_storage.storage[1481] ),
    .S(net641),
    .X(_03874_));
 sg13g2_and2_1 _09779_ (.A(net343),
    .B(_03874_),
    .X(_00638_));
 sg13g2_mux2_1 _09780_ (.A0(\shift_storage.storage[1483] ),
    .A1(\shift_storage.storage[1482] ),
    .S(net642),
    .X(_03875_));
 sg13g2_and2_1 _09781_ (.A(net343),
    .B(_03875_),
    .X(_00639_));
 sg13g2_mux2_1 _09782_ (.A0(\shift_storage.storage[1484] ),
    .A1(\shift_storage.storage[1483] ),
    .S(net642),
    .X(_03876_));
 sg13g2_and2_1 _09783_ (.A(net345),
    .B(_03876_),
    .X(_00640_));
 sg13g2_mux2_1 _09784_ (.A0(\shift_storage.storage[1485] ),
    .A1(\shift_storage.storage[1484] ),
    .S(net642),
    .X(_03877_));
 sg13g2_and2_1 _09785_ (.A(net345),
    .B(_03877_),
    .X(_00641_));
 sg13g2_mux2_1 _09786_ (.A0(\shift_storage.storage[1486] ),
    .A1(\shift_storage.storage[1485] ),
    .S(net642),
    .X(_03878_));
 sg13g2_and2_1 _09787_ (.A(net345),
    .B(_03878_),
    .X(_00642_));
 sg13g2_buf_1 fanout252 (.A(net255),
    .X(net252));
 sg13g2_mux2_1 _09789_ (.A0(\shift_storage.storage[1487] ),
    .A1(\shift_storage.storage[1486] ),
    .S(net643),
    .X(_03880_));
 sg13g2_and2_1 _09790_ (.A(net345),
    .B(_03880_),
    .X(_00643_));
 sg13g2_mux2_1 _09791_ (.A0(\shift_storage.storage[1488] ),
    .A1(\shift_storage.storage[1487] ),
    .S(net642),
    .X(_03881_));
 sg13g2_and2_1 _09792_ (.A(net345),
    .B(_03881_),
    .X(_00644_));
 sg13g2_mux2_1 _09793_ (.A0(\shift_storage.storage[1489] ),
    .A1(\shift_storage.storage[1488] ),
    .S(net647),
    .X(_03882_));
 sg13g2_and2_1 _09794_ (.A(net349),
    .B(_03882_),
    .X(_00645_));
 sg13g2_buf_2 fanout251 (.A(net255),
    .X(net251));
 sg13g2_mux2_1 _09796_ (.A0(\shift_storage.storage[148] ),
    .A1(\shift_storage.storage[147] ),
    .S(net573),
    .X(_03884_));
 sg13g2_and2_1 _09797_ (.A(net321),
    .B(_03884_),
    .X(_00646_));
 sg13g2_mux2_1 _09798_ (.A0(\shift_storage.storage[1490] ),
    .A1(\shift_storage.storage[1489] ),
    .S(net647),
    .X(_03885_));
 sg13g2_and2_1 _09799_ (.A(net349),
    .B(_03885_),
    .X(_00647_));
 sg13g2_mux2_1 _09800_ (.A0(\shift_storage.storage[1491] ),
    .A1(\shift_storage.storage[1490] ),
    .S(net647),
    .X(_03886_));
 sg13g2_and2_1 _09801_ (.A(net349),
    .B(_03886_),
    .X(_00648_));
 sg13g2_mux2_1 _09802_ (.A0(\shift_storage.storage[1492] ),
    .A1(\shift_storage.storage[1491] ),
    .S(net647),
    .X(_03887_));
 sg13g2_and2_1 _09803_ (.A(net349),
    .B(_03887_),
    .X(_00649_));
 sg13g2_mux2_1 _09804_ (.A0(\shift_storage.storage[1493] ),
    .A1(\shift_storage.storage[1492] ),
    .S(net647),
    .X(_03888_));
 sg13g2_and2_1 _09805_ (.A(net349),
    .B(_03888_),
    .X(_00650_));
 sg13g2_mux2_1 _09806_ (.A0(\shift_storage.storage[1494] ),
    .A1(\shift_storage.storage[1493] ),
    .S(net648),
    .X(_03889_));
 sg13g2_and2_1 _09807_ (.A(net338),
    .B(_03889_),
    .X(_00651_));
 sg13g2_mux2_1 _09808_ (.A0(\shift_storage.storage[1495] ),
    .A1(\shift_storage.storage[1494] ),
    .S(net636),
    .X(_03890_));
 sg13g2_and2_1 _09809_ (.A(net338),
    .B(_03890_),
    .X(_00652_));
 sg13g2_buf_1 fanout250 (.A(net256),
    .X(net250));
 sg13g2_mux2_1 _09811_ (.A0(\shift_storage.storage[1496] ),
    .A1(\shift_storage.storage[1495] ),
    .S(net636),
    .X(_03892_));
 sg13g2_and2_1 _09812_ (.A(net338),
    .B(_03892_),
    .X(_00653_));
 sg13g2_mux2_1 _09813_ (.A0(\shift_storage.storage[1497] ),
    .A1(\shift_storage.storage[1496] ),
    .S(net639),
    .X(_03893_));
 sg13g2_and2_1 _09814_ (.A(net339),
    .B(_03893_),
    .X(_00654_));
 sg13g2_mux2_1 _09815_ (.A0(\shift_storage.storage[1498] ),
    .A1(\shift_storage.storage[1497] ),
    .S(net636),
    .X(_03894_));
 sg13g2_and2_1 _09816_ (.A(net338),
    .B(_03894_),
    .X(_00655_));
 sg13g2_buf_2 fanout249 (.A(net250),
    .X(net249));
 sg13g2_mux2_1 _09818_ (.A0(\shift_storage.storage[1499] ),
    .A1(\shift_storage.storage[1498] ),
    .S(net635),
    .X(_03896_));
 sg13g2_and2_1 _09819_ (.A(net337),
    .B(_03896_),
    .X(_00656_));
 sg13g2_mux2_1 _09820_ (.A0(\shift_storage.storage[149] ),
    .A1(\shift_storage.storage[148] ),
    .S(net619),
    .X(_03897_));
 sg13g2_and2_1 _09821_ (.A(net321),
    .B(_03897_),
    .X(_00657_));
 sg13g2_mux2_1 _09822_ (.A0(\shift_storage.storage[14] ),
    .A1(\shift_storage.storage[13] ),
    .S(net610),
    .X(_03898_));
 sg13g2_and2_1 _09823_ (.A(net312),
    .B(_03898_),
    .X(_00658_));
 sg13g2_mux2_1 _09824_ (.A0(\shift_storage.storage[1500] ),
    .A1(\shift_storage.storage[1499] ),
    .S(net636),
    .X(_03899_));
 sg13g2_and2_1 _09825_ (.A(net339),
    .B(_03899_),
    .X(_00659_));
 sg13g2_mux2_1 _09826_ (.A0(\shift_storage.storage[1501] ),
    .A1(\shift_storage.storage[1500] ),
    .S(net635),
    .X(_03900_));
 sg13g2_and2_1 _09827_ (.A(net337),
    .B(_03900_),
    .X(_00660_));
 sg13g2_mux2_1 _09828_ (.A0(\shift_storage.storage[1502] ),
    .A1(\shift_storage.storage[1501] ),
    .S(net635),
    .X(_03901_));
 sg13g2_and2_1 _09829_ (.A(net337),
    .B(_03901_),
    .X(_00661_));
 sg13g2_mux2_1 _09830_ (.A0(\shift_storage.storage[1503] ),
    .A1(\shift_storage.storage[1502] ),
    .S(net635),
    .X(_03902_));
 sg13g2_and2_1 _09831_ (.A(net337),
    .B(_03902_),
    .X(_00662_));
 sg13g2_buf_2 fanout248 (.A(net250),
    .X(net248));
 sg13g2_buf_2 fanout247 (.A(net256),
    .X(net247));
 sg13g2_buf_2 fanout246 (.A(net247),
    .X(net246));
 sg13g2_mux2_1 _09835_ (.A0(\shift_storage.storage[1504] ),
    .A1(\shift_storage.storage[1503] ),
    .S(net635),
    .X(_03906_));
 sg13g2_and2_1 _09836_ (.A(net337),
    .B(_03906_),
    .X(_00663_));
 sg13g2_mux2_1 _09837_ (.A0(\shift_storage.storage[1505] ),
    .A1(\shift_storage.storage[1504] ),
    .S(net636),
    .X(_03907_));
 sg13g2_and2_1 _09838_ (.A(net339),
    .B(_03907_),
    .X(_00664_));
 sg13g2_mux2_1 _09839_ (.A0(\shift_storage.storage[1506] ),
    .A1(\shift_storage.storage[1505] ),
    .S(net631),
    .X(_03908_));
 sg13g2_and2_1 _09840_ (.A(net333),
    .B(_03908_),
    .X(_00665_));
 sg13g2_buf_1 fanout245 (.A(net289),
    .X(net245));
 sg13g2_buf_1 fanout244 (.A(net245),
    .X(net244));
 sg13g2_buf_1 fanout243 (.A(net244),
    .X(net243));
 sg13g2_mux2_1 _09844_ (.A0(\shift_storage.storage[1507] ),
    .A1(\shift_storage.storage[1506] ),
    .S(net632),
    .X(_03912_));
 sg13g2_and2_1 _09845_ (.A(net334),
    .B(_03912_),
    .X(_00666_));
 sg13g2_mux2_1 _09846_ (.A0(\shift_storage.storage[1508] ),
    .A1(\shift_storage.storage[1507] ),
    .S(net632),
    .X(_03913_));
 sg13g2_and2_1 _09847_ (.A(net334),
    .B(_03913_),
    .X(_00667_));
 sg13g2_mux2_1 _09848_ (.A0(\shift_storage.storage[1509] ),
    .A1(\shift_storage.storage[1508] ),
    .S(net632),
    .X(_03914_));
 sg13g2_and2_1 _09849_ (.A(net334),
    .B(_03914_),
    .X(_00668_));
 sg13g2_mux2_1 _09850_ (.A0(\shift_storage.storage[150] ),
    .A1(\shift_storage.storage[149] ),
    .S(net619),
    .X(_03915_));
 sg13g2_and2_1 _09851_ (.A(net321),
    .B(_03915_),
    .X(_00669_));
 sg13g2_mux2_1 _09852_ (.A0(\shift_storage.storage[1510] ),
    .A1(\shift_storage.storage[1509] ),
    .S(net632),
    .X(_03916_));
 sg13g2_and2_1 _09853_ (.A(net334),
    .B(_03916_),
    .X(_00670_));
 sg13g2_mux2_1 _09854_ (.A0(\shift_storage.storage[1511] ),
    .A1(\shift_storage.storage[1510] ),
    .S(net632),
    .X(_03917_));
 sg13g2_and2_1 _09855_ (.A(net334),
    .B(_03917_),
    .X(_00671_));
 sg13g2_mux2_1 _09856_ (.A0(\shift_storage.storage[1512] ),
    .A1(\shift_storage.storage[1511] ),
    .S(net632),
    .X(_03918_));
 sg13g2_and2_1 _09857_ (.A(net334),
    .B(_03918_),
    .X(_00672_));
 sg13g2_buf_1 fanout242 (.A(net243),
    .X(net242));
 sg13g2_mux2_1 _09859_ (.A0(\shift_storage.storage[1513] ),
    .A1(\shift_storage.storage[1512] ),
    .S(net630),
    .X(_03920_));
 sg13g2_and2_1 _09860_ (.A(net332),
    .B(_03920_),
    .X(_00673_));
 sg13g2_mux2_1 _09861_ (.A0(\shift_storage.storage[1514] ),
    .A1(\shift_storage.storage[1513] ),
    .S(net630),
    .X(_03921_));
 sg13g2_and2_1 _09862_ (.A(net332),
    .B(_03921_),
    .X(_00674_));
 sg13g2_mux2_1 _09863_ (.A0(\shift_storage.storage[1515] ),
    .A1(\shift_storage.storage[1514] ),
    .S(net630),
    .X(_03922_));
 sg13g2_and2_1 _09864_ (.A(net332),
    .B(_03922_),
    .X(_00675_));
 sg13g2_buf_1 fanout241 (.A(net244),
    .X(net241));
 sg13g2_mux2_1 _09866_ (.A0(\shift_storage.storage[1516] ),
    .A1(\shift_storage.storage[1515] ),
    .S(net633),
    .X(_03924_));
 sg13g2_and2_1 _09867_ (.A(net335),
    .B(_03924_),
    .X(_00676_));
 sg13g2_mux2_1 _09868_ (.A0(\shift_storage.storage[1517] ),
    .A1(\shift_storage.storage[1516] ),
    .S(net633),
    .X(_03925_));
 sg13g2_and2_1 _09869_ (.A(net335),
    .B(_03925_),
    .X(_00677_));
 sg13g2_mux2_1 _09870_ (.A0(\shift_storage.storage[1518] ),
    .A1(\shift_storage.storage[1517] ),
    .S(net633),
    .X(_03926_));
 sg13g2_and2_1 _09871_ (.A(net335),
    .B(_03926_),
    .X(_00678_));
 sg13g2_mux2_1 _09872_ (.A0(\shift_storage.storage[1519] ),
    .A1(\shift_storage.storage[1518] ),
    .S(net633),
    .X(_03927_));
 sg13g2_and2_1 _09873_ (.A(net335),
    .B(_03927_),
    .X(_00679_));
 sg13g2_mux2_1 _09874_ (.A0(\shift_storage.storage[151] ),
    .A1(\shift_storage.storage[150] ),
    .S(net619),
    .X(_03928_));
 sg13g2_and2_1 _09875_ (.A(net321),
    .B(_03928_),
    .X(_00680_));
 sg13g2_mux2_1 _09876_ (.A0(\shift_storage.storage[1520] ),
    .A1(\shift_storage.storage[1519] ),
    .S(net633),
    .X(_03929_));
 sg13g2_and2_1 _09877_ (.A(net286),
    .B(_03929_),
    .X(_00681_));
 sg13g2_mux2_1 _09878_ (.A0(\shift_storage.storage[1521] ),
    .A1(\shift_storage.storage[1520] ),
    .S(net586),
    .X(_03930_));
 sg13g2_and2_1 _09879_ (.A(net285),
    .B(_03930_),
    .X(_00682_));
 sg13g2_buf_2 fanout240 (.A(net241),
    .X(net240));
 sg13g2_mux2_1 _09881_ (.A0(\shift_storage.storage[1522] ),
    .A1(\shift_storage.storage[1521] ),
    .S(net676),
    .X(_03932_));
 sg13g2_and2_1 _09882_ (.A(net382),
    .B(_03932_),
    .X(_00683_));
 sg13g2_mux2_1 _09883_ (.A0(\shift_storage.storage[1523] ),
    .A1(\shift_storage.storage[1522] ),
    .S(net676),
    .X(_03933_));
 sg13g2_and2_1 _09884_ (.A(net382),
    .B(_03933_),
    .X(_00684_));
 sg13g2_mux2_1 _09885_ (.A0(\shift_storage.storage[1524] ),
    .A1(\shift_storage.storage[1523] ),
    .S(net680),
    .X(_03934_));
 sg13g2_and2_1 _09886_ (.A(net386),
    .B(_03934_),
    .X(_00685_));
 sg13g2_buf_1 fanout239 (.A(net241),
    .X(net239));
 sg13g2_mux2_1 _09888_ (.A0(\shift_storage.storage[1525] ),
    .A1(\shift_storage.storage[1524] ),
    .S(net680),
    .X(_03936_));
 sg13g2_and2_1 _09889_ (.A(net382),
    .B(_03936_),
    .X(_00686_));
 sg13g2_mux2_1 _09890_ (.A0(\shift_storage.storage[1526] ),
    .A1(\shift_storage.storage[1525] ),
    .S(net676),
    .X(_03937_));
 sg13g2_and2_1 _09891_ (.A(net386),
    .B(_03937_),
    .X(_00687_));
 sg13g2_mux2_1 _09892_ (.A0(\shift_storage.storage[1527] ),
    .A1(\shift_storage.storage[1526] ),
    .S(net676),
    .X(_03938_));
 sg13g2_and2_1 _09893_ (.A(net382),
    .B(_03938_),
    .X(_00688_));
 sg13g2_mux2_1 _09894_ (.A0(\shift_storage.storage[1528] ),
    .A1(\shift_storage.storage[1527] ),
    .S(net676),
    .X(_03939_));
 sg13g2_and2_1 _09895_ (.A(net382),
    .B(_03939_),
    .X(_00689_));
 sg13g2_mux2_1 _09896_ (.A0(\shift_storage.storage[1529] ),
    .A1(\shift_storage.storage[1528] ),
    .S(net676),
    .X(_03940_));
 sg13g2_and2_1 _09897_ (.A(net382),
    .B(_03940_),
    .X(_00690_));
 sg13g2_mux2_1 _09898_ (.A0(\shift_storage.storage[152] ),
    .A1(\shift_storage.storage[151] ),
    .S(net619),
    .X(_03941_));
 sg13g2_and2_1 _09899_ (.A(net321),
    .B(_03941_),
    .X(_00691_));
 sg13g2_mux2_1 _09900_ (.A0(\shift_storage.storage[1530] ),
    .A1(\shift_storage.storage[1529] ),
    .S(net676),
    .X(_03942_));
 sg13g2_and2_1 _09901_ (.A(net382),
    .B(_03942_),
    .X(_00692_));
 sg13g2_buf_1 fanout238 (.A(net244),
    .X(net238));
 sg13g2_mux2_1 _09903_ (.A0(\shift_storage.storage[1531] ),
    .A1(\shift_storage.storage[1530] ),
    .S(net676),
    .X(_03944_));
 sg13g2_and2_1 _09904_ (.A(net382),
    .B(_03944_),
    .X(_00693_));
 sg13g2_mux2_1 _09905_ (.A0(\shift_storage.storage[1532] ),
    .A1(\shift_storage.storage[1531] ),
    .S(net585),
    .X(_03945_));
 sg13g2_and2_1 _09906_ (.A(net285),
    .B(_03945_),
    .X(_00694_));
 sg13g2_mux2_1 _09907_ (.A0(\shift_storage.storage[1533] ),
    .A1(\shift_storage.storage[1532] ),
    .S(net586),
    .X(_03946_));
 sg13g2_and2_1 _09908_ (.A(net285),
    .B(_03946_),
    .X(_00695_));
 sg13g2_buf_2 fanout237 (.A(net238),
    .X(net237));
 sg13g2_mux2_1 _09910_ (.A0(\shift_storage.storage[1534] ),
    .A1(\shift_storage.storage[1533] ),
    .S(net586),
    .X(_03948_));
 sg13g2_and2_1 _09911_ (.A(net286),
    .B(_03948_),
    .X(_00696_));
 sg13g2_mux2_1 _09912_ (.A0(\shift_storage.storage[1535] ),
    .A1(\shift_storage.storage[1534] ),
    .S(net584),
    .X(_03949_));
 sg13g2_and2_1 _09913_ (.A(net284),
    .B(_03949_),
    .X(_00697_));
 sg13g2_mux2_1 _09914_ (.A0(\shift_storage.storage[1536] ),
    .A1(\shift_storage.storage[1535] ),
    .S(net584),
    .X(_03950_));
 sg13g2_and2_1 _09915_ (.A(net284),
    .B(_03950_),
    .X(_00698_));
 sg13g2_mux2_1 _09916_ (.A0(\shift_storage.storage[1537] ),
    .A1(\shift_storage.storage[1536] ),
    .S(net586),
    .X(_03951_));
 sg13g2_and2_1 _09917_ (.A(net284),
    .B(_03951_),
    .X(_00699_));
 sg13g2_mux2_1 _09918_ (.A0(\shift_storage.storage[1538] ),
    .A1(\shift_storage.storage[1537] ),
    .S(net677),
    .X(_03952_));
 sg13g2_and2_1 _09919_ (.A(net383),
    .B(_03952_),
    .X(_00700_));
 sg13g2_mux2_1 _09920_ (.A0(\shift_storage.storage[1539] ),
    .A1(\shift_storage.storage[1538] ),
    .S(net677),
    .X(_03953_));
 sg13g2_and2_1 _09921_ (.A(net383),
    .B(_03953_),
    .X(_00701_));
 sg13g2_mux2_1 _09922_ (.A0(\shift_storage.storage[153] ),
    .A1(\shift_storage.storage[152] ),
    .S(net619),
    .X(_03954_));
 sg13g2_and2_1 _09923_ (.A(net321),
    .B(_03954_),
    .X(_00702_));
 sg13g2_buf_1 fanout236 (.A(net244),
    .X(net236));
 sg13g2_mux2_1 _09925_ (.A0(\shift_storage.storage[1540] ),
    .A1(\shift_storage.storage[1539] ),
    .S(net677),
    .X(_03956_));
 sg13g2_and2_1 _09926_ (.A(net383),
    .B(_03956_),
    .X(_00703_));
 sg13g2_mux2_1 _09927_ (.A0(\shift_storage.storage[1541] ),
    .A1(\shift_storage.storage[1540] ),
    .S(net677),
    .X(_03957_));
 sg13g2_and2_1 _09928_ (.A(net383),
    .B(_03957_),
    .X(_00704_));
 sg13g2_mux2_1 _09929_ (.A0(\shift_storage.storage[1542] ),
    .A1(\shift_storage.storage[1541] ),
    .S(net677),
    .X(_03958_));
 sg13g2_and2_1 _09930_ (.A(net383),
    .B(_03958_),
    .X(_00705_));
 sg13g2_buf_1 fanout235 (.A(net236),
    .X(net235));
 sg13g2_mux2_1 _09932_ (.A0(\shift_storage.storage[1543] ),
    .A1(\shift_storage.storage[1542] ),
    .S(net677),
    .X(_03960_));
 sg13g2_and2_1 _09933_ (.A(net383),
    .B(_03960_),
    .X(_00706_));
 sg13g2_mux2_1 _09934_ (.A0(\shift_storage.storage[1544] ),
    .A1(\shift_storage.storage[1543] ),
    .S(net678),
    .X(_03961_));
 sg13g2_and2_1 _09935_ (.A(net384),
    .B(_03961_),
    .X(_00707_));
 sg13g2_mux2_1 _09936_ (.A0(\shift_storage.storage[1545] ),
    .A1(\shift_storage.storage[1544] ),
    .S(net678),
    .X(_03962_));
 sg13g2_and2_1 _09937_ (.A(net384),
    .B(_03962_),
    .X(_00708_));
 sg13g2_mux2_1 _09938_ (.A0(\shift_storage.storage[1546] ),
    .A1(\shift_storage.storage[1545] ),
    .S(net678),
    .X(_03963_));
 sg13g2_and2_1 _09939_ (.A(net384),
    .B(_03963_),
    .X(_00709_));
 sg13g2_mux2_1 _09940_ (.A0(\shift_storage.storage[1547] ),
    .A1(\shift_storage.storage[1546] ),
    .S(net678),
    .X(_03964_));
 sg13g2_and2_1 _09941_ (.A(net384),
    .B(_03964_),
    .X(_00710_));
 sg13g2_mux2_1 _09942_ (.A0(\shift_storage.storage[1548] ),
    .A1(\shift_storage.storage[1547] ),
    .S(net687),
    .X(_03965_));
 sg13g2_and2_1 _09943_ (.A(net393),
    .B(_03965_),
    .X(_00711_));
 sg13g2_mux2_1 _09944_ (.A0(\shift_storage.storage[1549] ),
    .A1(\shift_storage.storage[1548] ),
    .S(net687),
    .X(_03966_));
 sg13g2_and2_1 _09945_ (.A(net393),
    .B(_03966_),
    .X(_00712_));
 sg13g2_buf_1 fanout234 (.A(net245),
    .X(net234));
 sg13g2_mux2_1 _09947_ (.A0(\shift_storage.storage[154] ),
    .A1(\shift_storage.storage[153] ),
    .S(net620),
    .X(_03968_));
 sg13g2_and2_1 _09948_ (.A(net326),
    .B(_03968_),
    .X(_00713_));
 sg13g2_mux2_1 _09949_ (.A0(\shift_storage.storage[1550] ),
    .A1(\shift_storage.storage[1549] ),
    .S(net687),
    .X(_03969_));
 sg13g2_and2_1 _09950_ (.A(net393),
    .B(_03969_),
    .X(_00714_));
 sg13g2_mux2_1 _09951_ (.A0(\shift_storage.storage[1551] ),
    .A1(\shift_storage.storage[1550] ),
    .S(net687),
    .X(_03970_));
 sg13g2_and2_1 _09952_ (.A(net393),
    .B(_03970_),
    .X(_00715_));
 sg13g2_buf_2 fanout233 (.A(net234),
    .X(net233));
 sg13g2_mux2_1 _09954_ (.A0(\shift_storage.storage[1552] ),
    .A1(\shift_storage.storage[1551] ),
    .S(net687),
    .X(_03972_));
 sg13g2_and2_1 _09955_ (.A(net393),
    .B(_03972_),
    .X(_00716_));
 sg13g2_mux2_1 _09956_ (.A0(\shift_storage.storage[1553] ),
    .A1(\shift_storage.storage[1552] ),
    .S(net692),
    .X(_03973_));
 sg13g2_and2_1 _09957_ (.A(net393),
    .B(_03973_),
    .X(_00717_));
 sg13g2_mux2_1 _09958_ (.A0(\shift_storage.storage[1554] ),
    .A1(\shift_storage.storage[1553] ),
    .S(net690),
    .X(_03974_));
 sg13g2_and2_1 _09959_ (.A(net394),
    .B(_03974_),
    .X(_00718_));
 sg13g2_mux2_1 _09960_ (.A0(\shift_storage.storage[1555] ),
    .A1(\shift_storage.storage[1554] ),
    .S(net690),
    .X(_03975_));
 sg13g2_and2_1 _09961_ (.A(net394),
    .B(_03975_),
    .X(_00719_));
 sg13g2_mux2_1 _09962_ (.A0(\shift_storage.storage[1556] ),
    .A1(\shift_storage.storage[1555] ),
    .S(net742),
    .X(_03976_));
 sg13g2_and2_1 _09963_ (.A(net446),
    .B(_03976_),
    .X(_00720_));
 sg13g2_mux2_1 _09964_ (.A0(\shift_storage.storage[1557] ),
    .A1(\shift_storage.storage[1556] ),
    .S(net742),
    .X(_03977_));
 sg13g2_and2_1 _09965_ (.A(net449),
    .B(_03977_),
    .X(_00721_));
 sg13g2_mux2_1 _09966_ (.A0(\shift_storage.storage[1558] ),
    .A1(\shift_storage.storage[1557] ),
    .S(net742),
    .X(_03978_));
 sg13g2_and2_1 _09967_ (.A(net449),
    .B(_03978_),
    .X(_00722_));
 sg13g2_buf_2 fanout232 (.A(net233),
    .X(net232));
 sg13g2_mux2_1 _09969_ (.A0(\shift_storage.storage[1559] ),
    .A1(\shift_storage.storage[1558] ),
    .S(net742),
    .X(_03980_));
 sg13g2_and2_1 _09970_ (.A(net449),
    .B(_03980_),
    .X(_00723_));
 sg13g2_mux2_1 _09971_ (.A0(\shift_storage.storage[155] ),
    .A1(\shift_storage.storage[154] ),
    .S(net620),
    .X(_03981_));
 sg13g2_and2_1 _09972_ (.A(net302),
    .B(_03981_),
    .X(_00724_));
 sg13g2_mux2_1 _09973_ (.A0(\shift_storage.storage[1560] ),
    .A1(\shift_storage.storage[1559] ),
    .S(net742),
    .X(_03982_));
 sg13g2_and2_1 _09974_ (.A(net449),
    .B(_03982_),
    .X(_00725_));
 sg13g2_buf_1 fanout231 (.A(net234),
    .X(net231));
 sg13g2_mux2_1 _09976_ (.A0(\shift_storage.storage[1561] ),
    .A1(\shift_storage.storage[1560] ),
    .S(net743),
    .X(_03984_));
 sg13g2_and2_1 _09977_ (.A(net450),
    .B(_03984_),
    .X(_00726_));
 sg13g2_mux2_1 _09978_ (.A0(\shift_storage.storage[1562] ),
    .A1(\shift_storage.storage[1561] ),
    .S(net743),
    .X(_03985_));
 sg13g2_and2_1 _09979_ (.A(net450),
    .B(_03985_),
    .X(_00727_));
 sg13g2_mux2_1 _09980_ (.A0(\shift_storage.storage[1563] ),
    .A1(\shift_storage.storage[1562] ),
    .S(net743),
    .X(_03986_));
 sg13g2_and2_1 _09981_ (.A(net450),
    .B(_03986_),
    .X(_00728_));
 sg13g2_mux2_1 _09982_ (.A0(\shift_storage.storage[1564] ),
    .A1(\shift_storage.storage[1563] ),
    .S(net743),
    .X(_03987_));
 sg13g2_and2_1 _09983_ (.A(net450),
    .B(_03987_),
    .X(_00729_));
 sg13g2_mux2_1 _09984_ (.A0(\shift_storage.storage[1565] ),
    .A1(\shift_storage.storage[1564] ),
    .S(net762),
    .X(_03988_));
 sg13g2_and2_1 _09985_ (.A(net475),
    .B(_03988_),
    .X(_00730_));
 sg13g2_mux2_1 _09986_ (.A0(\shift_storage.storage[1566] ),
    .A1(\shift_storage.storage[1565] ),
    .S(net759),
    .X(_03989_));
 sg13g2_and2_1 _09987_ (.A(net472),
    .B(_03989_),
    .X(_00731_));
 sg13g2_mux2_1 _09988_ (.A0(\shift_storage.storage[1567] ),
    .A1(\shift_storage.storage[1566] ),
    .S(net763),
    .X(_03990_));
 sg13g2_and2_1 _09989_ (.A(net452),
    .B(_03990_),
    .X(_00732_));
 sg13g2_buf_1 fanout230 (.A(net234),
    .X(net230));
 sg13g2_buf_1 fanout229 (.A(net245),
    .X(net229));
 sg13g2_mux2_1 _09992_ (.A0(\shift_storage.storage[1568] ),
    .A1(\shift_storage.storage[1567] ),
    .S(net763),
    .X(_03993_));
 sg13g2_and2_1 _09993_ (.A(net476),
    .B(_03993_),
    .X(_00733_));
 sg13g2_mux2_1 _09994_ (.A0(\shift_storage.storage[1569] ),
    .A1(\shift_storage.storage[1568] ),
    .S(net763),
    .X(_03994_));
 sg13g2_and2_1 _09995_ (.A(net476),
    .B(_03994_),
    .X(_00734_));
 sg13g2_mux2_1 _09996_ (.A0(\shift_storage.storage[156] ),
    .A1(\shift_storage.storage[155] ),
    .S(net620),
    .X(_03995_));
 sg13g2_and2_1 _09997_ (.A(net304),
    .B(_03995_),
    .X(_00735_));
 sg13g2_buf_2 fanout228 (.A(net229),
    .X(net228));
 sg13g2_buf_1 fanout227 (.A(net228),
    .X(net227));
 sg13g2_mux2_1 _10000_ (.A0(\shift_storage.storage[1570] ),
    .A1(\shift_storage.storage[1569] ),
    .S(net763),
    .X(_03998_));
 sg13g2_and2_1 _10001_ (.A(net476),
    .B(_03998_),
    .X(_00736_));
 sg13g2_mux2_1 _10002_ (.A0(\shift_storage.storage[1571] ),
    .A1(\shift_storage.storage[1570] ),
    .S(net763),
    .X(_03999_));
 sg13g2_and2_1 _10003_ (.A(net476),
    .B(_03999_),
    .X(_00737_));
 sg13g2_mux2_1 _10004_ (.A0(\shift_storage.storage[1572] ),
    .A1(\shift_storage.storage[1571] ),
    .S(net764),
    .X(_04000_));
 sg13g2_and2_1 _10005_ (.A(net478),
    .B(_04000_),
    .X(_00738_));
 sg13g2_mux2_1 _10006_ (.A0(\shift_storage.storage[1573] ),
    .A1(\shift_storage.storage[1572] ),
    .S(net764),
    .X(_04001_));
 sg13g2_and2_1 _10007_ (.A(net478),
    .B(_04001_),
    .X(_00739_));
 sg13g2_mux2_1 _10008_ (.A0(\shift_storage.storage[1574] ),
    .A1(\shift_storage.storage[1573] ),
    .S(net763),
    .X(_04002_));
 sg13g2_and2_1 _10009_ (.A(net478),
    .B(_04002_),
    .X(_00740_));
 sg13g2_mux2_1 _10010_ (.A0(\shift_storage.storage[1575] ),
    .A1(\shift_storage.storage[1574] ),
    .S(net763),
    .X(_04003_));
 sg13g2_and2_1 _10011_ (.A(net478),
    .B(_04003_),
    .X(_00741_));
 sg13g2_mux2_1 _10012_ (.A0(\shift_storage.storage[1576] ),
    .A1(\shift_storage.storage[1575] ),
    .S(net763),
    .X(_04004_));
 sg13g2_and2_1 _10013_ (.A(net478),
    .B(_04004_),
    .X(_00742_));
 sg13g2_buf_1 fanout226 (.A(net229),
    .X(net226));
 sg13g2_mux2_1 _10015_ (.A0(\shift_storage.storage[1577] ),
    .A1(\shift_storage.storage[1576] ),
    .S(net766),
    .X(_04006_));
 sg13g2_and2_1 _10016_ (.A(net482),
    .B(_04006_),
    .X(_00743_));
 sg13g2_mux2_1 _10017_ (.A0(\shift_storage.storage[1578] ),
    .A1(\shift_storage.storage[1577] ),
    .S(net766),
    .X(_04007_));
 sg13g2_and2_1 _10018_ (.A(net482),
    .B(_04007_),
    .X(_00744_));
 sg13g2_mux2_1 _10019_ (.A0(\shift_storage.storage[1579] ),
    .A1(\shift_storage.storage[1578] ),
    .S(net766),
    .X(_04008_));
 sg13g2_and2_1 _10020_ (.A(net482),
    .B(_04008_),
    .X(_00745_));
 sg13g2_buf_1 fanout225 (.A(net245),
    .X(net225));
 sg13g2_mux2_1 _10022_ (.A0(\shift_storage.storage[157] ),
    .A1(\shift_storage.storage[156] ),
    .S(net620),
    .X(_04010_));
 sg13g2_and2_1 _10023_ (.A(net326),
    .B(_04010_),
    .X(_00746_));
 sg13g2_mux2_1 _10024_ (.A0(\shift_storage.storage[1580] ),
    .A1(\shift_storage.storage[1579] ),
    .S(net766),
    .X(_04011_));
 sg13g2_and2_1 _10025_ (.A(net482),
    .B(_04011_),
    .X(_00747_));
 sg13g2_mux2_1 _10026_ (.A0(\shift_storage.storage[1581] ),
    .A1(\shift_storage.storage[1580] ),
    .S(net766),
    .X(_04012_));
 sg13g2_and2_1 _10027_ (.A(net482),
    .B(_04012_),
    .X(_00748_));
 sg13g2_mux2_1 _10028_ (.A0(\shift_storage.storage[1582] ),
    .A1(\shift_storage.storage[1581] ),
    .S(net766),
    .X(_04013_));
 sg13g2_and2_1 _10029_ (.A(net482),
    .B(_04013_),
    .X(_00749_));
 sg13g2_mux2_1 _10030_ (.A0(\shift_storage.storage[1583] ),
    .A1(\shift_storage.storage[1582] ),
    .S(net766),
    .X(_04014_));
 sg13g2_and2_1 _10031_ (.A(net482),
    .B(_04014_),
    .X(_00750_));
 sg13g2_mux2_1 _10032_ (.A0(\shift_storage.storage[1584] ),
    .A1(\shift_storage.storage[1583] ),
    .S(net766),
    .X(_04015_));
 sg13g2_and2_1 _10033_ (.A(net482),
    .B(_04015_),
    .X(_00751_));
 sg13g2_mux2_1 _10034_ (.A0(\shift_storage.storage[1585] ),
    .A1(\shift_storage.storage[1584] ),
    .S(net767),
    .X(_04016_));
 sg13g2_and2_1 _10035_ (.A(net483),
    .B(_04016_),
    .X(_00752_));
 sg13g2_buf_2 fanout224 (.A(net225),
    .X(net224));
 sg13g2_mux2_1 _10037_ (.A0(\shift_storage.storage[1586] ),
    .A1(\shift_storage.storage[1585] ),
    .S(net767),
    .X(_04018_));
 sg13g2_and2_1 _10038_ (.A(net483),
    .B(_04018_),
    .X(_00753_));
 sg13g2_mux2_1 _10039_ (.A0(\shift_storage.storage[1587] ),
    .A1(\shift_storage.storage[1586] ),
    .S(net772),
    .X(_04019_));
 sg13g2_and2_1 _10040_ (.A(net491),
    .B(_04019_),
    .X(_00754_));
 sg13g2_mux2_1 _10041_ (.A0(\shift_storage.storage[1588] ),
    .A1(\shift_storage.storage[1587] ),
    .S(net772),
    .X(_04020_));
 sg13g2_and2_1 _10042_ (.A(net487),
    .B(_04020_),
    .X(_00755_));
 sg13g2_buf_1 fanout223 (.A(net224),
    .X(net223));
 sg13g2_mux2_1 _10044_ (.A0(\shift_storage.storage[1589] ),
    .A1(\shift_storage.storage[1588] ),
    .S(net772),
    .X(_04022_));
 sg13g2_and2_1 _10045_ (.A(net487),
    .B(_04022_),
    .X(_00756_));
 sg13g2_mux2_1 _10046_ (.A0(\shift_storage.storage[158] ),
    .A1(\shift_storage.storage[157] ),
    .S(net625),
    .X(_04023_));
 sg13g2_and2_1 _10047_ (.A(net327),
    .B(_04023_),
    .X(_00757_));
 sg13g2_mux2_1 _10048_ (.A0(\shift_storage.storage[1590] ),
    .A1(\shift_storage.storage[1589] ),
    .S(net772),
    .X(_04024_));
 sg13g2_and2_1 _10049_ (.A(net491),
    .B(_04024_),
    .X(_00758_));
 sg13g2_mux2_1 _10050_ (.A0(\shift_storage.storage[1591] ),
    .A1(\shift_storage.storage[1590] ),
    .S(net772),
    .X(_04025_));
 sg13g2_and2_1 _10051_ (.A(net487),
    .B(_04025_),
    .X(_00759_));
 sg13g2_mux2_1 _10052_ (.A0(\shift_storage.storage[1592] ),
    .A1(\shift_storage.storage[1591] ),
    .S(net772),
    .X(_04026_));
 sg13g2_and2_1 _10053_ (.A(net487),
    .B(_04026_),
    .X(_00760_));
 sg13g2_mux2_1 _10054_ (.A0(\shift_storage.storage[1593] ),
    .A1(\shift_storage.storage[1592] ),
    .S(net772),
    .X(_04027_));
 sg13g2_and2_1 _10055_ (.A(net487),
    .B(_04027_),
    .X(_00761_));
 sg13g2_mux2_1 _10056_ (.A0(\shift_storage.storage[1594] ),
    .A1(\shift_storage.storage[1593] ),
    .S(net772),
    .X(_04028_));
 sg13g2_and2_1 _10057_ (.A(net487),
    .B(_04028_),
    .X(_00762_));
 sg13g2_buf_1 fanout222 (.A(net225),
    .X(net222));
 sg13g2_mux2_1 _10059_ (.A0(\shift_storage.storage[1595] ),
    .A1(\shift_storage.storage[1594] ),
    .S(net770),
    .X(_04030_));
 sg13g2_and2_1 _10060_ (.A(net489),
    .B(_04030_),
    .X(_00763_));
 sg13g2_mux2_1 _10061_ (.A0(\shift_storage.storage[1596] ),
    .A1(\shift_storage.storage[1595] ),
    .S(net770),
    .X(_04031_));
 sg13g2_and2_1 _10062_ (.A(net489),
    .B(_04031_),
    .X(_00764_));
 sg13g2_mux2_1 _10063_ (.A0(\shift_storage.storage[1597] ),
    .A1(\shift_storage.storage[1596] ),
    .S(net770),
    .X(_04032_));
 sg13g2_and2_1 _10064_ (.A(net489),
    .B(_04032_),
    .X(_00765_));
 sg13g2_buf_2 fanout221 (.A(net225),
    .X(net221));
 sg13g2_mux2_1 _10066_ (.A0(\shift_storage.storage[1598] ),
    .A1(\shift_storage.storage[1597] ),
    .S(net770),
    .X(_04034_));
 sg13g2_and2_1 _10067_ (.A(net489),
    .B(_04034_),
    .X(_00766_));
 sg13g2_mux2_1 _10068_ (.A0(\shift_storage.shreg_out ),
    .A1(\shift_storage.storage[1598] ),
    .S(net769),
    .X(_04035_));
 sg13g2_and2_1 _10069_ (.A(net488),
    .B(_04035_),
    .X(_00767_));
 sg13g2_mux2_1 _10070_ (.A0(\shift_storage.storage[159] ),
    .A1(\shift_storage.storage[158] ),
    .S(net625),
    .X(_04036_));
 sg13g2_and2_1 _10071_ (.A(net327),
    .B(_04036_),
    .X(_00768_));
 sg13g2_mux2_1 _10072_ (.A0(\shift_storage.storage[15] ),
    .A1(\shift_storage.storage[14] ),
    .S(net614),
    .X(_04037_));
 sg13g2_and2_1 _10073_ (.A(net316),
    .B(_04037_),
    .X(_00769_));
 sg13g2_mux2_1 _10074_ (.A0(\shift_storage.storage[160] ),
    .A1(\shift_storage.storage[159] ),
    .S(net625),
    .X(_04038_));
 sg13g2_and2_1 _10075_ (.A(net327),
    .B(_04038_),
    .X(_00770_));
 sg13g2_mux2_1 _10076_ (.A0(\shift_storage.storage[161] ),
    .A1(\shift_storage.storage[160] ),
    .S(net607),
    .X(_04039_));
 sg13g2_and2_1 _10077_ (.A(net309),
    .B(_04039_),
    .X(_00771_));
 sg13g2_mux2_1 _10078_ (.A0(\shift_storage.storage[162] ),
    .A1(\shift_storage.storage[161] ),
    .S(net607),
    .X(_04040_));
 sg13g2_and2_1 _10079_ (.A(net308),
    .B(_04040_),
    .X(_00772_));
 sg13g2_buf_2 fanout220 (.A(net225),
    .X(net220));
 sg13g2_mux2_1 _10081_ (.A0(\shift_storage.storage[163] ),
    .A1(\shift_storage.storage[162] ),
    .S(net601),
    .X(_04042_));
 sg13g2_and2_1 _10082_ (.A(net302),
    .B(_04042_),
    .X(_00773_));
 sg13g2_mux2_1 _10083_ (.A0(\shift_storage.storage[164] ),
    .A1(\shift_storage.storage[163] ),
    .S(net601),
    .X(_04043_));
 sg13g2_and2_1 _10084_ (.A(net304),
    .B(_04043_),
    .X(_00774_));
 sg13g2_mux2_1 _10085_ (.A0(\shift_storage.storage[165] ),
    .A1(\shift_storage.storage[164] ),
    .S(net601),
    .X(_04044_));
 sg13g2_and2_1 _10086_ (.A(net302),
    .B(_04044_),
    .X(_00775_));
 sg13g2_buf_1 fanout219 (.A(net220),
    .X(net219));
 sg13g2_mux2_1 _10088_ (.A0(\shift_storage.storage[166] ),
    .A1(\shift_storage.storage[165] ),
    .S(net601),
    .X(_04046_));
 sg13g2_and2_1 _10089_ (.A(net302),
    .B(_04046_),
    .X(_00776_));
 sg13g2_mux2_1 _10090_ (.A0(\shift_storage.storage[167] ),
    .A1(\shift_storage.storage[166] ),
    .S(net601),
    .X(_04047_));
 sg13g2_and2_1 _10091_ (.A(net302),
    .B(_04047_),
    .X(_00777_));
 sg13g2_mux2_1 _10092_ (.A0(\shift_storage.storage[168] ),
    .A1(\shift_storage.storage[167] ),
    .S(net601),
    .X(_04048_));
 sg13g2_and2_1 _10093_ (.A(net302),
    .B(_04048_),
    .X(_00778_));
 sg13g2_mux2_1 _10094_ (.A0(\shift_storage.storage[169] ),
    .A1(\shift_storage.storage[168] ),
    .S(net601),
    .X(_04049_));
 sg13g2_and2_1 _10095_ (.A(net302),
    .B(_04049_),
    .X(_00779_));
 sg13g2_mux2_1 _10096_ (.A0(\shift_storage.storage[16] ),
    .A1(\shift_storage.storage[15] ),
    .S(net614),
    .X(_04050_));
 sg13g2_and2_1 _10097_ (.A(net316),
    .B(_04050_),
    .X(_00780_));
 sg13g2_mux2_1 _10098_ (.A0(\shift_storage.storage[170] ),
    .A1(\shift_storage.storage[169] ),
    .S(net601),
    .X(_04051_));
 sg13g2_and2_1 _10099_ (.A(net302),
    .B(_04051_),
    .X(_00781_));
 sg13g2_mux2_1 _10100_ (.A0(\shift_storage.storage[171] ),
    .A1(\shift_storage.storage[170] ),
    .S(net603),
    .X(_04052_));
 sg13g2_and2_1 _10101_ (.A(net304),
    .B(_04052_),
    .X(_00782_));
 sg13g2_buf_1 fanout218 (.A(net225),
    .X(net218));
 sg13g2_mux2_1 _10103_ (.A0(\shift_storage.storage[172] ),
    .A1(\shift_storage.storage[171] ),
    .S(net602),
    .X(_04054_));
 sg13g2_and2_1 _10104_ (.A(net303),
    .B(_04054_),
    .X(_00783_));
 sg13g2_mux2_1 _10105_ (.A0(\shift_storage.storage[173] ),
    .A1(\shift_storage.storage[172] ),
    .S(net602),
    .X(_04055_));
 sg13g2_and2_1 _10106_ (.A(net303),
    .B(_04055_),
    .X(_00784_));
 sg13g2_mux2_1 _10107_ (.A0(\shift_storage.storage[174] ),
    .A1(\shift_storage.storage[173] ),
    .S(net602),
    .X(_04056_));
 sg13g2_and2_1 _10108_ (.A(net303),
    .B(_04056_),
    .X(_00785_));
 sg13g2_buf_1 fanout217 (.A(net218),
    .X(net217));
 sg13g2_mux2_1 _10110_ (.A0(\shift_storage.storage[175] ),
    .A1(\shift_storage.storage[174] ),
    .S(net602),
    .X(_04058_));
 sg13g2_and2_1 _10111_ (.A(net303),
    .B(_04058_),
    .X(_00786_));
 sg13g2_mux2_1 _10112_ (.A0(\shift_storage.storage[176] ),
    .A1(\shift_storage.storage[175] ),
    .S(net602),
    .X(_04059_));
 sg13g2_and2_1 _10113_ (.A(net303),
    .B(_04059_),
    .X(_00787_));
 sg13g2_mux2_1 _10114_ (.A0(\shift_storage.storage[177] ),
    .A1(\shift_storage.storage[176] ),
    .S(net602),
    .X(_04060_));
 sg13g2_and2_1 _10115_ (.A(net303),
    .B(_04060_),
    .X(_00788_));
 sg13g2_mux2_1 _10116_ (.A0(\shift_storage.storage[178] ),
    .A1(\shift_storage.storage[177] ),
    .S(net602),
    .X(_04061_));
 sg13g2_and2_1 _10117_ (.A(net303),
    .B(_04061_),
    .X(_00789_));
 sg13g2_mux2_1 _10118_ (.A0(\shift_storage.storage[179] ),
    .A1(\shift_storage.storage[178] ),
    .S(net544),
    .X(_04062_));
 sg13g2_and2_1 _10119_ (.A(net243),
    .B(_04062_),
    .X(_00790_));
 sg13g2_mux2_1 _10120_ (.A0(\shift_storage.storage[17] ),
    .A1(\shift_storage.storage[16] ),
    .S(net615),
    .X(_04063_));
 sg13g2_and2_1 _10121_ (.A(net316),
    .B(_04063_),
    .X(_00791_));
 sg13g2_mux2_1 _10122_ (.A0(\shift_storage.storage[180] ),
    .A1(\shift_storage.storage[179] ),
    .S(net542),
    .X(_04064_));
 sg13g2_and2_1 _10123_ (.A(net242),
    .B(_04064_),
    .X(_00792_));
 sg13g2_buf_1 fanout216 (.A(net218),
    .X(net216));
 sg13g2_mux2_1 _10125_ (.A0(\shift_storage.storage[181] ),
    .A1(\shift_storage.storage[180] ),
    .S(net542),
    .X(_04066_));
 sg13g2_and2_1 _10126_ (.A(net242),
    .B(_04066_),
    .X(_00793_));
 sg13g2_mux2_1 _10127_ (.A0(\shift_storage.storage[182] ),
    .A1(\shift_storage.storage[181] ),
    .S(net544),
    .X(_04067_));
 sg13g2_and2_1 _10128_ (.A(net242),
    .B(_04067_),
    .X(_00794_));
 sg13g2_mux2_1 _10129_ (.A0(\shift_storage.storage[183] ),
    .A1(\shift_storage.storage[182] ),
    .S(net542),
    .X(_04068_));
 sg13g2_and2_1 _10130_ (.A(net242),
    .B(_04068_),
    .X(_00795_));
 sg13g2_buf_1 fanout215 (.A(net245),
    .X(net215));
 sg13g2_mux2_1 _10132_ (.A0(\shift_storage.storage[184] ),
    .A1(\shift_storage.storage[183] ),
    .S(net542),
    .X(_04070_));
 sg13g2_and2_1 _10133_ (.A(net242),
    .B(_04070_),
    .X(_00796_));
 sg13g2_mux2_1 _10134_ (.A0(\shift_storage.storage[185] ),
    .A1(\shift_storage.storage[184] ),
    .S(net542),
    .X(_04071_));
 sg13g2_and2_1 _10135_ (.A(net240),
    .B(_04071_),
    .X(_00797_));
 sg13g2_mux2_1 _10136_ (.A0(\shift_storage.storage[186] ),
    .A1(\shift_storage.storage[185] ),
    .S(net541),
    .X(_04072_));
 sg13g2_and2_1 _10137_ (.A(net241),
    .B(_04072_),
    .X(_00798_));
 sg13g2_mux2_1 _10138_ (.A0(\shift_storage.storage[187] ),
    .A1(\shift_storage.storage[186] ),
    .S(net541),
    .X(_04073_));
 sg13g2_and2_1 _10139_ (.A(net240),
    .B(_04073_),
    .X(_00799_));
 sg13g2_mux2_1 _10140_ (.A0(\shift_storage.storage[188] ),
    .A1(\shift_storage.storage[187] ),
    .S(net541),
    .X(_04074_));
 sg13g2_and2_1 _10141_ (.A(net240),
    .B(_04074_),
    .X(_00800_));
 sg13g2_mux2_1 _10142_ (.A0(\shift_storage.storage[189] ),
    .A1(\shift_storage.storage[188] ),
    .S(net541),
    .X(_04075_));
 sg13g2_and2_1 _10143_ (.A(net240),
    .B(_04075_),
    .X(_00801_));
 sg13g2_mux2_1 _10144_ (.A0(\shift_storage.storage[18] ),
    .A1(\shift_storage.storage[17] ),
    .S(net614),
    .X(_04076_));
 sg13g2_and2_1 _10145_ (.A(net317),
    .B(_04076_),
    .X(_00802_));
 sg13g2_buf_1 fanout214 (.A(net215),
    .X(net214));
 sg13g2_buf_2 fanout213 (.A(net215),
    .X(net213));
 sg13g2_mux2_1 _10148_ (.A0(\shift_storage.storage[190] ),
    .A1(\shift_storage.storage[189] ),
    .S(net598),
    .X(_04079_));
 sg13g2_and2_1 _10149_ (.A(net300),
    .B(_04079_),
    .X(_00803_));
 sg13g2_mux2_1 _10150_ (.A0(\shift_storage.storage[191] ),
    .A1(\shift_storage.storage[190] ),
    .S(net600),
    .X(_04080_));
 sg13g2_and2_1 _10151_ (.A(net300),
    .B(_04080_),
    .X(_00804_));
 sg13g2_mux2_1 _10152_ (.A0(\shift_storage.storage[192] ),
    .A1(\shift_storage.storage[191] ),
    .S(net598),
    .X(_04081_));
 sg13g2_and2_1 _10153_ (.A(net300),
    .B(_04081_),
    .X(_00805_));
 sg13g2_buf_1 fanout212 (.A(net215),
    .X(net212));
 sg13g2_buf_1 fanout211 (.A(net215),
    .X(net211));
 sg13g2_mux2_1 _10156_ (.A0(\shift_storage.storage[193] ),
    .A1(\shift_storage.storage[192] ),
    .S(net598),
    .X(_04084_));
 sg13g2_and2_1 _10157_ (.A(net300),
    .B(_04084_),
    .X(_00806_));
 sg13g2_mux2_1 _10158_ (.A0(\shift_storage.storage[194] ),
    .A1(\shift_storage.storage[193] ),
    .S(net602),
    .X(_04085_));
 sg13g2_and2_1 _10159_ (.A(net303),
    .B(_04085_),
    .X(_00807_));
 sg13g2_mux2_1 _10160_ (.A0(\shift_storage.storage[195] ),
    .A1(\shift_storage.storage[194] ),
    .S(net598),
    .X(_04086_));
 sg13g2_and2_1 _10161_ (.A(net301),
    .B(_04086_),
    .X(_00808_));
 sg13g2_mux2_1 _10162_ (.A0(\shift_storage.storage[196] ),
    .A1(\shift_storage.storage[195] ),
    .S(net598),
    .X(_04087_));
 sg13g2_and2_1 _10163_ (.A(net300),
    .B(_04087_),
    .X(_00809_));
 sg13g2_mux2_1 _10164_ (.A0(\shift_storage.storage[197] ),
    .A1(\shift_storage.storage[196] ),
    .S(net600),
    .X(_04088_));
 sg13g2_and2_1 _10165_ (.A(net301),
    .B(_04088_),
    .X(_00810_));
 sg13g2_mux2_1 _10166_ (.A0(\shift_storage.storage[198] ),
    .A1(\shift_storage.storage[197] ),
    .S(net600),
    .X(_04089_));
 sg13g2_and2_1 _10167_ (.A(net301),
    .B(_04089_),
    .X(_00811_));
 sg13g2_mux2_1 _10168_ (.A0(\shift_storage.storage[199] ),
    .A1(\shift_storage.storage[198] ),
    .S(net599),
    .X(_04090_));
 sg13g2_and2_1 _10169_ (.A(net301),
    .B(_04090_),
    .X(_00812_));
 sg13g2_buf_1 fanout210 (.A(net245),
    .X(net210));
 sg13g2_mux2_1 _10171_ (.A0(\shift_storage.storage[19] ),
    .A1(\shift_storage.storage[18] ),
    .S(net615),
    .X(_04092_));
 sg13g2_and2_1 _10172_ (.A(net316),
    .B(_04092_),
    .X(_00813_));
 sg13g2_mux2_1 _10173_ (.A0(\shift_storage.storage[1] ),
    .A1(\shift_storage.storage[0] ),
    .S(net612),
    .X(_04093_));
 sg13g2_and2_1 _10174_ (.A(net314),
    .B(_04093_),
    .X(_00814_));
 sg13g2_mux2_1 _10175_ (.A0(\shift_storage.storage[200] ),
    .A1(\shift_storage.storage[199] ),
    .S(net599),
    .X(_04094_));
 sg13g2_and2_1 _10176_ (.A(net301),
    .B(_04094_),
    .X(_00815_));
 sg13g2_buf_2 fanout209 (.A(net210),
    .X(net209));
 sg13g2_mux2_1 _10178_ (.A0(\shift_storage.storage[201] ),
    .A1(\shift_storage.storage[200] ),
    .S(net599),
    .X(_04096_));
 sg13g2_and2_1 _10179_ (.A(net301),
    .B(_04096_),
    .X(_00816_));
 sg13g2_mux2_1 _10180_ (.A0(\shift_storage.storage[202] ),
    .A1(\shift_storage.storage[201] ),
    .S(net604),
    .X(_04097_));
 sg13g2_and2_1 _10181_ (.A(net307),
    .B(_04097_),
    .X(_00817_));
 sg13g2_mux2_1 _10182_ (.A0(\shift_storage.storage[203] ),
    .A1(\shift_storage.storage[202] ),
    .S(net604),
    .X(_04098_));
 sg13g2_and2_1 _10183_ (.A(net307),
    .B(_04098_),
    .X(_00818_));
 sg13g2_mux2_1 _10184_ (.A0(\shift_storage.storage[204] ),
    .A1(\shift_storage.storage[203] ),
    .S(net604),
    .X(_04099_));
 sg13g2_and2_1 _10185_ (.A(net307),
    .B(_04099_),
    .X(_00819_));
 sg13g2_mux2_1 _10186_ (.A0(\shift_storage.storage[205] ),
    .A1(\shift_storage.storage[204] ),
    .S(net604),
    .X(_04100_));
 sg13g2_and2_1 _10187_ (.A(net307),
    .B(_04100_),
    .X(_00820_));
 sg13g2_mux2_1 _10188_ (.A0(\shift_storage.storage[206] ),
    .A1(\shift_storage.storage[205] ),
    .S(net596),
    .X(_04101_));
 sg13g2_and2_1 _10189_ (.A(net297),
    .B(_04101_),
    .X(_00821_));
 sg13g2_mux2_1 _10190_ (.A0(\shift_storage.storage[207] ),
    .A1(\shift_storage.storage[206] ),
    .S(net596),
    .X(_04102_));
 sg13g2_and2_1 _10191_ (.A(net298),
    .B(_04102_),
    .X(_00822_));
 sg13g2_buf_2 fanout208 (.A(net209),
    .X(net208));
 sg13g2_mux2_1 _10193_ (.A0(\shift_storage.storage[208] ),
    .A1(\shift_storage.storage[207] ),
    .S(net595),
    .X(_04104_));
 sg13g2_and2_1 _10194_ (.A(net297),
    .B(_04104_),
    .X(_00823_));
 sg13g2_mux2_1 _10195_ (.A0(\shift_storage.storage[209] ),
    .A1(\shift_storage.storage[208] ),
    .S(net595),
    .X(_04105_));
 sg13g2_and2_1 _10196_ (.A(net297),
    .B(_04105_),
    .X(_00824_));
 sg13g2_mux2_1 _10197_ (.A0(\shift_storage.storage[20] ),
    .A1(\shift_storage.storage[19] ),
    .S(net615),
    .X(_04106_));
 sg13g2_and2_1 _10198_ (.A(net317),
    .B(_04106_),
    .X(_00825_));
 sg13g2_buf_1 fanout207 (.A(net210),
    .X(net207));
 sg13g2_mux2_1 _10200_ (.A0(\shift_storage.storage[210] ),
    .A1(\shift_storage.storage[209] ),
    .S(net595),
    .X(_04108_));
 sg13g2_and2_1 _10201_ (.A(net297),
    .B(_04108_),
    .X(_00826_));
 sg13g2_mux2_1 _10202_ (.A0(\shift_storage.storage[211] ),
    .A1(\shift_storage.storage[210] ),
    .S(net595),
    .X(_04109_));
 sg13g2_and2_1 _10203_ (.A(net297),
    .B(_04109_),
    .X(_00827_));
 sg13g2_mux2_1 _10204_ (.A0(\shift_storage.storage[212] ),
    .A1(\shift_storage.storage[211] ),
    .S(net595),
    .X(_04110_));
 sg13g2_and2_1 _10205_ (.A(net297),
    .B(_04110_),
    .X(_00828_));
 sg13g2_mux2_1 _10206_ (.A0(\shift_storage.storage[213] ),
    .A1(\shift_storage.storage[212] ),
    .S(net595),
    .X(_04111_));
 sg13g2_and2_1 _10207_ (.A(net293),
    .B(_04111_),
    .X(_00829_));
 sg13g2_mux2_1 _10208_ (.A0(\shift_storage.storage[214] ),
    .A1(\shift_storage.storage[213] ),
    .S(net592),
    .X(_04112_));
 sg13g2_and2_1 _10209_ (.A(net293),
    .B(_04112_),
    .X(_00830_));
 sg13g2_mux2_1 _10210_ (.A0(\shift_storage.storage[215] ),
    .A1(\shift_storage.storage[214] ),
    .S(net592),
    .X(_04113_));
 sg13g2_and2_1 _10211_ (.A(net293),
    .B(_04113_),
    .X(_00831_));
 sg13g2_mux2_1 _10212_ (.A0(\shift_storage.storage[216] ),
    .A1(\shift_storage.storage[215] ),
    .S(net592),
    .X(_04114_));
 sg13g2_and2_1 _10213_ (.A(net293),
    .B(_04114_),
    .X(_00832_));
 sg13g2_buf_1 fanout206 (.A(net207),
    .X(net206));
 sg13g2_mux2_1 _10215_ (.A0(\shift_storage.storage[217] ),
    .A1(\shift_storage.storage[216] ),
    .S(net592),
    .X(_04116_));
 sg13g2_and2_1 _10216_ (.A(net293),
    .B(_04116_),
    .X(_00833_));
 sg13g2_mux2_1 _10217_ (.A0(\shift_storage.storage[218] ),
    .A1(\shift_storage.storage[217] ),
    .S(net592),
    .X(_04117_));
 sg13g2_and2_1 _10218_ (.A(net293),
    .B(_04117_),
    .X(_00834_));
 sg13g2_mux2_1 _10219_ (.A0(\shift_storage.storage[219] ),
    .A1(\shift_storage.storage[218] ),
    .S(net591),
    .X(_04118_));
 sg13g2_and2_1 _10220_ (.A(net292),
    .B(_04118_),
    .X(_00835_));
 sg13g2_buf_1 fanout205 (.A(net207),
    .X(net205));
 sg13g2_mux2_1 _10222_ (.A0(\shift_storage.storage[21] ),
    .A1(\shift_storage.storage[20] ),
    .S(net614),
    .X(_04120_));
 sg13g2_and2_1 _10223_ (.A(net316),
    .B(_04120_),
    .X(_00836_));
 sg13g2_mux2_1 _10224_ (.A0(\shift_storage.storage[220] ),
    .A1(\shift_storage.storage[219] ),
    .S(net591),
    .X(_04121_));
 sg13g2_and2_1 _10225_ (.A(net292),
    .B(_04121_),
    .X(_00837_));
 sg13g2_mux2_1 _10226_ (.A0(\shift_storage.storage[221] ),
    .A1(\shift_storage.storage[220] ),
    .S(net591),
    .X(_04122_));
 sg13g2_and2_1 _10227_ (.A(net292),
    .B(_04122_),
    .X(_00838_));
 sg13g2_mux2_1 _10228_ (.A0(\shift_storage.storage[222] ),
    .A1(\shift_storage.storage[221] ),
    .S(net591),
    .X(_04123_));
 sg13g2_and2_1 _10229_ (.A(net290),
    .B(_04123_),
    .X(_00839_));
 sg13g2_mux2_1 _10230_ (.A0(\shift_storage.storage[223] ),
    .A1(\shift_storage.storage[222] ),
    .S(net591),
    .X(_04124_));
 sg13g2_and2_1 _10231_ (.A(net292),
    .B(_04124_),
    .X(_00840_));
 sg13g2_mux2_1 _10232_ (.A0(\shift_storage.storage[224] ),
    .A1(\shift_storage.storage[223] ),
    .S(net591),
    .X(_04125_));
 sg13g2_and2_1 _10233_ (.A(net292),
    .B(_04125_),
    .X(_00841_));
 sg13g2_mux2_1 _10234_ (.A0(\shift_storage.storage[225] ),
    .A1(\shift_storage.storage[224] ),
    .S(net533),
    .X(_04126_));
 sg13g2_and2_1 _10235_ (.A(net232),
    .B(_04126_),
    .X(_00842_));
 sg13g2_buf_2 fanout204 (.A(net207),
    .X(net204));
 sg13g2_mux2_1 _10237_ (.A0(\shift_storage.storage[226] ),
    .A1(\shift_storage.storage[225] ),
    .S(net533),
    .X(_04128_));
 sg13g2_and2_1 _10238_ (.A(net232),
    .B(_04128_),
    .X(_00843_));
 sg13g2_mux2_1 _10239_ (.A0(\shift_storage.storage[227] ),
    .A1(\shift_storage.storage[226] ),
    .S(net533),
    .X(_04129_));
 sg13g2_and2_1 _10240_ (.A(net232),
    .B(_04129_),
    .X(_00844_));
 sg13g2_mux2_1 _10241_ (.A0(\shift_storage.storage[228] ),
    .A1(\shift_storage.storage[227] ),
    .S(net533),
    .X(_04130_));
 sg13g2_and2_1 _10242_ (.A(net232),
    .B(_04130_),
    .X(_00845_));
 sg13g2_buf_1 fanout203 (.A(_03207_),
    .X(net203));
 sg13g2_mux2_1 _10244_ (.A0(\shift_storage.storage[229] ),
    .A1(\shift_storage.storage[228] ),
    .S(net533),
    .X(_04132_));
 sg13g2_and2_1 _10245_ (.A(net232),
    .B(_04132_),
    .X(_00846_));
 sg13g2_mux2_1 _10246_ (.A0(\shift_storage.storage[22] ),
    .A1(\shift_storage.storage[21] ),
    .S(net604),
    .X(_04133_));
 sg13g2_and2_1 _10247_ (.A(net308),
    .B(_04133_),
    .X(_00847_));
 sg13g2_mux2_1 _10248_ (.A0(\shift_storage.storage[230] ),
    .A1(\shift_storage.storage[229] ),
    .S(net533),
    .X(_04134_));
 sg13g2_and2_1 _10249_ (.A(net232),
    .B(_04134_),
    .X(_00848_));
 sg13g2_mux2_1 _10250_ (.A0(\shift_storage.storage[231] ),
    .A1(\shift_storage.storage[230] ),
    .S(net531),
    .X(_04135_));
 sg13g2_and2_1 _10251_ (.A(net230),
    .B(_04135_),
    .X(_00849_));
 sg13g2_mux2_1 _10252_ (.A0(\shift_storage.storage[232] ),
    .A1(\shift_storage.storage[231] ),
    .S(net531),
    .X(_04136_));
 sg13g2_and2_1 _10253_ (.A(net230),
    .B(_04136_),
    .X(_00850_));
 sg13g2_mux2_1 _10254_ (.A0(\shift_storage.storage[233] ),
    .A1(\shift_storage.storage[232] ),
    .S(net532),
    .X(_04137_));
 sg13g2_and2_1 _10255_ (.A(net230),
    .B(_04137_),
    .X(_00851_));
 sg13g2_mux2_1 _10256_ (.A0(\shift_storage.storage[234] ),
    .A1(\shift_storage.storage[233] ),
    .S(net532),
    .X(_04138_));
 sg13g2_and2_1 _10257_ (.A(net230),
    .B(_04138_),
    .X(_00852_));
 sg13g2_buf_2 fanout202 (.A(net203),
    .X(net202));
 sg13g2_mux2_1 _10259_ (.A0(\shift_storage.storage[235] ),
    .A1(\shift_storage.storage[234] ),
    .S(net531),
    .X(_04140_));
 sg13g2_and2_1 _10260_ (.A(net231),
    .B(_04140_),
    .X(_00853_));
 sg13g2_mux2_1 _10261_ (.A0(\shift_storage.storage[236] ),
    .A1(\shift_storage.storage[235] ),
    .S(net531),
    .X(_04141_));
 sg13g2_and2_1 _10262_ (.A(net231),
    .B(_04141_),
    .X(_00854_));
 sg13g2_mux2_1 _10263_ (.A0(\shift_storage.storage[237] ),
    .A1(\shift_storage.storage[236] ),
    .S(net531),
    .X(_04142_));
 sg13g2_and2_1 _10264_ (.A(net231),
    .B(_04142_),
    .X(_00855_));
 sg13g2_buf_2 fanout201 (.A(net203),
    .X(net201));
 sg13g2_mux2_1 _10266_ (.A0(\shift_storage.storage[238] ),
    .A1(\shift_storage.storage[237] ),
    .S(net531),
    .X(_04144_));
 sg13g2_and2_1 _10267_ (.A(net231),
    .B(_04144_),
    .X(_00856_));
 sg13g2_mux2_1 _10268_ (.A0(\shift_storage.storage[239] ),
    .A1(\shift_storage.storage[238] ),
    .S(net531),
    .X(_04145_));
 sg13g2_and2_1 _10269_ (.A(net231),
    .B(_04145_),
    .X(_00857_));
 sg13g2_mux2_1 _10270_ (.A0(\shift_storage.storage[23] ),
    .A1(\shift_storage.storage[22] ),
    .S(net605),
    .X(_04146_));
 sg13g2_and2_1 _10271_ (.A(net306),
    .B(_04146_),
    .X(_00858_));
 sg13g2_mux2_1 _10272_ (.A0(\shift_storage.storage[240] ),
    .A1(\shift_storage.storage[239] ),
    .S(net531),
    .X(_04147_));
 sg13g2_and2_1 _10273_ (.A(net231),
    .B(_04147_),
    .X(_00859_));
 sg13g2_mux2_1 _10274_ (.A0(\shift_storage.storage[241] ),
    .A1(\shift_storage.storage[240] ),
    .S(net589),
    .X(_04148_));
 sg13g2_and2_1 _10275_ (.A(net290),
    .B(_04148_),
    .X(_00860_));
 sg13g2_mux2_1 _10276_ (.A0(\shift_storage.storage[242] ),
    .A1(\shift_storage.storage[241] ),
    .S(net589),
    .X(_04149_));
 sg13g2_and2_1 _10277_ (.A(net290),
    .B(_04149_),
    .X(_00861_));
 sg13g2_mux2_1 _10278_ (.A0(\shift_storage.storage[243] ),
    .A1(\shift_storage.storage[242] ),
    .S(net589),
    .X(_04150_));
 sg13g2_and2_1 _10279_ (.A(net290),
    .B(_04150_),
    .X(_00862_));
 sg13g2_buf_1 fanout200 (.A(_03207_),
    .X(net200));
 sg13g2_mux2_1 _10281_ (.A0(\shift_storage.storage[244] ),
    .A1(\shift_storage.storage[243] ),
    .S(net589),
    .X(_04152_));
 sg13g2_and2_1 _10282_ (.A(net290),
    .B(_04152_),
    .X(_00863_));
 sg13g2_mux2_1 _10283_ (.A0(\shift_storage.storage[245] ),
    .A1(\shift_storage.storage[244] ),
    .S(net589),
    .X(_04153_));
 sg13g2_and2_1 _10284_ (.A(net290),
    .B(_04153_),
    .X(_00864_));
 sg13g2_mux2_1 _10285_ (.A0(\shift_storage.storage[246] ),
    .A1(\shift_storage.storage[245] ),
    .S(net589),
    .X(_04154_));
 sg13g2_and2_1 _10286_ (.A(net290),
    .B(_04154_),
    .X(_00865_));
 sg13g2_buf_2 fanout199 (.A(net200),
    .X(net199));
 sg13g2_mux2_1 _10288_ (.A0(\shift_storage.storage[247] ),
    .A1(\shift_storage.storage[246] ),
    .S(net589),
    .X(_04156_));
 sg13g2_and2_1 _10289_ (.A(net290),
    .B(_04156_),
    .X(_00866_));
 sg13g2_mux2_1 _10290_ (.A0(\shift_storage.storage[248] ),
    .A1(\shift_storage.storage[247] ),
    .S(net590),
    .X(_04157_));
 sg13g2_and2_1 _10291_ (.A(net291),
    .B(_04157_),
    .X(_00867_));
 sg13g2_mux2_1 _10292_ (.A0(\shift_storage.storage[249] ),
    .A1(\shift_storage.storage[248] ),
    .S(net590),
    .X(_04158_));
 sg13g2_and2_1 _10293_ (.A(net291),
    .B(_04158_),
    .X(_00868_));
 sg13g2_mux2_1 _10294_ (.A0(\shift_storage.storage[24] ),
    .A1(\shift_storage.storage[23] ),
    .S(net605),
    .X(_04159_));
 sg13g2_and2_1 _10295_ (.A(net306),
    .B(_04159_),
    .X(_00869_));
 sg13g2_mux2_1 _10296_ (.A0(\shift_storage.storage[250] ),
    .A1(\shift_storage.storage[249] ),
    .S(net590),
    .X(_04160_));
 sg13g2_and2_1 _10297_ (.A(net291),
    .B(_04160_),
    .X(_00870_));
 sg13g2_mux2_1 _10298_ (.A0(\shift_storage.storage[251] ),
    .A1(\shift_storage.storage[250] ),
    .S(net590),
    .X(_04161_));
 sg13g2_and2_1 _10299_ (.A(net291),
    .B(_04161_),
    .X(_00871_));
 sg13g2_mux2_1 _10300_ (.A0(\shift_storage.storage[252] ),
    .A1(\shift_storage.storage[251] ),
    .S(net590),
    .X(_04162_));
 sg13g2_and2_1 _10301_ (.A(net291),
    .B(_04162_),
    .X(_00872_));
 sg13g2_buf_2 fanout198 (.A(_05183_),
    .X(net198));
 sg13g2_buf_1 fanout197 (.A(\median_processor.input_storage[0] ),
    .X(net197));
 sg13g2_mux2_1 _10304_ (.A0(\shift_storage.storage[253] ),
    .A1(\shift_storage.storage[252] ),
    .S(net590),
    .X(_04165_));
 sg13g2_and2_1 _10305_ (.A(net291),
    .B(_04165_),
    .X(_00873_));
 sg13g2_mux2_1 _10306_ (.A0(\shift_storage.storage[254] ),
    .A1(\shift_storage.storage[253] ),
    .S(net589),
    .X(_04166_));
 sg13g2_and2_1 _10307_ (.A(net291),
    .B(_04166_),
    .X(_00874_));
 sg13g2_mux2_1 _10308_ (.A0(\shift_storage.storage[255] ),
    .A1(\shift_storage.storage[254] ),
    .S(net590),
    .X(_04167_));
 sg13g2_and2_1 _10309_ (.A(net291),
    .B(_04167_),
    .X(_00875_));
 sg13g2_buf_2 fanout196 (.A(net197),
    .X(net196));
 sg13g2_buf_1 fanout195 (.A(\median_processor.input_storage[10] ),
    .X(net195));
 sg13g2_mux2_1 _10312_ (.A0(\shift_storage.storage[256] ),
    .A1(\shift_storage.storage[255] ),
    .S(net593),
    .X(_04170_));
 sg13g2_and2_1 _10313_ (.A(net295),
    .B(_04170_),
    .X(_00876_));
 sg13g2_mux2_1 _10314_ (.A0(\shift_storage.storage[257] ),
    .A1(\shift_storage.storage[256] ),
    .S(net593),
    .X(_04171_));
 sg13g2_and2_1 _10315_ (.A(net295),
    .B(_04171_),
    .X(_00877_));
 sg13g2_mux2_1 _10316_ (.A0(\shift_storage.storage[258] ),
    .A1(\shift_storage.storage[257] ),
    .S(net593),
    .X(_04172_));
 sg13g2_and2_1 _10317_ (.A(net295),
    .B(_04172_),
    .X(_00878_));
 sg13g2_mux2_1 _10318_ (.A0(\shift_storage.storage[259] ),
    .A1(\shift_storage.storage[258] ),
    .S(net593),
    .X(_04173_));
 sg13g2_and2_1 _10319_ (.A(net295),
    .B(_04173_),
    .X(_00879_));
 sg13g2_mux2_1 _10320_ (.A0(\shift_storage.storage[25] ),
    .A1(\shift_storage.storage[24] ),
    .S(net605),
    .X(_04174_));
 sg13g2_and2_1 _10321_ (.A(net306),
    .B(_04174_),
    .X(_00880_));
 sg13g2_mux2_1 _10322_ (.A0(\shift_storage.storage[260] ),
    .A1(\shift_storage.storage[259] ),
    .S(net593),
    .X(_04175_));
 sg13g2_and2_1 _10323_ (.A(net295),
    .B(_04175_),
    .X(_00881_));
 sg13g2_mux2_1 _10324_ (.A0(\shift_storage.storage[261] ),
    .A1(\shift_storage.storage[260] ),
    .S(net593),
    .X(_04176_));
 sg13g2_and2_1 _10325_ (.A(net295),
    .B(_04176_),
    .X(_00882_));
 sg13g2_buf_2 fanout194 (.A(\median_processor.input_storage[10] ),
    .X(net194));
 sg13g2_mux2_1 _10327_ (.A0(\shift_storage.storage[262] ),
    .A1(\shift_storage.storage[261] ),
    .S(net593),
    .X(_04178_));
 sg13g2_and2_1 _10328_ (.A(net296),
    .B(_04178_),
    .X(_00883_));
 sg13g2_mux2_1 _10329_ (.A0(\shift_storage.storage[263] ),
    .A1(\shift_storage.storage[262] ),
    .S(net594),
    .X(_04179_));
 sg13g2_and2_1 _10330_ (.A(net295),
    .B(_04179_),
    .X(_00884_));
 sg13g2_mux2_1 _10331_ (.A0(\shift_storage.storage[264] ),
    .A1(\shift_storage.storage[263] ),
    .S(net593),
    .X(_04180_));
 sg13g2_and2_1 _10332_ (.A(net295),
    .B(_04180_),
    .X(_00885_));
 sg13g2_buf_1 fanout193 (.A(\median_processor.input_storage[11] ),
    .X(net193));
 sg13g2_mux2_1 _10334_ (.A0(\shift_storage.storage[265] ),
    .A1(\shift_storage.storage[264] ),
    .S(net594),
    .X(_04182_));
 sg13g2_and2_1 _10335_ (.A(net296),
    .B(_04182_),
    .X(_00886_));
 sg13g2_mux2_1 _10336_ (.A0(\shift_storage.storage[266] ),
    .A1(\shift_storage.storage[265] ),
    .S(net594),
    .X(_04183_));
 sg13g2_and2_1 _10337_ (.A(net296),
    .B(_04183_),
    .X(_00887_));
 sg13g2_mux2_1 _10338_ (.A0(\shift_storage.storage[267] ),
    .A1(\shift_storage.storage[266] ),
    .S(net594),
    .X(_04184_));
 sg13g2_and2_1 _10339_ (.A(net296),
    .B(_04184_),
    .X(_00888_));
 sg13g2_mux2_1 _10340_ (.A0(\shift_storage.storage[268] ),
    .A1(\shift_storage.storage[267] ),
    .S(net596),
    .X(_04185_));
 sg13g2_and2_1 _10341_ (.A(net298),
    .B(_04185_),
    .X(_00889_));
 sg13g2_mux2_1 _10342_ (.A0(\shift_storage.storage[269] ),
    .A1(\shift_storage.storage[268] ),
    .S(net609),
    .X(_04186_));
 sg13g2_and2_1 _10343_ (.A(net312),
    .B(_04186_),
    .X(_00890_));
 sg13g2_mux2_1 _10344_ (.A0(\shift_storage.storage[26] ),
    .A1(\shift_storage.storage[25] ),
    .S(net606),
    .X(_04187_));
 sg13g2_and2_1 _10345_ (.A(net306),
    .B(_04187_),
    .X(_00891_));
 sg13g2_mux2_1 _10346_ (.A0(\shift_storage.storage[270] ),
    .A1(\shift_storage.storage[269] ),
    .S(net609),
    .X(_04188_));
 sg13g2_and2_1 _10347_ (.A(net312),
    .B(_04188_),
    .X(_00892_));
 sg13g2_buf_1 fanout192 (.A(net193),
    .X(net192));
 sg13g2_mux2_1 _10349_ (.A0(\shift_storage.storage[271] ),
    .A1(\shift_storage.storage[270] ),
    .S(net608),
    .X(_04190_));
 sg13g2_and2_1 _10350_ (.A(net310),
    .B(_04190_),
    .X(_00893_));
 sg13g2_mux2_1 _10351_ (.A0(\shift_storage.storage[272] ),
    .A1(\shift_storage.storage[271] ),
    .S(net608),
    .X(_04191_));
 sg13g2_and2_1 _10352_ (.A(net310),
    .B(_04191_),
    .X(_00894_));
 sg13g2_mux2_1 _10353_ (.A0(\shift_storage.storage[273] ),
    .A1(\shift_storage.storage[272] ),
    .S(net608),
    .X(_04192_));
 sg13g2_and2_1 _10354_ (.A(net310),
    .B(_04192_),
    .X(_00895_));
 sg13g2_buf_2 fanout191 (.A(net193),
    .X(net191));
 sg13g2_mux2_1 _10356_ (.A0(\shift_storage.storage[274] ),
    .A1(\shift_storage.storage[273] ),
    .S(net608),
    .X(_04194_));
 sg13g2_and2_1 _10357_ (.A(net310),
    .B(_04194_),
    .X(_00896_));
 sg13g2_mux2_1 _10358_ (.A0(\shift_storage.storage[275] ),
    .A1(\shift_storage.storage[274] ),
    .S(net608),
    .X(_04195_));
 sg13g2_and2_1 _10359_ (.A(net310),
    .B(_04195_),
    .X(_00897_));
 sg13g2_mux2_1 _10360_ (.A0(\shift_storage.storage[276] ),
    .A1(\shift_storage.storage[275] ),
    .S(net611),
    .X(_04196_));
 sg13g2_and2_1 _10361_ (.A(net313),
    .B(_04196_),
    .X(_00898_));
 sg13g2_mux2_1 _10362_ (.A0(\shift_storage.storage[277] ),
    .A1(\shift_storage.storage[276] ),
    .S(net608),
    .X(_04197_));
 sg13g2_and2_1 _10363_ (.A(net310),
    .B(_04197_),
    .X(_00899_));
 sg13g2_mux2_1 _10364_ (.A0(\shift_storage.storage[278] ),
    .A1(\shift_storage.storage[277] ),
    .S(net612),
    .X(_04198_));
 sg13g2_and2_1 _10365_ (.A(net314),
    .B(_04198_),
    .X(_00900_));
 sg13g2_mux2_1 _10366_ (.A0(\shift_storage.storage[279] ),
    .A1(\shift_storage.storage[278] ),
    .S(net612),
    .X(_04199_));
 sg13g2_and2_1 _10367_ (.A(net314),
    .B(_04199_),
    .X(_00901_));
 sg13g2_mux2_1 _10368_ (.A0(\shift_storage.storage[27] ),
    .A1(\shift_storage.storage[26] ),
    .S(net606),
    .X(_04200_));
 sg13g2_and2_1 _10369_ (.A(net308),
    .B(_04200_),
    .X(_00902_));
 sg13g2_buf_2 fanout190 (.A(\median_processor.input_storage[12] ),
    .X(net190));
 sg13g2_mux2_1 _10371_ (.A0(\shift_storage.storage[280] ),
    .A1(\shift_storage.storage[279] ),
    .S(net613),
    .X(_04202_));
 sg13g2_and2_1 _10372_ (.A(net315),
    .B(_04202_),
    .X(_00903_));
 sg13g2_mux2_1 _10373_ (.A0(\shift_storage.storage[281] ),
    .A1(\shift_storage.storage[280] ),
    .S(net613),
    .X(_04203_));
 sg13g2_and2_1 _10374_ (.A(net315),
    .B(_04203_),
    .X(_00904_));
 sg13g2_mux2_1 _10375_ (.A0(\shift_storage.storage[282] ),
    .A1(\shift_storage.storage[281] ),
    .S(net613),
    .X(_04204_));
 sg13g2_and2_1 _10376_ (.A(net315),
    .B(_04204_),
    .X(_00905_));
 sg13g2_buf_2 fanout189 (.A(\median_processor.input_storage[12] ),
    .X(net189));
 sg13g2_mux2_1 _10378_ (.A0(\shift_storage.storage[283] ),
    .A1(\shift_storage.storage[282] ),
    .S(net609),
    .X(_04206_));
 sg13g2_and2_1 _10379_ (.A(net311),
    .B(_04206_),
    .X(_00906_));
 sg13g2_mux2_1 _10380_ (.A0(\shift_storage.storage[284] ),
    .A1(\shift_storage.storage[283] ),
    .S(net610),
    .X(_04207_));
 sg13g2_and2_1 _10381_ (.A(net311),
    .B(_04207_),
    .X(_00907_));
 sg13g2_mux2_1 _10382_ (.A0(\shift_storage.storage[285] ),
    .A1(\shift_storage.storage[284] ),
    .S(net616),
    .X(_04208_));
 sg13g2_and2_1 _10383_ (.A(net311),
    .B(_04208_),
    .X(_00908_));
 sg13g2_mux2_1 _10384_ (.A0(\shift_storage.storage[286] ),
    .A1(\shift_storage.storage[285] ),
    .S(net616),
    .X(_04209_));
 sg13g2_and2_1 _10385_ (.A(net317),
    .B(_04209_),
    .X(_00909_));
 sg13g2_mux2_1 _10386_ (.A0(\shift_storage.storage[287] ),
    .A1(\shift_storage.storage[286] ),
    .S(net617),
    .X(_04210_));
 sg13g2_and2_1 _10387_ (.A(net319),
    .B(_04210_),
    .X(_00910_));
 sg13g2_mux2_1 _10388_ (.A0(\shift_storage.storage[288] ),
    .A1(\shift_storage.storage[287] ),
    .S(net617),
    .X(_04211_));
 sg13g2_and2_1 _10389_ (.A(net319),
    .B(_04211_),
    .X(_00911_));
 sg13g2_mux2_1 _10390_ (.A0(\shift_storage.storage[289] ),
    .A1(\shift_storage.storage[288] ),
    .S(net617),
    .X(_04212_));
 sg13g2_and2_1 _10391_ (.A(net319),
    .B(_04212_),
    .X(_00912_));
 sg13g2_buf_2 fanout188 (.A(\median_processor.input_storage[13] ),
    .X(net188));
 sg13g2_mux2_1 _10393_ (.A0(\shift_storage.storage[28] ),
    .A1(\shift_storage.storage[27] ),
    .S(net606),
    .X(_04214_));
 sg13g2_and2_1 _10394_ (.A(net308),
    .B(_04214_),
    .X(_00913_));
 sg13g2_mux2_1 _10395_ (.A0(\shift_storage.storage[290] ),
    .A1(\shift_storage.storage[289] ),
    .S(net617),
    .X(_04215_));
 sg13g2_and2_1 _10396_ (.A(net319),
    .B(_04215_),
    .X(_00914_));
 sg13g2_mux2_1 _10397_ (.A0(\shift_storage.storage[291] ),
    .A1(\shift_storage.storage[290] ),
    .S(net617),
    .X(_04216_));
 sg13g2_and2_1 _10398_ (.A(net319),
    .B(_04216_),
    .X(_00915_));
 sg13g2_buf_2 fanout187 (.A(net188),
    .X(net187));
 sg13g2_mux2_1 _10400_ (.A0(\shift_storage.storage[292] ),
    .A1(\shift_storage.storage[291] ),
    .S(net616),
    .X(_04218_));
 sg13g2_and2_1 _10401_ (.A(net318),
    .B(_04218_),
    .X(_00916_));
 sg13g2_mux2_1 _10402_ (.A0(\shift_storage.storage[293] ),
    .A1(\shift_storage.storage[292] ),
    .S(net616),
    .X(_04219_));
 sg13g2_and2_1 _10403_ (.A(net318),
    .B(_04219_),
    .X(_00917_));
 sg13g2_mux2_1 _10404_ (.A0(\shift_storage.storage[294] ),
    .A1(\shift_storage.storage[293] ),
    .S(net616),
    .X(_04220_));
 sg13g2_and2_1 _10405_ (.A(net318),
    .B(_04220_),
    .X(_00918_));
 sg13g2_mux2_1 _10406_ (.A0(\shift_storage.storage[295] ),
    .A1(\shift_storage.storage[294] ),
    .S(net615),
    .X(_04221_));
 sg13g2_and2_1 _10407_ (.A(net317),
    .B(_04221_),
    .X(_00919_));
 sg13g2_mux2_1 _10408_ (.A0(\shift_storage.storage[296] ),
    .A1(\shift_storage.storage[295] ),
    .S(net616),
    .X(_04222_));
 sg13g2_and2_1 _10409_ (.A(net317),
    .B(_04222_),
    .X(_00920_));
 sg13g2_mux2_1 _10410_ (.A0(\shift_storage.storage[297] ),
    .A1(\shift_storage.storage[296] ),
    .S(net615),
    .X(_04223_));
 sg13g2_and2_1 _10411_ (.A(net318),
    .B(_04223_),
    .X(_00921_));
 sg13g2_mux2_1 _10412_ (.A0(\shift_storage.storage[298] ),
    .A1(\shift_storage.storage[297] ),
    .S(net615),
    .X(_04224_));
 sg13g2_and2_1 _10413_ (.A(net317),
    .B(_04224_),
    .X(_00922_));
 sg13g2_buf_2 fanout186 (.A(net187),
    .X(net186));
 sg13g2_mux2_1 _10415_ (.A0(\shift_storage.storage[299] ),
    .A1(\shift_storage.storage[298] ),
    .S(net615),
    .X(_04226_));
 sg13g2_and2_1 _10416_ (.A(net317),
    .B(_04226_),
    .X(_00923_));
 sg13g2_mux2_1 _10417_ (.A0(\shift_storage.storage[29] ),
    .A1(\shift_storage.storage[28] ),
    .S(net606),
    .X(_04227_));
 sg13g2_and2_1 _10418_ (.A(net308),
    .B(_04227_),
    .X(_00924_));
 sg13g2_mux2_1 _10419_ (.A0(\shift_storage.storage[2] ),
    .A1(\shift_storage.storage[1] ),
    .S(net612),
    .X(_04228_));
 sg13g2_and2_1 _10420_ (.A(net314),
    .B(_04228_),
    .X(_00925_));
 sg13g2_buf_1 fanout185 (.A(\median_processor.input_storage[14] ),
    .X(net185));
 sg13g2_mux2_1 _10422_ (.A0(\shift_storage.storage[300] ),
    .A1(\shift_storage.storage[299] ),
    .S(net614),
    .X(_04230_));
 sg13g2_and2_1 _10423_ (.A(net312),
    .B(_04230_),
    .X(_00926_));
 sg13g2_mux2_1 _10424_ (.A0(\shift_storage.storage[301] ),
    .A1(\shift_storage.storage[300] ),
    .S(net609),
    .X(_04231_));
 sg13g2_and2_1 _10425_ (.A(net312),
    .B(_04231_),
    .X(_00927_));
 sg13g2_mux2_1 _10426_ (.A0(\shift_storage.storage[302] ),
    .A1(\shift_storage.storage[301] ),
    .S(net609),
    .X(_04232_));
 sg13g2_and2_1 _10427_ (.A(net312),
    .B(_04232_),
    .X(_00928_));
 sg13g2_mux2_1 _10428_ (.A0(\shift_storage.storage[303] ),
    .A1(\shift_storage.storage[302] ),
    .S(net614),
    .X(_04233_));
 sg13g2_and2_1 _10429_ (.A(net316),
    .B(_04233_),
    .X(_00929_));
 sg13g2_mux2_1 _10430_ (.A0(\shift_storage.storage[304] ),
    .A1(\shift_storage.storage[303] ),
    .S(net614),
    .X(_04234_));
 sg13g2_and2_1 _10431_ (.A(net316),
    .B(_04234_),
    .X(_00930_));
 sg13g2_mux2_1 _10432_ (.A0(\shift_storage.storage[305] ),
    .A1(\shift_storage.storage[304] ),
    .S(net614),
    .X(_04235_));
 sg13g2_and2_1 _10433_ (.A(net316),
    .B(_04235_),
    .X(_00931_));
 sg13g2_mux2_1 _10434_ (.A0(\shift_storage.storage[306] ),
    .A1(\shift_storage.storage[305] ),
    .S(net605),
    .X(_04236_));
 sg13g2_and2_1 _10435_ (.A(net306),
    .B(_04236_),
    .X(_00932_));
 sg13g2_buf_1 fanout184 (.A(net185),
    .X(net184));
 sg13g2_mux2_1 _10437_ (.A0(\shift_storage.storage[307] ),
    .A1(\shift_storage.storage[306] ),
    .S(net605),
    .X(_04238_));
 sg13g2_and2_1 _10438_ (.A(net306),
    .B(_04238_),
    .X(_00933_));
 sg13g2_mux2_1 _10439_ (.A0(\shift_storage.storage[308] ),
    .A1(\shift_storage.storage[307] ),
    .S(net605),
    .X(_04239_));
 sg13g2_and2_1 _10440_ (.A(net306),
    .B(_04239_),
    .X(_00934_));
 sg13g2_mux2_1 _10441_ (.A0(\shift_storage.storage[309] ),
    .A1(\shift_storage.storage[308] ),
    .S(net605),
    .X(_04240_));
 sg13g2_and2_1 _10442_ (.A(net306),
    .B(_04240_),
    .X(_00935_));
 sg13g2_buf_2 fanout183 (.A(net185),
    .X(net183));
 sg13g2_mux2_1 _10444_ (.A0(\shift_storage.storage[30] ),
    .A1(\shift_storage.storage[29] ),
    .S(net606),
    .X(_04242_));
 sg13g2_and2_1 _10445_ (.A(net308),
    .B(_04242_),
    .X(_00936_));
 sg13g2_mux2_1 _10446_ (.A0(\shift_storage.storage[310] ),
    .A1(\shift_storage.storage[309] ),
    .S(net604),
    .X(_04243_));
 sg13g2_and2_1 _10447_ (.A(net307),
    .B(_04243_),
    .X(_00937_));
 sg13g2_mux2_1 _10448_ (.A0(\shift_storage.storage[311] ),
    .A1(\shift_storage.storage[310] ),
    .S(net604),
    .X(_04244_));
 sg13g2_and2_1 _10449_ (.A(net307),
    .B(_04244_),
    .X(_00938_));
 sg13g2_mux2_1 _10450_ (.A0(\shift_storage.storage[312] ),
    .A1(\shift_storage.storage[311] ),
    .S(net604),
    .X(_04245_));
 sg13g2_and2_1 _10451_ (.A(net307),
    .B(_04245_),
    .X(_00939_));
 sg13g2_mux2_1 _10452_ (.A0(\shift_storage.storage[313] ),
    .A1(\shift_storage.storage[312] ),
    .S(net595),
    .X(_04246_));
 sg13g2_and2_1 _10453_ (.A(net298),
    .B(_04246_),
    .X(_00940_));
 sg13g2_mux2_1 _10454_ (.A0(\shift_storage.storage[314] ),
    .A1(\shift_storage.storage[313] ),
    .S(net596),
    .X(_04247_));
 sg13g2_and2_1 _10455_ (.A(net297),
    .B(_04247_),
    .X(_00941_));
 sg13g2_mux2_1 _10456_ (.A0(\shift_storage.storage[315] ),
    .A1(\shift_storage.storage[314] ),
    .S(net595),
    .X(_04248_));
 sg13g2_and2_1 _10457_ (.A(net297),
    .B(_04248_),
    .X(_00942_));
 sg13g2_buf_2 fanout182 (.A(\median_processor.input_storage[15] ),
    .X(net182));
 sg13g2_buf_2 fanout181 (.A(net182),
    .X(net181));
 sg13g2_mux2_1 _10460_ (.A0(\shift_storage.storage[316] ),
    .A1(\shift_storage.storage[315] ),
    .S(net599),
    .X(_04251_));
 sg13g2_and2_1 _10461_ (.A(net305),
    .B(_04251_),
    .X(_00943_));
 sg13g2_mux2_1 _10462_ (.A0(\shift_storage.storage[317] ),
    .A1(\shift_storage.storage[316] ),
    .S(net599),
    .X(_04252_));
 sg13g2_and2_1 _10463_ (.A(net305),
    .B(_04252_),
    .X(_00944_));
 sg13g2_mux2_1 _10464_ (.A0(\shift_storage.storage[318] ),
    .A1(\shift_storage.storage[317] ),
    .S(net599),
    .X(_04253_));
 sg13g2_and2_1 _10465_ (.A(net301),
    .B(_04253_),
    .X(_00945_));
 sg13g2_buf_2 fanout180 (.A(net182),
    .X(net180));
 sg13g2_buf_2 fanout179 (.A(\median_processor.input_storage[16] ),
    .X(net179));
 sg13g2_mux2_1 _10468_ (.A0(\shift_storage.storage[319] ),
    .A1(\shift_storage.storage[318] ),
    .S(net599),
    .X(_04256_));
 sg13g2_and2_1 _10469_ (.A(net293),
    .B(_04256_),
    .X(_00946_));
 sg13g2_mux2_1 _10470_ (.A0(\shift_storage.storage[31] ),
    .A1(\shift_storage.storage[30] ),
    .S(net606),
    .X(_04257_));
 sg13g2_and2_1 _10471_ (.A(net308),
    .B(_04257_),
    .X(_00947_));
 sg13g2_mux2_1 _10472_ (.A0(\shift_storage.storage[320] ),
    .A1(\shift_storage.storage[319] ),
    .S(net599),
    .X(_04258_));
 sg13g2_and2_1 _10473_ (.A(net293),
    .B(_04258_),
    .X(_00948_));
 sg13g2_mux2_1 _10474_ (.A0(\shift_storage.storage[321] ),
    .A1(\shift_storage.storage[320] ),
    .S(net598),
    .X(_04259_));
 sg13g2_and2_1 _10475_ (.A(net300),
    .B(_04259_),
    .X(_00949_));
 sg13g2_mux2_1 _10476_ (.A0(\shift_storage.storage[322] ),
    .A1(\shift_storage.storage[321] ),
    .S(net598),
    .X(_04260_));
 sg13g2_and2_1 _10477_ (.A(net300),
    .B(_04260_),
    .X(_00950_));
 sg13g2_mux2_1 _10478_ (.A0(\shift_storage.storage[323] ),
    .A1(\shift_storage.storage[322] ),
    .S(net598),
    .X(_04261_));
 sg13g2_and2_1 _10479_ (.A(net300),
    .B(_04261_),
    .X(_00951_));
 sg13g2_mux2_1 _10480_ (.A0(\shift_storage.storage[324] ),
    .A1(\shift_storage.storage[323] ),
    .S(net591),
    .X(_04262_));
 sg13g2_and2_1 _10481_ (.A(net292),
    .B(_04262_),
    .X(_00952_));
 sg13g2_buf_2 fanout178 (.A(net179),
    .X(net178));
 sg13g2_mux2_1 _10483_ (.A0(\shift_storage.storage[325] ),
    .A1(\shift_storage.storage[324] ),
    .S(net592),
    .X(_04264_));
 sg13g2_and2_1 _10484_ (.A(net292),
    .B(_04264_),
    .X(_00953_));
 sg13g2_mux2_1 _10485_ (.A0(\shift_storage.storage[326] ),
    .A1(\shift_storage.storage[325] ),
    .S(net591),
    .X(_04265_));
 sg13g2_and2_1 _10486_ (.A(net292),
    .B(_04265_),
    .X(_00954_));
 sg13g2_mux2_1 _10487_ (.A0(\shift_storage.storage[327] ),
    .A1(\shift_storage.storage[326] ),
    .S(net535),
    .X(_04266_));
 sg13g2_and2_1 _10488_ (.A(net234),
    .B(_04266_),
    .X(_00955_));
 sg13g2_buf_2 fanout177 (.A(\median_processor.input_storage[17] ),
    .X(net177));
 sg13g2_mux2_1 _10490_ (.A0(\shift_storage.storage[328] ),
    .A1(\shift_storage.storage[327] ),
    .S(net533),
    .X(_04268_));
 sg13g2_and2_1 _10491_ (.A(net232),
    .B(_04268_),
    .X(_00956_));
 sg13g2_mux2_1 _10492_ (.A0(\shift_storage.storage[329] ),
    .A1(\shift_storage.storage[328] ),
    .S(net535),
    .X(_04269_));
 sg13g2_and2_1 _10493_ (.A(net232),
    .B(_04269_),
    .X(_00957_));
 sg13g2_mux2_1 _10494_ (.A0(\shift_storage.storage[32] ),
    .A1(\shift_storage.storage[31] ),
    .S(net626),
    .X(_04270_));
 sg13g2_and2_1 _10495_ (.A(net328),
    .B(_04270_),
    .X(_00958_));
 sg13g2_mux2_1 _10496_ (.A0(\shift_storage.storage[330] ),
    .A1(\shift_storage.storage[329] ),
    .S(net533),
    .X(_04271_));
 sg13g2_and2_1 _10497_ (.A(net234),
    .B(_04271_),
    .X(_00959_));
 sg13g2_mux2_1 _10498_ (.A0(\shift_storage.storage[331] ),
    .A1(\shift_storage.storage[330] ),
    .S(net541),
    .X(_04272_));
 sg13g2_and2_1 _10499_ (.A(net240),
    .B(_04272_),
    .X(_00960_));
 sg13g2_mux2_1 _10500_ (.A0(\shift_storage.storage[332] ),
    .A1(\shift_storage.storage[331] ),
    .S(net541),
    .X(_04273_));
 sg13g2_and2_1 _10501_ (.A(net240),
    .B(_04273_),
    .X(_00961_));
 sg13g2_mux2_1 _10502_ (.A0(\shift_storage.storage[333] ),
    .A1(\shift_storage.storage[332] ),
    .S(net541),
    .X(_04274_));
 sg13g2_and2_1 _10503_ (.A(net241),
    .B(_04274_),
    .X(_00962_));
 sg13g2_buf_2 fanout176 (.A(\median_processor.input_storage[18] ),
    .X(net176));
 sg13g2_mux2_1 _10505_ (.A0(\shift_storage.storage[334] ),
    .A1(\shift_storage.storage[333] ),
    .S(net541),
    .X(_04276_));
 sg13g2_and2_1 _10506_ (.A(net240),
    .B(_04276_),
    .X(_00963_));
 sg13g2_mux2_1 _10507_ (.A0(\shift_storage.storage[335] ),
    .A1(\shift_storage.storage[334] ),
    .S(net540),
    .X(_04277_));
 sg13g2_and2_1 _10508_ (.A(net239),
    .B(_04277_),
    .X(_00964_));
 sg13g2_mux2_1 _10509_ (.A0(\shift_storage.storage[336] ),
    .A1(\shift_storage.storage[335] ),
    .S(net540),
    .X(_04278_));
 sg13g2_and2_1 _10510_ (.A(net239),
    .B(_04278_),
    .X(_00965_));
 sg13g2_buf_2 fanout175 (.A(net176),
    .X(net175));
 sg13g2_mux2_1 _10512_ (.A0(\shift_storage.storage[337] ),
    .A1(\shift_storage.storage[336] ),
    .S(net540),
    .X(_04280_));
 sg13g2_and2_1 _10513_ (.A(net233),
    .B(_04280_),
    .X(_00966_));
 sg13g2_mux2_1 _10514_ (.A0(\shift_storage.storage[338] ),
    .A1(\shift_storage.storage[337] ),
    .S(net534),
    .X(_04281_));
 sg13g2_and2_1 _10515_ (.A(net233),
    .B(_04281_),
    .X(_00967_));
 sg13g2_mux2_1 _10516_ (.A0(\shift_storage.storage[339] ),
    .A1(\shift_storage.storage[338] ),
    .S(net534),
    .X(_04282_));
 sg13g2_and2_1 _10517_ (.A(net233),
    .B(_04282_),
    .X(_00968_));
 sg13g2_mux2_1 _10518_ (.A0(\shift_storage.storage[33] ),
    .A1(\shift_storage.storage[32] ),
    .S(net626),
    .X(_04283_));
 sg13g2_and2_1 _10519_ (.A(net328),
    .B(_04283_),
    .X(_00969_));
 sg13g2_mux2_1 _10520_ (.A0(\shift_storage.storage[340] ),
    .A1(\shift_storage.storage[339] ),
    .S(net534),
    .X(_04284_));
 sg13g2_and2_1 _10521_ (.A(net233),
    .B(_04284_),
    .X(_00970_));
 sg13g2_mux2_1 _10522_ (.A0(\shift_storage.storage[341] ),
    .A1(\shift_storage.storage[340] ),
    .S(net534),
    .X(_04285_));
 sg13g2_and2_1 _10523_ (.A(net233),
    .B(_04285_),
    .X(_00971_));
 sg13g2_mux2_1 _10524_ (.A0(\shift_storage.storage[342] ),
    .A1(\shift_storage.storage[341] ),
    .S(net534),
    .X(_04286_));
 sg13g2_and2_1 _10525_ (.A(net233),
    .B(_04286_),
    .X(_00972_));
 sg13g2_buf_2 fanout174 (.A(\median_processor.input_storage[19] ),
    .X(net174));
 sg13g2_mux2_1 _10527_ (.A0(\shift_storage.storage[343] ),
    .A1(\shift_storage.storage[342] ),
    .S(net534),
    .X(_04288_));
 sg13g2_and2_1 _10528_ (.A(net230),
    .B(_04288_),
    .X(_00973_));
 sg13g2_mux2_1 _10529_ (.A0(\shift_storage.storage[344] ),
    .A1(\shift_storage.storage[343] ),
    .S(net532),
    .X(_04289_));
 sg13g2_and2_1 _10530_ (.A(net230),
    .B(_04289_),
    .X(_00974_));
 sg13g2_mux2_1 _10531_ (.A0(\shift_storage.storage[345] ),
    .A1(\shift_storage.storage[344] ),
    .S(net532),
    .X(_04290_));
 sg13g2_and2_1 _10532_ (.A(net230),
    .B(_04290_),
    .X(_00975_));
 sg13g2_buf_2 fanout173 (.A(net174),
    .X(net173));
 sg13g2_mux2_1 _10534_ (.A0(\shift_storage.storage[346] ),
    .A1(\shift_storage.storage[345] ),
    .S(net532),
    .X(_04292_));
 sg13g2_and2_1 _10535_ (.A(net230),
    .B(_04292_),
    .X(_00976_));
 sg13g2_mux2_1 _10536_ (.A0(\shift_storage.storage[347] ),
    .A1(\shift_storage.storage[346] ),
    .S(net527),
    .X(_04293_));
 sg13g2_and2_1 _10537_ (.A(net226),
    .B(_04293_),
    .X(_00977_));
 sg13g2_mux2_1 _10538_ (.A0(\shift_storage.storage[348] ),
    .A1(\shift_storage.storage[347] ),
    .S(net530),
    .X(_04294_));
 sg13g2_and2_1 _10539_ (.A(net229),
    .B(_04294_),
    .X(_00978_));
 sg13g2_mux2_1 _10540_ (.A0(\shift_storage.storage[349] ),
    .A1(\shift_storage.storage[348] ),
    .S(net527),
    .X(_04295_));
 sg13g2_and2_1 _10541_ (.A(net229),
    .B(_04295_),
    .X(_00979_));
 sg13g2_mux2_1 _10542_ (.A0(\shift_storage.storage[34] ),
    .A1(\shift_storage.storage[33] ),
    .S(net629),
    .X(_04296_));
 sg13g2_and2_1 _10543_ (.A(net331),
    .B(_04296_),
    .X(_00980_));
 sg13g2_mux2_1 _10544_ (.A0(\shift_storage.storage[350] ),
    .A1(\shift_storage.storage[349] ),
    .S(net530),
    .X(_04297_));
 sg13g2_and2_1 _10545_ (.A(net226),
    .B(_04297_),
    .X(_00981_));
 sg13g2_mux2_1 _10546_ (.A0(\shift_storage.storage[351] ),
    .A1(\shift_storage.storage[350] ),
    .S(net527),
    .X(_04298_));
 sg13g2_and2_1 _10547_ (.A(net226),
    .B(_04298_),
    .X(_00982_));
 sg13g2_buf_1 fanout172 (.A(\median_processor.input_storage[20] ),
    .X(net172));
 sg13g2_mux2_1 _10549_ (.A0(\shift_storage.storage[352] ),
    .A1(\shift_storage.storage[351] ),
    .S(net527),
    .X(_04300_));
 sg13g2_and2_1 _10550_ (.A(net226),
    .B(_04300_),
    .X(_00983_));
 sg13g2_mux2_1 _10551_ (.A0(\shift_storage.storage[353] ),
    .A1(\shift_storage.storage[352] ),
    .S(net527),
    .X(_04301_));
 sg13g2_and2_1 _10552_ (.A(net226),
    .B(_04301_),
    .X(_00984_));
 sg13g2_mux2_1 _10553_ (.A0(\shift_storage.storage[354] ),
    .A1(\shift_storage.storage[353] ),
    .S(net527),
    .X(_04302_));
 sg13g2_and2_1 _10554_ (.A(net226),
    .B(_04302_),
    .X(_00985_));
 sg13g2_buf_2 fanout171 (.A(\median_processor.input_storage[20] ),
    .X(net171));
 sg13g2_mux2_1 _10556_ (.A0(\shift_storage.storage[355] ),
    .A1(\shift_storage.storage[354] ),
    .S(net527),
    .X(_04304_));
 sg13g2_and2_1 _10557_ (.A(net226),
    .B(_04304_),
    .X(_00986_));
 sg13g2_mux2_1 _10558_ (.A0(\shift_storage.storage[356] ),
    .A1(\shift_storage.storage[355] ),
    .S(net527),
    .X(_04305_));
 sg13g2_and2_1 _10559_ (.A(net226),
    .B(_04305_),
    .X(_00987_));
 sg13g2_mux2_1 _10560_ (.A0(\shift_storage.storage[357] ),
    .A1(\shift_storage.storage[356] ),
    .S(net529),
    .X(_04306_));
 sg13g2_and2_1 _10561_ (.A(net228),
    .B(_04306_),
    .X(_00988_));
 sg13g2_mux2_1 _10562_ (.A0(\shift_storage.storage[358] ),
    .A1(\shift_storage.storage[357] ),
    .S(net529),
    .X(_04307_));
 sg13g2_and2_1 _10563_ (.A(net228),
    .B(_04307_),
    .X(_00989_));
 sg13g2_mux2_1 _10564_ (.A0(\shift_storage.storage[359] ),
    .A1(\shift_storage.storage[358] ),
    .S(net529),
    .X(_04308_));
 sg13g2_and2_1 _10565_ (.A(net228),
    .B(_04308_),
    .X(_00990_));
 sg13g2_mux2_1 _10566_ (.A0(\shift_storage.storage[35] ),
    .A1(\shift_storage.storage[34] ),
    .S(net626),
    .X(_04309_));
 sg13g2_and2_1 _10567_ (.A(net328),
    .B(_04309_),
    .X(_00991_));
 sg13g2_mux2_1 _10568_ (.A0(\shift_storage.storage[360] ),
    .A1(\shift_storage.storage[359] ),
    .S(net529),
    .X(_04310_));
 sg13g2_and2_1 _10569_ (.A(net228),
    .B(_04310_),
    .X(_00992_));
 sg13g2_buf_2 fanout170 (.A(\median_processor.input_storage[21] ),
    .X(net170));
 sg13g2_mux2_1 _10571_ (.A0(\shift_storage.storage[361] ),
    .A1(\shift_storage.storage[360] ),
    .S(net529),
    .X(_04312_));
 sg13g2_and2_1 _10572_ (.A(net228),
    .B(_04312_),
    .X(_00993_));
 sg13g2_mux2_1 _10573_ (.A0(\shift_storage.storage[362] ),
    .A1(\shift_storage.storage[361] ),
    .S(net537),
    .X(_04313_));
 sg13g2_and2_1 _10574_ (.A(net236),
    .B(_04313_),
    .X(_00994_));
 sg13g2_mux2_1 _10575_ (.A0(\shift_storage.storage[363] ),
    .A1(\shift_storage.storage[362] ),
    .S(net537),
    .X(_04314_));
 sg13g2_and2_1 _10576_ (.A(net236),
    .B(_04314_),
    .X(_00995_));
 sg13g2_buf_2 fanout169 (.A(net170),
    .X(net169));
 sg13g2_mux2_1 _10578_ (.A0(\shift_storage.storage[364] ),
    .A1(\shift_storage.storage[363] ),
    .S(net537),
    .X(_04316_));
 sg13g2_and2_1 _10579_ (.A(net236),
    .B(_04316_),
    .X(_00996_));
 sg13g2_mux2_1 _10580_ (.A0(\shift_storage.storage[365] ),
    .A1(\shift_storage.storage[364] ),
    .S(net529),
    .X(_04317_));
 sg13g2_and2_1 _10581_ (.A(net228),
    .B(_04317_),
    .X(_00997_));
 sg13g2_mux2_1 _10582_ (.A0(\shift_storage.storage[366] ),
    .A1(\shift_storage.storage[365] ),
    .S(net529),
    .X(_04318_));
 sg13g2_and2_1 _10583_ (.A(net228),
    .B(_04318_),
    .X(_00998_));
 sg13g2_mux2_1 _10584_ (.A0(\shift_storage.storage[367] ),
    .A1(\shift_storage.storage[366] ),
    .S(net530),
    .X(_04319_));
 sg13g2_and2_1 _10585_ (.A(net229),
    .B(_04319_),
    .X(_00999_));
 sg13g2_mux2_1 _10586_ (.A0(\shift_storage.storage[368] ),
    .A1(\shift_storage.storage[367] ),
    .S(net528),
    .X(_04320_));
 sg13g2_and2_1 _10587_ (.A(net229),
    .B(_04320_),
    .X(_01000_));
 sg13g2_mux2_1 _10588_ (.A0(\shift_storage.storage[369] ),
    .A1(\shift_storage.storage[368] ),
    .S(net528),
    .X(_04321_));
 sg13g2_and2_1 _10589_ (.A(net227),
    .B(_04321_),
    .X(_01001_));
 sg13g2_mux2_1 _10590_ (.A0(\shift_storage.storage[36] ),
    .A1(\shift_storage.storage[35] ),
    .S(net628),
    .X(_04322_));
 sg13g2_and2_1 _10591_ (.A(net330),
    .B(_04322_),
    .X(_01002_));
 sg13g2_buf_2 fanout168 (.A(\median_processor.input_storage[22] ),
    .X(net168));
 sg13g2_mux2_1 _10593_ (.A0(\shift_storage.storage[370] ),
    .A1(\shift_storage.storage[369] ),
    .S(net528),
    .X(_04324_));
 sg13g2_and2_1 _10594_ (.A(net227),
    .B(_04324_),
    .X(_01003_));
 sg13g2_mux2_1 _10595_ (.A0(\shift_storage.storage[371] ),
    .A1(\shift_storage.storage[370] ),
    .S(net528),
    .X(_04325_));
 sg13g2_and2_1 _10596_ (.A(net227),
    .B(_04325_),
    .X(_01004_));
 sg13g2_mux2_1 _10597_ (.A0(\shift_storage.storage[372] ),
    .A1(\shift_storage.storage[371] ),
    .S(net528),
    .X(_04326_));
 sg13g2_and2_1 _10598_ (.A(net227),
    .B(_04326_),
    .X(_01005_));
 sg13g2_buf_2 fanout167 (.A(\median_processor.input_storage[22] ),
    .X(net167));
 sg13g2_mux2_1 _10600_ (.A0(\shift_storage.storage[373] ),
    .A1(\shift_storage.storage[372] ),
    .S(net528),
    .X(_04328_));
 sg13g2_and2_1 _10601_ (.A(net227),
    .B(_04328_),
    .X(_01006_));
 sg13g2_mux2_1 _10602_ (.A0(\shift_storage.storage[374] ),
    .A1(\shift_storage.storage[373] ),
    .S(net528),
    .X(_04329_));
 sg13g2_and2_1 _10603_ (.A(net227),
    .B(_04329_),
    .X(_01007_));
 sg13g2_mux2_1 _10604_ (.A0(\shift_storage.storage[375] ),
    .A1(\shift_storage.storage[374] ),
    .S(net528),
    .X(_04330_));
 sg13g2_and2_1 _10605_ (.A(net227),
    .B(_04330_),
    .X(_01008_));
 sg13g2_mux2_1 _10606_ (.A0(\shift_storage.storage[376] ),
    .A1(\shift_storage.storage[375] ),
    .S(net530),
    .X(_04331_));
 sg13g2_and2_1 _10607_ (.A(net227),
    .B(_04331_),
    .X(_01009_));
 sg13g2_mux2_1 _10608_ (.A0(\shift_storage.storage[377] ),
    .A1(\shift_storage.storage[376] ),
    .S(net534),
    .X(_04332_));
 sg13g2_and2_1 _10609_ (.A(net233),
    .B(_04332_),
    .X(_01010_));
 sg13g2_mux2_1 _10610_ (.A0(\shift_storage.storage[378] ),
    .A1(\shift_storage.storage[377] ),
    .S(net540),
    .X(_04333_));
 sg13g2_and2_1 _10611_ (.A(net239),
    .B(_04333_),
    .X(_01011_));
 sg13g2_mux2_1 _10612_ (.A0(\shift_storage.storage[379] ),
    .A1(\shift_storage.storage[378] ),
    .S(net540),
    .X(_04334_));
 sg13g2_and2_1 _10613_ (.A(net239),
    .B(_04334_),
    .X(_01012_));
 sg13g2_buf_1 fanout166 (.A(\median_processor.input_storage[23] ),
    .X(net166));
 sg13g2_buf_2 fanout165 (.A(\median_processor.input_storage[23] ),
    .X(net165));
 sg13g2_mux2_1 _10616_ (.A0(\shift_storage.storage[37] ),
    .A1(\shift_storage.storage[36] ),
    .S(net628),
    .X(_04337_));
 sg13g2_and2_1 _10617_ (.A(net330),
    .B(_04337_),
    .X(_01013_));
 sg13g2_mux2_1 _10618_ (.A0(\shift_storage.storage[380] ),
    .A1(\shift_storage.storage[379] ),
    .S(net540),
    .X(_04338_));
 sg13g2_and2_1 _10619_ (.A(net239),
    .B(_04338_),
    .X(_01014_));
 sg13g2_mux2_1 _10620_ (.A0(\shift_storage.storage[381] ),
    .A1(\shift_storage.storage[380] ),
    .S(net540),
    .X(_04339_));
 sg13g2_and2_1 _10621_ (.A(net239),
    .B(_04339_),
    .X(_01015_));
 sg13g2_buf_1 fanout164 (.A(\median_processor.input_storage[24] ),
    .X(net164));
 sg13g2_buf_2 fanout163 (.A(\median_processor.input_storage[24] ),
    .X(net163));
 sg13g2_mux2_1 _10624_ (.A0(\shift_storage.storage[382] ),
    .A1(\shift_storage.storage[381] ),
    .S(net540),
    .X(_04342_));
 sg13g2_and2_1 _10625_ (.A(net241),
    .B(_04342_),
    .X(_01016_));
 sg13g2_mux2_1 _10626_ (.A0(\shift_storage.storage[383] ),
    .A1(\shift_storage.storage[382] ),
    .S(net543),
    .X(_04343_));
 sg13g2_and2_1 _10627_ (.A(net239),
    .B(_04343_),
    .X(_01017_));
 sg13g2_mux2_1 _10628_ (.A0(\shift_storage.storage[384] ),
    .A1(\shift_storage.storage[383] ),
    .S(net543),
    .X(_04344_));
 sg13g2_and2_1 _10629_ (.A(net239),
    .B(_04344_),
    .X(_01018_));
 sg13g2_mux2_1 _10630_ (.A0(\shift_storage.storage[385] ),
    .A1(\shift_storage.storage[384] ),
    .S(net543),
    .X(_04345_));
 sg13g2_and2_1 _10631_ (.A(net240),
    .B(_04345_),
    .X(_01019_));
 sg13g2_mux2_1 _10632_ (.A0(\shift_storage.storage[386] ),
    .A1(\shift_storage.storage[385] ),
    .S(net542),
    .X(_04346_));
 sg13g2_and2_1 _10633_ (.A(net242),
    .B(_04346_),
    .X(_01020_));
 sg13g2_mux2_1 _10634_ (.A0(\shift_storage.storage[387] ),
    .A1(\shift_storage.storage[386] ),
    .S(net542),
    .X(_04347_));
 sg13g2_and2_1 _10635_ (.A(net242),
    .B(_04347_),
    .X(_01021_));
 sg13g2_mux2_1 _10636_ (.A0(\shift_storage.storage[388] ),
    .A1(\shift_storage.storage[387] ),
    .S(net542),
    .X(_04348_));
 sg13g2_and2_1 _10637_ (.A(net242),
    .B(_04348_),
    .X(_01022_));
 sg13g2_buf_1 fanout162 (.A(\median_processor.input_storage[25] ),
    .X(net162));
 sg13g2_mux2_1 _10639_ (.A0(\shift_storage.storage[389] ),
    .A1(\shift_storage.storage[388] ),
    .S(net543),
    .X(_04350_));
 sg13g2_and2_1 _10640_ (.A(net243),
    .B(_04350_),
    .X(_01023_));
 sg13g2_mux2_1 _10641_ (.A0(\shift_storage.storage[38] ),
    .A1(\shift_storage.storage[37] ),
    .S(net627),
    .X(_04351_));
 sg13g2_and2_1 _10642_ (.A(net329),
    .B(_04351_),
    .X(_01024_));
 sg13g2_mux2_1 _10643_ (.A0(\shift_storage.storage[390] ),
    .A1(\shift_storage.storage[389] ),
    .S(net543),
    .X(_04352_));
 sg13g2_and2_1 _10644_ (.A(net243),
    .B(_04352_),
    .X(_01025_));
 sg13g2_buf_2 fanout161 (.A(\median_processor.input_storage[25] ),
    .X(net161));
 sg13g2_mux2_1 _10646_ (.A0(\shift_storage.storage[391] ),
    .A1(\shift_storage.storage[390] ),
    .S(net543),
    .X(_04354_));
 sg13g2_and2_1 _10647_ (.A(net243),
    .B(_04354_),
    .X(_01026_));
 sg13g2_mux2_1 _10648_ (.A0(\shift_storage.storage[392] ),
    .A1(\shift_storage.storage[391] ),
    .S(net543),
    .X(_04355_));
 sg13g2_and2_1 _10649_ (.A(net243),
    .B(_04355_),
    .X(_01027_));
 sg13g2_mux2_1 _10650_ (.A0(\shift_storage.storage[393] ),
    .A1(\shift_storage.storage[392] ),
    .S(net543),
    .X(_04356_));
 sg13g2_and2_1 _10651_ (.A(net243),
    .B(_04356_),
    .X(_01028_));
 sg13g2_mux2_1 _10652_ (.A0(\shift_storage.storage[394] ),
    .A1(\shift_storage.storage[393] ),
    .S(net572),
    .X(_04357_));
 sg13g2_and2_1 _10653_ (.A(net272),
    .B(_04357_),
    .X(_01029_));
 sg13g2_mux2_1 _10654_ (.A0(\shift_storage.storage[395] ),
    .A1(\shift_storage.storage[394] ),
    .S(net572),
    .X(_04358_));
 sg13g2_and2_1 _10655_ (.A(net272),
    .B(_04358_),
    .X(_01030_));
 sg13g2_mux2_1 _10656_ (.A0(\shift_storage.storage[396] ),
    .A1(\shift_storage.storage[395] ),
    .S(net572),
    .X(_04359_));
 sg13g2_and2_1 _10657_ (.A(net272),
    .B(_04359_),
    .X(_01031_));
 sg13g2_mux2_1 _10658_ (.A0(\shift_storage.storage[397] ),
    .A1(\shift_storage.storage[396] ),
    .S(net569),
    .X(_04360_));
 sg13g2_and2_1 _10659_ (.A(net269),
    .B(_04360_),
    .X(_01032_));
 sg13g2_buf_2 fanout160 (.A(\median_processor.input_storage[26] ),
    .X(net160));
 sg13g2_mux2_1 _10661_ (.A0(\shift_storage.storage[398] ),
    .A1(\shift_storage.storage[397] ),
    .S(net569),
    .X(_04362_));
 sg13g2_and2_1 _10662_ (.A(net269),
    .B(_04362_),
    .X(_01033_));
 sg13g2_mux2_1 _10663_ (.A0(\shift_storage.storage[399] ),
    .A1(\shift_storage.storage[398] ),
    .S(net569),
    .X(_04363_));
 sg13g2_and2_1 _10664_ (.A(net269),
    .B(_04363_),
    .X(_01034_));
 sg13g2_mux2_1 _10665_ (.A0(\shift_storage.storage[39] ),
    .A1(\shift_storage.storage[38] ),
    .S(net627),
    .X(_04364_));
 sg13g2_and2_1 _10666_ (.A(net329),
    .B(_04364_),
    .X(_01035_));
 sg13g2_buf_2 fanout159 (.A(\median_processor.input_storage[26] ),
    .X(net159));
 sg13g2_mux2_1 _10668_ (.A0(\shift_storage.storage[3] ),
    .A1(\shift_storage.storage[2] ),
    .S(net612),
    .X(_04366_));
 sg13g2_and2_1 _10669_ (.A(net314),
    .B(_04366_),
    .X(_01036_));
 sg13g2_mux2_1 _10670_ (.A0(\shift_storage.storage[400] ),
    .A1(\shift_storage.storage[399] ),
    .S(net568),
    .X(_04367_));
 sg13g2_and2_1 _10671_ (.A(net268),
    .B(_04367_),
    .X(_01037_));
 sg13g2_mux2_1 _10672_ (.A0(\shift_storage.storage[401] ),
    .A1(\shift_storage.storage[400] ),
    .S(net572),
    .X(_04368_));
 sg13g2_and2_1 _10673_ (.A(net272),
    .B(_04368_),
    .X(_01038_));
 sg13g2_mux2_1 _10674_ (.A0(\shift_storage.storage[402] ),
    .A1(\shift_storage.storage[401] ),
    .S(net575),
    .X(_04369_));
 sg13g2_and2_1 _10675_ (.A(net275),
    .B(_04369_),
    .X(_01039_));
 sg13g2_mux2_1 _10676_ (.A0(\shift_storage.storage[403] ),
    .A1(\shift_storage.storage[402] ),
    .S(net575),
    .X(_04370_));
 sg13g2_and2_1 _10677_ (.A(net275),
    .B(_04370_),
    .X(_01040_));
 sg13g2_mux2_1 _10678_ (.A0(\shift_storage.storage[404] ),
    .A1(\shift_storage.storage[403] ),
    .S(net575),
    .X(_04371_));
 sg13g2_and2_1 _10679_ (.A(net275),
    .B(_04371_),
    .X(_01041_));
 sg13g2_mux2_1 _10680_ (.A0(\shift_storage.storage[405] ),
    .A1(\shift_storage.storage[404] ),
    .S(net575),
    .X(_04372_));
 sg13g2_and2_1 _10681_ (.A(net275),
    .B(_04372_),
    .X(_01042_));
 sg13g2_buf_2 fanout158 (.A(\median_processor.input_storage[27] ),
    .X(net158));
 sg13g2_mux2_1 _10683_ (.A0(\shift_storage.storage[406] ),
    .A1(\shift_storage.storage[405] ),
    .S(net575),
    .X(_04374_));
 sg13g2_and2_1 _10684_ (.A(net275),
    .B(_04374_),
    .X(_01043_));
 sg13g2_mux2_1 _10685_ (.A0(\shift_storage.storage[407] ),
    .A1(\shift_storage.storage[406] ),
    .S(net582),
    .X(_04375_));
 sg13g2_and2_1 _10686_ (.A(net282),
    .B(_04375_),
    .X(_01044_));
 sg13g2_mux2_1 _10687_ (.A0(\shift_storage.storage[408] ),
    .A1(\shift_storage.storage[407] ),
    .S(net582),
    .X(_04376_));
 sg13g2_and2_1 _10688_ (.A(net282),
    .B(_04376_),
    .X(_01045_));
 sg13g2_buf_2 fanout157 (.A(net158),
    .X(net157));
 sg13g2_mux2_1 _10690_ (.A0(\shift_storage.storage[409] ),
    .A1(\shift_storage.storage[408] ),
    .S(net582),
    .X(_04378_));
 sg13g2_and2_1 _10691_ (.A(net282),
    .B(_04378_),
    .X(_01046_));
 sg13g2_mux2_1 _10692_ (.A0(\shift_storage.storage[40] ),
    .A1(\shift_storage.storage[39] ),
    .S(net627),
    .X(_04379_));
 sg13g2_and2_1 _10693_ (.A(net329),
    .B(_04379_),
    .X(_01047_));
 sg13g2_mux2_1 _10694_ (.A0(\shift_storage.storage[410] ),
    .A1(\shift_storage.storage[409] ),
    .S(net582),
    .X(_04380_));
 sg13g2_and2_1 _10695_ (.A(net282),
    .B(_04380_),
    .X(_01048_));
 sg13g2_mux2_1 _10696_ (.A0(\shift_storage.storage[411] ),
    .A1(\shift_storage.storage[410] ),
    .S(net583),
    .X(_04381_));
 sg13g2_and2_1 _10697_ (.A(net282),
    .B(_04381_),
    .X(_01049_));
 sg13g2_mux2_1 _10698_ (.A0(\shift_storage.storage[412] ),
    .A1(\shift_storage.storage[411] ),
    .S(net582),
    .X(_04382_));
 sg13g2_and2_1 _10699_ (.A(net283),
    .B(_04382_),
    .X(_01050_));
 sg13g2_mux2_1 _10700_ (.A0(\shift_storage.storage[413] ),
    .A1(\shift_storage.storage[412] ),
    .S(net582),
    .X(_04383_));
 sg13g2_and2_1 _10701_ (.A(net283),
    .B(_04383_),
    .X(_01051_));
 sg13g2_mux2_1 _10702_ (.A0(\shift_storage.storage[414] ),
    .A1(\shift_storage.storage[413] ),
    .S(net584),
    .X(_04384_));
 sg13g2_and2_1 _10703_ (.A(net284),
    .B(_04384_),
    .X(_01052_));
 sg13g2_buf_2 fanout156 (.A(\median_processor.input_storage[28] ),
    .X(net156));
 sg13g2_mux2_1 _10705_ (.A0(\shift_storage.storage[415] ),
    .A1(\shift_storage.storage[414] ),
    .S(net584),
    .X(_04386_));
 sg13g2_and2_1 _10706_ (.A(net284),
    .B(_04386_),
    .X(_01053_));
 sg13g2_mux2_1 _10707_ (.A0(\shift_storage.storage[416] ),
    .A1(\shift_storage.storage[415] ),
    .S(net584),
    .X(_04387_));
 sg13g2_and2_1 _10708_ (.A(net284),
    .B(_04387_),
    .X(_01054_));
 sg13g2_mux2_1 _10709_ (.A0(\shift_storage.storage[417] ),
    .A1(\shift_storage.storage[416] ),
    .S(net584),
    .X(_04388_));
 sg13g2_and2_1 _10710_ (.A(net284),
    .B(_04388_),
    .X(_01055_));
 sg13g2_buf_2 fanout155 (.A(net156),
    .X(net155));
 sg13g2_mux2_1 _10712_ (.A0(\shift_storage.storage[418] ),
    .A1(\shift_storage.storage[417] ),
    .S(net584),
    .X(_04390_));
 sg13g2_and2_1 _10713_ (.A(net284),
    .B(_04390_),
    .X(_01056_));
 sg13g2_mux2_1 _10714_ (.A0(\shift_storage.storage[419] ),
    .A1(\shift_storage.storage[418] ),
    .S(net584),
    .X(_04391_));
 sg13g2_and2_1 _10715_ (.A(net282),
    .B(_04391_),
    .X(_01057_));
 sg13g2_mux2_1 _10716_ (.A0(\shift_storage.storage[41] ),
    .A1(\shift_storage.storage[40] ),
    .S(net627),
    .X(_04392_));
 sg13g2_and2_1 _10717_ (.A(net329),
    .B(_04392_),
    .X(_01058_));
 sg13g2_mux2_1 _10718_ (.A0(\shift_storage.storage[420] ),
    .A1(\shift_storage.storage[419] ),
    .S(net577),
    .X(_04393_));
 sg13g2_and2_1 _10719_ (.A(net277),
    .B(_04393_),
    .X(_01059_));
 sg13g2_mux2_1 _10720_ (.A0(\shift_storage.storage[421] ),
    .A1(\shift_storage.storage[420] ),
    .S(net577),
    .X(_04394_));
 sg13g2_and2_1 _10721_ (.A(net277),
    .B(_04394_),
    .X(_01060_));
 sg13g2_mux2_1 _10722_ (.A0(\shift_storage.storage[422] ),
    .A1(\shift_storage.storage[421] ),
    .S(net577),
    .X(_04395_));
 sg13g2_and2_1 _10723_ (.A(net277),
    .B(_04395_),
    .X(_01061_));
 sg13g2_mux2_1 _10724_ (.A0(\shift_storage.storage[423] ),
    .A1(\shift_storage.storage[422] ),
    .S(net577),
    .X(_04396_));
 sg13g2_and2_1 _10725_ (.A(net277),
    .B(_04396_),
    .X(_01062_));
 sg13g2_buf_2 fanout154 (.A(\median_processor.input_storage[29] ),
    .X(net154));
 sg13g2_mux2_1 _10727_ (.A0(\shift_storage.storage[424] ),
    .A1(\shift_storage.storage[423] ),
    .S(net577),
    .X(_04398_));
 sg13g2_and2_1 _10728_ (.A(net277),
    .B(_04398_),
    .X(_01063_));
 sg13g2_mux2_1 _10729_ (.A0(\shift_storage.storage[425] ),
    .A1(\shift_storage.storage[424] ),
    .S(net577),
    .X(_04399_));
 sg13g2_and2_1 _10730_ (.A(net277),
    .B(_04399_),
    .X(_01064_));
 sg13g2_mux2_1 _10731_ (.A0(\shift_storage.storage[426] ),
    .A1(\shift_storage.storage[425] ),
    .S(net577),
    .X(_04400_));
 sg13g2_and2_1 _10732_ (.A(net277),
    .B(_04400_),
    .X(_01065_));
 sg13g2_buf_1 fanout153 (.A(net154),
    .X(net153));
 sg13g2_mux2_1 _10734_ (.A0(\shift_storage.storage[427] ),
    .A1(\shift_storage.storage[426] ),
    .S(net571),
    .X(_04402_));
 sg13g2_and2_1 _10735_ (.A(net271),
    .B(_04402_),
    .X(_01066_));
 sg13g2_mux2_1 _10736_ (.A0(\shift_storage.storage[428] ),
    .A1(\shift_storage.storage[427] ),
    .S(net571),
    .X(_04403_));
 sg13g2_and2_1 _10737_ (.A(net271),
    .B(_04403_),
    .X(_01067_));
 sg13g2_mux2_1 _10738_ (.A0(\shift_storage.storage[429] ),
    .A1(\shift_storage.storage[428] ),
    .S(net570),
    .X(_04404_));
 sg13g2_and2_1 _10739_ (.A(net270),
    .B(_04404_),
    .X(_01068_));
 sg13g2_mux2_1 _10740_ (.A0(\shift_storage.storage[42] ),
    .A1(\shift_storage.storage[41] ),
    .S(net627),
    .X(_04405_));
 sg13g2_and2_1 _10741_ (.A(net329),
    .B(_04405_),
    .X(_01069_));
 sg13g2_mux2_1 _10742_ (.A0(\shift_storage.storage[430] ),
    .A1(\shift_storage.storage[429] ),
    .S(net570),
    .X(_04406_));
 sg13g2_and2_1 _10743_ (.A(net270),
    .B(_04406_),
    .X(_01070_));
 sg13g2_mux2_1 _10744_ (.A0(\shift_storage.storage[431] ),
    .A1(\shift_storage.storage[430] ),
    .S(net570),
    .X(_04407_));
 sg13g2_and2_1 _10745_ (.A(net270),
    .B(_04407_),
    .X(_01071_));
 sg13g2_mux2_1 _10746_ (.A0(\shift_storage.storage[432] ),
    .A1(\shift_storage.storage[431] ),
    .S(net570),
    .X(_04408_));
 sg13g2_and2_1 _10747_ (.A(net270),
    .B(_04408_),
    .X(_01072_));
 sg13g2_buf_2 fanout152 (.A(net154),
    .X(net152));
 sg13g2_mux2_1 _10749_ (.A0(\shift_storage.storage[433] ),
    .A1(\shift_storage.storage[432] ),
    .S(net571),
    .X(_04410_));
 sg13g2_and2_1 _10750_ (.A(net271),
    .B(_04410_),
    .X(_01073_));
 sg13g2_mux2_1 _10751_ (.A0(\shift_storage.storage[434] ),
    .A1(\shift_storage.storage[433] ),
    .S(net569),
    .X(_04411_));
 sg13g2_and2_1 _10752_ (.A(net269),
    .B(_04411_),
    .X(_01074_));
 sg13g2_mux2_1 _10753_ (.A0(\shift_storage.storage[435] ),
    .A1(\shift_storage.storage[434] ),
    .S(net569),
    .X(_04412_));
 sg13g2_and2_1 _10754_ (.A(net268),
    .B(_04412_),
    .X(_01075_));
 sg13g2_buf_1 fanout151 (.A(\median_processor.input_storage[2] ),
    .X(net151));
 sg13g2_mux2_1 _10756_ (.A0(\shift_storage.storage[436] ),
    .A1(\shift_storage.storage[435] ),
    .S(net568),
    .X(_04414_));
 sg13g2_and2_1 _10757_ (.A(net269),
    .B(_04414_),
    .X(_01076_));
 sg13g2_mux2_1 _10758_ (.A0(\shift_storage.storage[437] ),
    .A1(\shift_storage.storage[436] ),
    .S(net569),
    .X(_04415_));
 sg13g2_and2_1 _10759_ (.A(net269),
    .B(_04415_),
    .X(_01077_));
 sg13g2_mux2_1 _10760_ (.A0(\shift_storage.storage[438] ),
    .A1(\shift_storage.storage[437] ),
    .S(net568),
    .X(_04416_));
 sg13g2_and2_1 _10761_ (.A(net268),
    .B(_04416_),
    .X(_01078_));
 sg13g2_mux2_1 _10762_ (.A0(\shift_storage.storage[439] ),
    .A1(\shift_storage.storage[438] ),
    .S(net538),
    .X(_04417_));
 sg13g2_and2_1 _10763_ (.A(net237),
    .B(_04417_),
    .X(_01079_));
 sg13g2_mux2_1 _10764_ (.A0(\shift_storage.storage[43] ),
    .A1(\shift_storage.storage[42] ),
    .S(net627),
    .X(_04418_));
 sg13g2_and2_1 _10765_ (.A(net329),
    .B(_04418_),
    .X(_01080_));
 sg13g2_mux2_1 _10766_ (.A0(\shift_storage.storage[440] ),
    .A1(\shift_storage.storage[439] ),
    .S(net538),
    .X(_04419_));
 sg13g2_and2_1 _10767_ (.A(net237),
    .B(_04419_),
    .X(_01081_));
 sg13g2_mux2_1 _10768_ (.A0(\shift_storage.storage[441] ),
    .A1(\shift_storage.storage[440] ),
    .S(net538),
    .X(_04420_));
 sg13g2_and2_1 _10769_ (.A(net237),
    .B(_04420_),
    .X(_01082_));
 sg13g2_buf_2 fanout150 (.A(net151),
    .X(net150));
 sg13g2_buf_2 fanout149 (.A(\median_processor.input_storage[30] ),
    .X(net149));
 sg13g2_mux2_1 _10772_ (.A0(\shift_storage.storage[442] ),
    .A1(\shift_storage.storage[441] ),
    .S(net538),
    .X(_04423_));
 sg13g2_and2_1 _10773_ (.A(net237),
    .B(_04423_),
    .X(_01083_));
 sg13g2_mux2_1 _10774_ (.A0(\shift_storage.storage[443] ),
    .A1(\shift_storage.storage[442] ),
    .S(net539),
    .X(_04424_));
 sg13g2_and2_1 _10775_ (.A(net238),
    .B(_04424_),
    .X(_01084_));
 sg13g2_mux2_1 _10776_ (.A0(\shift_storage.storage[444] ),
    .A1(\shift_storage.storage[443] ),
    .S(net539),
    .X(_04425_));
 sg13g2_and2_1 _10777_ (.A(net238),
    .B(_04425_),
    .X(_01085_));
 sg13g2_buf_2 fanout148 (.A(net149),
    .X(net148));
 sg13g2_buf_2 fanout147 (.A(\median_processor.input_storage[31] ),
    .X(net147));
 sg13g2_mux2_1 _10780_ (.A0(\shift_storage.storage[445] ),
    .A1(\shift_storage.storage[444] ),
    .S(net539),
    .X(_04428_));
 sg13g2_and2_1 _10781_ (.A(net235),
    .B(_04428_),
    .X(_01086_));
 sg13g2_mux2_1 _10782_ (.A0(\shift_storage.storage[446] ),
    .A1(\shift_storage.storage[445] ),
    .S(net536),
    .X(_04429_));
 sg13g2_and2_1 _10783_ (.A(net235),
    .B(_04429_),
    .X(_01087_));
 sg13g2_mux2_1 _10784_ (.A0(\shift_storage.storage[447] ),
    .A1(\shift_storage.storage[446] ),
    .S(net536),
    .X(_04430_));
 sg13g2_and2_1 _10785_ (.A(net235),
    .B(_04430_),
    .X(_01088_));
 sg13g2_mux2_1 _10786_ (.A0(\shift_storage.storage[448] ),
    .A1(\shift_storage.storage[447] ),
    .S(net536),
    .X(_04431_));
 sg13g2_and2_1 _10787_ (.A(net235),
    .B(_04431_),
    .X(_01089_));
 sg13g2_mux2_1 _10788_ (.A0(\shift_storage.storage[449] ),
    .A1(\shift_storage.storage[448] ),
    .S(net536),
    .X(_04432_));
 sg13g2_and2_1 _10789_ (.A(net235),
    .B(_04432_),
    .X(_01090_));
 sg13g2_mux2_1 _10790_ (.A0(\shift_storage.storage[44] ),
    .A1(\shift_storage.storage[43] ),
    .S(net621),
    .X(_04433_));
 sg13g2_and2_1 _10791_ (.A(net324),
    .B(_04433_),
    .X(_01091_));
 sg13g2_mux2_1 _10792_ (.A0(\shift_storage.storage[450] ),
    .A1(\shift_storage.storage[449] ),
    .S(net536),
    .X(_04434_));
 sg13g2_and2_1 _10793_ (.A(net235),
    .B(_04434_),
    .X(_01092_));
 sg13g2_buf_2 fanout146 (.A(\median_processor.input_storage[31] ),
    .X(net146));
 sg13g2_mux2_1 _10795_ (.A0(\shift_storage.storage[451] ),
    .A1(\shift_storage.storage[450] ),
    .S(net536),
    .X(_04436_));
 sg13g2_and2_1 _10796_ (.A(net235),
    .B(_04436_),
    .X(_01093_));
 sg13g2_mux2_1 _10797_ (.A0(\shift_storage.storage[452] ),
    .A1(\shift_storage.storage[451] ),
    .S(net536),
    .X(_04437_));
 sg13g2_and2_1 _10798_ (.A(net235),
    .B(_04437_),
    .X(_01094_));
 sg13g2_mux2_1 _10799_ (.A0(\shift_storage.storage[453] ),
    .A1(\shift_storage.storage[452] ),
    .S(net537),
    .X(_04438_));
 sg13g2_and2_1 _10800_ (.A(net236),
    .B(_04438_),
    .X(_01095_));
 sg13g2_buf_2 fanout145 (.A(\median_processor.input_storage[32] ),
    .X(net145));
 sg13g2_mux2_1 _10802_ (.A0(\shift_storage.storage[454] ),
    .A1(\shift_storage.storage[453] ),
    .S(net536),
    .X(_04440_));
 sg13g2_and2_1 _10803_ (.A(net236),
    .B(_04440_),
    .X(_01096_));
 sg13g2_mux2_1 _10804_ (.A0(\shift_storage.storage[455] ),
    .A1(\shift_storage.storage[454] ),
    .S(net537),
    .X(_04441_));
 sg13g2_and2_1 _10805_ (.A(net236),
    .B(_04441_),
    .X(_01097_));
 sg13g2_mux2_1 _10806_ (.A0(\shift_storage.storage[456] ),
    .A1(\shift_storage.storage[455] ),
    .S(net537),
    .X(_04442_));
 sg13g2_and2_1 _10807_ (.A(net236),
    .B(_04442_),
    .X(_01098_));
 sg13g2_mux2_1 _10808_ (.A0(\shift_storage.storage[457] ),
    .A1(\shift_storage.storage[456] ),
    .S(net538),
    .X(_04443_));
 sg13g2_and2_1 _10809_ (.A(net237),
    .B(_04443_),
    .X(_01099_));
 sg13g2_mux2_1 _10810_ (.A0(\shift_storage.storage[458] ),
    .A1(\shift_storage.storage[457] ),
    .S(net538),
    .X(_04444_));
 sg13g2_and2_1 _10811_ (.A(net237),
    .B(_04444_),
    .X(_01100_));
 sg13g2_mux2_1 _10812_ (.A0(\shift_storage.storage[459] ),
    .A1(\shift_storage.storage[458] ),
    .S(net538),
    .X(_04445_));
 sg13g2_and2_1 _10813_ (.A(net237),
    .B(_04445_),
    .X(_01101_));
 sg13g2_mux2_1 _10814_ (.A0(\shift_storage.storage[45] ),
    .A1(\shift_storage.storage[44] ),
    .S(net621),
    .X(_04446_));
 sg13g2_and2_1 _10815_ (.A(net324),
    .B(_04446_),
    .X(_01102_));
 sg13g2_buf_2 fanout144 (.A(net145),
    .X(net144));
 sg13g2_mux2_1 _10817_ (.A0(\shift_storage.storage[460] ),
    .A1(\shift_storage.storage[459] ),
    .S(net539),
    .X(_04448_));
 sg13g2_and2_1 _10818_ (.A(net238),
    .B(_04448_),
    .X(_01103_));
 sg13g2_mux2_1 _10819_ (.A0(\shift_storage.storage[461] ),
    .A1(\shift_storage.storage[460] ),
    .S(net538),
    .X(_04449_));
 sg13g2_and2_1 _10820_ (.A(net237),
    .B(_04449_),
    .X(_01104_));
 sg13g2_mux2_1 _10821_ (.A0(\shift_storage.storage[462] ),
    .A1(\shift_storage.storage[461] ),
    .S(net568),
    .X(_04450_));
 sg13g2_and2_1 _10822_ (.A(net268),
    .B(_04450_),
    .X(_01105_));
 sg13g2_buf_2 fanout143 (.A(\median_processor.input_storage[33] ),
    .X(net143));
 sg13g2_mux2_1 _10824_ (.A0(\shift_storage.storage[463] ),
    .A1(\shift_storage.storage[462] ),
    .S(net568),
    .X(_04452_));
 sg13g2_and2_1 _10825_ (.A(net268),
    .B(_04452_),
    .X(_01106_));
 sg13g2_mux2_1 _10826_ (.A0(\shift_storage.storage[464] ),
    .A1(\shift_storage.storage[463] ),
    .S(net568),
    .X(_04453_));
 sg13g2_and2_1 _10827_ (.A(net268),
    .B(_04453_),
    .X(_01107_));
 sg13g2_mux2_1 _10828_ (.A0(\shift_storage.storage[465] ),
    .A1(\shift_storage.storage[464] ),
    .S(net568),
    .X(_04454_));
 sg13g2_and2_1 _10829_ (.A(net268),
    .B(_04454_),
    .X(_01108_));
 sg13g2_mux2_1 _10830_ (.A0(\shift_storage.storage[466] ),
    .A1(\shift_storage.storage[465] ),
    .S(net568),
    .X(_04455_));
 sg13g2_and2_1 _10831_ (.A(net268),
    .B(_04455_),
    .X(_01109_));
 sg13g2_mux2_1 _10832_ (.A0(\shift_storage.storage[467] ),
    .A1(\shift_storage.storage[466] ),
    .S(net570),
    .X(_04456_));
 sg13g2_and2_1 _10833_ (.A(net270),
    .B(_04456_),
    .X(_01110_));
 sg13g2_mux2_1 _10834_ (.A0(\shift_storage.storage[468] ),
    .A1(\shift_storage.storage[467] ),
    .S(net570),
    .X(_04457_));
 sg13g2_and2_1 _10835_ (.A(net270),
    .B(_04457_),
    .X(_01111_));
 sg13g2_mux2_1 _10836_ (.A0(\shift_storage.storage[469] ),
    .A1(\shift_storage.storage[468] ),
    .S(net570),
    .X(_04458_));
 sg13g2_and2_1 _10837_ (.A(net270),
    .B(_04458_),
    .X(_01112_));
 sg13g2_buf_2 fanout142 (.A(\median_processor.input_storage[33] ),
    .X(net142));
 sg13g2_mux2_1 _10839_ (.A0(\shift_storage.storage[46] ),
    .A1(\shift_storage.storage[45] ),
    .S(net621),
    .X(_04460_));
 sg13g2_and2_1 _10840_ (.A(net322),
    .B(_04460_),
    .X(_01113_));
 sg13g2_mux2_1 _10841_ (.A0(\shift_storage.storage[470] ),
    .A1(\shift_storage.storage[469] ),
    .S(net570),
    .X(_04461_));
 sg13g2_and2_1 _10842_ (.A(net270),
    .B(_04461_),
    .X(_01114_));
 sg13g2_mux2_1 _10843_ (.A0(\shift_storage.storage[471] ),
    .A1(\shift_storage.storage[470] ),
    .S(net554),
    .X(_04462_));
 sg13g2_and2_1 _10844_ (.A(net254),
    .B(_04462_),
    .X(_01115_));
 sg13g2_buf_2 fanout141 (.A(\median_processor.input_storage[34] ),
    .X(net141));
 sg13g2_mux2_1 _10846_ (.A0(\shift_storage.storage[472] ),
    .A1(\shift_storage.storage[471] ),
    .S(net563),
    .X(_04464_));
 sg13g2_and2_1 _10847_ (.A(net263),
    .B(_04464_),
    .X(_01116_));
 sg13g2_mux2_1 _10848_ (.A0(\shift_storage.storage[473] ),
    .A1(\shift_storage.storage[472] ),
    .S(net578),
    .X(_04465_));
 sg13g2_and2_1 _10849_ (.A(net278),
    .B(_04465_),
    .X(_01117_));
 sg13g2_mux2_1 _10850_ (.A0(\shift_storage.storage[474] ),
    .A1(\shift_storage.storage[473] ),
    .S(net578),
    .X(_04466_));
 sg13g2_and2_1 _10851_ (.A(net278),
    .B(_04466_),
    .X(_01118_));
 sg13g2_mux2_1 _10852_ (.A0(\shift_storage.storage[475] ),
    .A1(\shift_storage.storage[474] ),
    .S(net578),
    .X(_04467_));
 sg13g2_and2_1 _10853_ (.A(net278),
    .B(_04467_),
    .X(_01119_));
 sg13g2_mux2_1 _10854_ (.A0(\shift_storage.storage[476] ),
    .A1(\shift_storage.storage[475] ),
    .S(net578),
    .X(_04468_));
 sg13g2_and2_1 _10855_ (.A(net278),
    .B(_04468_),
    .X(_01120_));
 sg13g2_mux2_1 _10856_ (.A0(\shift_storage.storage[477] ),
    .A1(\shift_storage.storage[476] ),
    .S(net578),
    .X(_04469_));
 sg13g2_and2_1 _10857_ (.A(net278),
    .B(_04469_),
    .X(_01121_));
 sg13g2_mux2_1 _10858_ (.A0(\shift_storage.storage[478] ),
    .A1(\shift_storage.storage[477] ),
    .S(net581),
    .X(_04470_));
 sg13g2_and2_1 _10859_ (.A(net281),
    .B(_04470_),
    .X(_01122_));
 sg13g2_buf_2 fanout140 (.A(net141),
    .X(net140));
 sg13g2_mux2_1 _10861_ (.A0(\shift_storage.storage[479] ),
    .A1(\shift_storage.storage[478] ),
    .S(net581),
    .X(_04472_));
 sg13g2_and2_1 _10862_ (.A(net277),
    .B(_04472_),
    .X(_01123_));
 sg13g2_mux2_1 _10863_ (.A0(\shift_storage.storage[47] ),
    .A1(\shift_storage.storage[46] ),
    .S(net621),
    .X(_04473_));
 sg13g2_and2_1 _10864_ (.A(net324),
    .B(_04473_),
    .X(_01124_));
 sg13g2_mux2_1 _10865_ (.A0(\shift_storage.storage[480] ),
    .A1(\shift_storage.storage[479] ),
    .S(net577),
    .X(_04474_));
 sg13g2_and2_1 _10866_ (.A(net281),
    .B(_04474_),
    .X(_01125_));
 sg13g2_buf_2 fanout139 (.A(\median_processor.input_storage[35] ),
    .X(net139));
 sg13g2_mux2_1 _10868_ (.A0(\shift_storage.storage[481] ),
    .A1(\shift_storage.storage[480] ),
    .S(net579),
    .X(_04476_));
 sg13g2_and2_1 _10869_ (.A(net279),
    .B(_04476_),
    .X(_01126_));
 sg13g2_mux2_1 _10870_ (.A0(\shift_storage.storage[482] ),
    .A1(\shift_storage.storage[481] ),
    .S(net579),
    .X(_04477_));
 sg13g2_and2_1 _10871_ (.A(net279),
    .B(_04477_),
    .X(_01127_));
 sg13g2_mux2_1 _10872_ (.A0(\shift_storage.storage[483] ),
    .A1(\shift_storage.storage[482] ),
    .S(net579),
    .X(_04478_));
 sg13g2_and2_1 _10873_ (.A(net279),
    .B(_04478_),
    .X(_01128_));
 sg13g2_mux2_1 _10874_ (.A0(\shift_storage.storage[484] ),
    .A1(\shift_storage.storage[483] ),
    .S(net579),
    .X(_04479_));
 sg13g2_and2_1 _10875_ (.A(net279),
    .B(_04479_),
    .X(_01129_));
 sg13g2_mux2_1 _10876_ (.A0(\shift_storage.storage[485] ),
    .A1(\shift_storage.storage[484] ),
    .S(net581),
    .X(_04480_));
 sg13g2_and2_1 _10877_ (.A(net281),
    .B(_04480_),
    .X(_01130_));
 sg13g2_mux2_1 _10878_ (.A0(\shift_storage.storage[486] ),
    .A1(\shift_storage.storage[485] ),
    .S(net579),
    .X(_04481_));
 sg13g2_and2_1 _10879_ (.A(net279),
    .B(_04481_),
    .X(_01131_));
 sg13g2_mux2_1 _10880_ (.A0(\shift_storage.storage[487] ),
    .A1(\shift_storage.storage[486] ),
    .S(net579),
    .X(_04482_));
 sg13g2_and2_1 _10881_ (.A(net279),
    .B(_04482_),
    .X(_01132_));
 sg13g2_buf_2 fanout138 (.A(net139),
    .X(net138));
 sg13g2_mux2_1 _10883_ (.A0(\shift_storage.storage[488] ),
    .A1(\shift_storage.storage[487] ),
    .S(net579),
    .X(_04484_));
 sg13g2_and2_1 _10884_ (.A(net279),
    .B(_04484_),
    .X(_01133_));
 sg13g2_mux2_1 _10885_ (.A0(\shift_storage.storage[489] ),
    .A1(\shift_storage.storage[488] ),
    .S(net579),
    .X(_04485_));
 sg13g2_and2_1 _10886_ (.A(net279),
    .B(_04485_),
    .X(_01134_));
 sg13g2_mux2_1 _10887_ (.A0(\shift_storage.storage[48] ),
    .A1(\shift_storage.storage[47] ),
    .S(net621),
    .X(_04486_));
 sg13g2_and2_1 _10888_ (.A(net324),
    .B(_04486_),
    .X(_01135_));
 sg13g2_buf_2 fanout137 (.A(\median_processor.input_storage[36] ),
    .X(net137));
 sg13g2_mux2_1 _10890_ (.A0(\shift_storage.storage[490] ),
    .A1(\shift_storage.storage[489] ),
    .S(net580),
    .X(_04488_));
 sg13g2_and2_1 _10891_ (.A(net280),
    .B(_04488_),
    .X(_01136_));
 sg13g2_mux2_1 _10892_ (.A0(\shift_storage.storage[491] ),
    .A1(\shift_storage.storage[490] ),
    .S(net580),
    .X(_04489_));
 sg13g2_and2_1 _10893_ (.A(net280),
    .B(_04489_),
    .X(_01137_));
 sg13g2_mux2_1 _10894_ (.A0(\shift_storage.storage[492] ),
    .A1(\shift_storage.storage[491] ),
    .S(net580),
    .X(_04490_));
 sg13g2_and2_1 _10895_ (.A(net280),
    .B(_04490_),
    .X(_01138_));
 sg13g2_mux2_1 _10896_ (.A0(\shift_storage.storage[493] ),
    .A1(\shift_storage.storage[492] ),
    .S(net580),
    .X(_04491_));
 sg13g2_and2_1 _10897_ (.A(net280),
    .B(_04491_),
    .X(_01139_));
 sg13g2_mux2_1 _10898_ (.A0(\shift_storage.storage[494] ),
    .A1(\shift_storage.storage[493] ),
    .S(net580),
    .X(_04492_));
 sg13g2_and2_1 _10899_ (.A(net280),
    .B(_04492_),
    .X(_01140_));
 sg13g2_mux2_1 _10900_ (.A0(\shift_storage.storage[495] ),
    .A1(\shift_storage.storage[494] ),
    .S(net580),
    .X(_04493_));
 sg13g2_and2_1 _10901_ (.A(net280),
    .B(_04493_),
    .X(_01141_));
 sg13g2_mux2_1 _10902_ (.A0(\shift_storage.storage[496] ),
    .A1(\shift_storage.storage[495] ),
    .S(net580),
    .X(_04494_));
 sg13g2_and2_1 _10903_ (.A(net280),
    .B(_04494_),
    .X(_01142_));
 sg13g2_buf_2 fanout136 (.A(\median_processor.input_storage[36] ),
    .X(net136));
 sg13g2_mux2_1 _10905_ (.A0(\shift_storage.storage[497] ),
    .A1(\shift_storage.storage[496] ),
    .S(net578),
    .X(_04496_));
 sg13g2_and2_1 _10906_ (.A(net278),
    .B(_04496_),
    .X(_01143_));
 sg13g2_mux2_1 _10907_ (.A0(\shift_storage.storage[498] ),
    .A1(\shift_storage.storage[497] ),
    .S(net578),
    .X(_04497_));
 sg13g2_and2_1 _10908_ (.A(net278),
    .B(_04497_),
    .X(_01144_));
 sg13g2_mux2_1 _10909_ (.A0(\shift_storage.storage[499] ),
    .A1(\shift_storage.storage[498] ),
    .S(net578),
    .X(_04498_));
 sg13g2_and2_1 _10910_ (.A(net278),
    .B(_04498_),
    .X(_01145_));
 sg13g2_buf_2 fanout135 (.A(\median_processor.input_storage[37] ),
    .X(net135));
 sg13g2_mux2_1 _10912_ (.A0(\shift_storage.storage[49] ),
    .A1(\shift_storage.storage[48] ),
    .S(net621),
    .X(_04500_));
 sg13g2_and2_1 _10913_ (.A(net324),
    .B(_04500_),
    .X(_01146_));
 sg13g2_mux2_1 _10914_ (.A0(\shift_storage.storage[4] ),
    .A1(\shift_storage.storage[3] ),
    .S(net612),
    .X(_04501_));
 sg13g2_and2_1 _10915_ (.A(net314),
    .B(_04501_),
    .X(_01147_));
 sg13g2_mux2_1 _10916_ (.A0(\shift_storage.storage[500] ),
    .A1(\shift_storage.storage[499] ),
    .S(net563),
    .X(_04502_));
 sg13g2_and2_1 _10917_ (.A(net263),
    .B(_04502_),
    .X(_01148_));
 sg13g2_mux2_1 _10918_ (.A0(\shift_storage.storage[501] ),
    .A1(\shift_storage.storage[500] ),
    .S(net566),
    .X(_04503_));
 sg13g2_and2_1 _10919_ (.A(net263),
    .B(_04503_),
    .X(_01149_));
 sg13g2_mux2_1 _10920_ (.A0(\shift_storage.storage[502] ),
    .A1(\shift_storage.storage[501] ),
    .S(net563),
    .X(_04504_));
 sg13g2_and2_1 _10921_ (.A(net263),
    .B(_04504_),
    .X(_01150_));
 sg13g2_mux2_1 _10922_ (.A0(\shift_storage.storage[503] ),
    .A1(\shift_storage.storage[502] ),
    .S(net563),
    .X(_04505_));
 sg13g2_and2_1 _10923_ (.A(net263),
    .B(_04505_),
    .X(_01151_));
 sg13g2_mux2_1 _10924_ (.A0(\shift_storage.storage[504] ),
    .A1(\shift_storage.storage[503] ),
    .S(net563),
    .X(_04506_));
 sg13g2_and2_1 _10925_ (.A(net263),
    .B(_04506_),
    .X(_01152_));
 sg13g2_buf_2 fanout134 (.A(\median_processor.input_storage[37] ),
    .X(net134));
 sg13g2_buf_1 fanout133 (.A(\median_processor.input_storage[38] ),
    .X(net133));
 sg13g2_buf_2 fanout132 (.A(\median_processor.input_storage[38] ),
    .X(net132));
 sg13g2_mux2_1 _10929_ (.A0(\shift_storage.storage[505] ),
    .A1(\shift_storage.storage[504] ),
    .S(net563),
    .X(_04510_));
 sg13g2_and2_1 _10930_ (.A(net266),
    .B(_04510_),
    .X(_01153_));
 sg13g2_mux2_1 _10931_ (.A0(\shift_storage.storage[506] ),
    .A1(\shift_storage.storage[505] ),
    .S(net566),
    .X(_04511_));
 sg13g2_and2_1 _10932_ (.A(net254),
    .B(_04511_),
    .X(_01154_));
 sg13g2_mux2_1 _10933_ (.A0(\shift_storage.storage[507] ),
    .A1(\shift_storage.storage[506] ),
    .S(net554),
    .X(_04512_));
 sg13g2_and2_1 _10934_ (.A(net254),
    .B(_04512_),
    .X(_01155_));
 sg13g2_buf_2 fanout131 (.A(\median_processor.input_storage[39] ),
    .X(net131));
 sg13g2_buf_2 fanout130 (.A(\median_processor.input_storage[39] ),
    .X(net130));
 sg13g2_buf_1 fanout129 (.A(\median_processor.input_storage[3] ),
    .X(net129));
 sg13g2_mux2_1 _10938_ (.A0(\shift_storage.storage[508] ),
    .A1(\shift_storage.storage[507] ),
    .S(net554),
    .X(_04516_));
 sg13g2_and2_1 _10939_ (.A(net254),
    .B(_04516_),
    .X(_01156_));
 sg13g2_mux2_1 _10940_ (.A0(\shift_storage.storage[509] ),
    .A1(\shift_storage.storage[508] ),
    .S(net554),
    .X(_04517_));
 sg13g2_and2_1 _10941_ (.A(net254),
    .B(_04517_),
    .X(_01157_));
 sg13g2_mux2_1 _10942_ (.A0(\shift_storage.storage[50] ),
    .A1(\shift_storage.storage[49] ),
    .S(net622),
    .X(_04518_));
 sg13g2_and2_1 _10943_ (.A(net323),
    .B(_04518_),
    .X(_01158_));
 sg13g2_mux2_1 _10944_ (.A0(\shift_storage.storage[510] ),
    .A1(\shift_storage.storage[509] ),
    .S(net554),
    .X(_04519_));
 sg13g2_and2_1 _10945_ (.A(net254),
    .B(_04519_),
    .X(_01159_));
 sg13g2_mux2_1 _10946_ (.A0(\shift_storage.storage[511] ),
    .A1(\shift_storage.storage[510] ),
    .S(net554),
    .X(_04520_));
 sg13g2_and2_1 _10947_ (.A(net254),
    .B(_04520_),
    .X(_01160_));
 sg13g2_mux2_1 _10948_ (.A0(\shift_storage.storage[512] ),
    .A1(\shift_storage.storage[511] ),
    .S(net555),
    .X(_04521_));
 sg13g2_and2_1 _10949_ (.A(net254),
    .B(_04521_),
    .X(_01161_));
 sg13g2_mux2_1 _10950_ (.A0(\shift_storage.storage[513] ),
    .A1(\shift_storage.storage[512] ),
    .S(net555),
    .X(_04522_));
 sg13g2_and2_1 _10951_ (.A(net252),
    .B(_04522_),
    .X(_01162_));
 sg13g2_buf_2 fanout128 (.A(net129),
    .X(net128));
 sg13g2_mux2_1 _10953_ (.A0(\shift_storage.storage[514] ),
    .A1(\shift_storage.storage[513] ),
    .S(net555),
    .X(_04524_));
 sg13g2_and2_1 _10954_ (.A(net252),
    .B(_04524_),
    .X(_01163_));
 sg13g2_mux2_1 _10955_ (.A0(\shift_storage.storage[515] ),
    .A1(\shift_storage.storage[514] ),
    .S(net555),
    .X(_04525_));
 sg13g2_and2_1 _10956_ (.A(net252),
    .B(_04525_),
    .X(_01164_));
 sg13g2_mux2_1 _10957_ (.A0(\shift_storage.storage[516] ),
    .A1(\shift_storage.storage[515] ),
    .S(net555),
    .X(_04526_));
 sg13g2_and2_1 _10958_ (.A(net252),
    .B(_04526_),
    .X(_01165_));
 sg13g2_buf_2 fanout127 (.A(\median_processor.input_storage[40] ),
    .X(net127));
 sg13g2_mux2_1 _10960_ (.A0(\shift_storage.storage[517] ),
    .A1(\shift_storage.storage[516] ),
    .S(net552),
    .X(_04528_));
 sg13g2_and2_1 _10961_ (.A(net252),
    .B(_04528_),
    .X(_01166_));
 sg13g2_mux2_1 _10962_ (.A0(\shift_storage.storage[518] ),
    .A1(\shift_storage.storage[517] ),
    .S(net552),
    .X(_04529_));
 sg13g2_and2_1 _10963_ (.A(net224),
    .B(_04529_),
    .X(_01167_));
 sg13g2_mux2_1 _10964_ (.A0(\shift_storage.storage[519] ),
    .A1(\shift_storage.storage[518] ),
    .S(net525),
    .X(_04530_));
 sg13g2_and2_1 _10965_ (.A(net224),
    .B(_04530_),
    .X(_01168_));
 sg13g2_mux2_1 _10966_ (.A0(\shift_storage.storage[51] ),
    .A1(\shift_storage.storage[50] ),
    .S(net622),
    .X(_04531_));
 sg13g2_and2_1 _10967_ (.A(net323),
    .B(_04531_),
    .X(_01169_));
 sg13g2_mux2_1 _10968_ (.A0(\shift_storage.storage[520] ),
    .A1(\shift_storage.storage[519] ),
    .S(net525),
    .X(_04532_));
 sg13g2_and2_1 _10969_ (.A(net224),
    .B(_04532_),
    .X(_01170_));
 sg13g2_mux2_1 _10970_ (.A0(\shift_storage.storage[521] ),
    .A1(\shift_storage.storage[520] ),
    .S(net525),
    .X(_04533_));
 sg13g2_and2_1 _10971_ (.A(net224),
    .B(_04533_),
    .X(_01171_));
 sg13g2_mux2_1 _10972_ (.A0(\shift_storage.storage[522] ),
    .A1(\shift_storage.storage[521] ),
    .S(net525),
    .X(_04534_));
 sg13g2_and2_1 _10973_ (.A(net224),
    .B(_04534_),
    .X(_01172_));
 sg13g2_buf_1 fanout126 (.A(\median_processor.input_storage[42] ),
    .X(net126));
 sg13g2_mux2_1 _10975_ (.A0(\shift_storage.storage[523] ),
    .A1(\shift_storage.storage[522] ),
    .S(net525),
    .X(_04536_));
 sg13g2_and2_1 _10976_ (.A(net224),
    .B(_04536_),
    .X(_01173_));
 sg13g2_mux2_1 _10977_ (.A0(\shift_storage.storage[524] ),
    .A1(\shift_storage.storage[523] ),
    .S(net523),
    .X(_04537_));
 sg13g2_and2_1 _10978_ (.A(net222),
    .B(_04537_),
    .X(_01174_));
 sg13g2_mux2_1 _10979_ (.A0(\shift_storage.storage[525] ),
    .A1(\shift_storage.storage[524] ),
    .S(net523),
    .X(_04538_));
 sg13g2_and2_1 _10980_ (.A(net222),
    .B(_04538_),
    .X(_01175_));
 sg13g2_buf_2 fanout125 (.A(\median_processor.input_storage[42] ),
    .X(net125));
 sg13g2_mux2_1 _10982_ (.A0(\shift_storage.storage[526] ),
    .A1(\shift_storage.storage[525] ),
    .S(net523),
    .X(_04540_));
 sg13g2_and2_1 _10983_ (.A(net222),
    .B(_04540_),
    .X(_01176_));
 sg13g2_mux2_1 _10984_ (.A0(\shift_storage.storage[527] ),
    .A1(\shift_storage.storage[526] ),
    .S(net523),
    .X(_04541_));
 sg13g2_and2_1 _10985_ (.A(net221),
    .B(_04541_),
    .X(_01177_));
 sg13g2_mux2_1 _10986_ (.A0(\shift_storage.storage[528] ),
    .A1(\shift_storage.storage[527] ),
    .S(net523),
    .X(_04542_));
 sg13g2_and2_1 _10987_ (.A(net221),
    .B(_04542_),
    .X(_01178_));
 sg13g2_mux2_1 _10988_ (.A0(\shift_storage.storage[529] ),
    .A1(\shift_storage.storage[528] ),
    .S(net523),
    .X(_04543_));
 sg13g2_and2_1 _10989_ (.A(net222),
    .B(_04543_),
    .X(_01179_));
 sg13g2_mux2_1 _10990_ (.A0(\shift_storage.storage[52] ),
    .A1(\shift_storage.storage[51] ),
    .S(net622),
    .X(_04544_));
 sg13g2_and2_1 _10991_ (.A(net323),
    .B(_04544_),
    .X(_01180_));
 sg13g2_mux2_1 _10992_ (.A0(\shift_storage.storage[530] ),
    .A1(\shift_storage.storage[529] ),
    .S(net523),
    .X(_04545_));
 sg13g2_and2_1 _10993_ (.A(net222),
    .B(_04545_),
    .X(_01181_));
 sg13g2_mux2_1 _10994_ (.A0(\shift_storage.storage[531] ),
    .A1(\shift_storage.storage[530] ),
    .S(net522),
    .X(_04546_));
 sg13g2_and2_1 _10995_ (.A(net222),
    .B(_04546_),
    .X(_01182_));
 sg13g2_buf_1 fanout124 (.A(\median_processor.input_storage[43] ),
    .X(net124));
 sg13g2_mux2_1 _10997_ (.A0(\shift_storage.storage[532] ),
    .A1(\shift_storage.storage[531] ),
    .S(net515),
    .X(_04548_));
 sg13g2_and2_1 _10998_ (.A(net214),
    .B(_04548_),
    .X(_01183_));
 sg13g2_mux2_1 _10999_ (.A0(\shift_storage.storage[533] ),
    .A1(\shift_storage.storage[532] ),
    .S(net515),
    .X(_04549_));
 sg13g2_and2_1 _11000_ (.A(net214),
    .B(_04549_),
    .X(_01184_));
 sg13g2_mux2_1 _11001_ (.A0(\shift_storage.storage[534] ),
    .A1(\shift_storage.storage[533] ),
    .S(net515),
    .X(_04550_));
 sg13g2_and2_1 _11002_ (.A(net213),
    .B(_04550_),
    .X(_01185_));
 sg13g2_buf_2 fanout123 (.A(net124),
    .X(net123));
 sg13g2_mux2_1 _11004_ (.A0(\shift_storage.storage[535] ),
    .A1(\shift_storage.storage[534] ),
    .S(net515),
    .X(_04552_));
 sg13g2_and2_1 _11005_ (.A(net213),
    .B(_04552_),
    .X(_01186_));
 sg13g2_mux2_1 _11006_ (.A0(\shift_storage.storage[536] ),
    .A1(\shift_storage.storage[535] ),
    .S(net514),
    .X(_04553_));
 sg13g2_and2_1 _11007_ (.A(net213),
    .B(_04553_),
    .X(_01187_));
 sg13g2_mux2_1 _11008_ (.A0(\shift_storage.storage[537] ),
    .A1(\shift_storage.storage[536] ),
    .S(net514),
    .X(_04554_));
 sg13g2_and2_1 _11009_ (.A(net212),
    .B(_04554_),
    .X(_01188_));
 sg13g2_mux2_1 _11010_ (.A0(\shift_storage.storage[538] ),
    .A1(\shift_storage.storage[537] ),
    .S(net516),
    .X(_04555_));
 sg13g2_and2_1 _11011_ (.A(net211),
    .B(_04555_),
    .X(_01189_));
 sg13g2_mux2_1 _11012_ (.A0(\shift_storage.storage[539] ),
    .A1(\shift_storage.storage[538] ),
    .S(net516),
    .X(_04556_));
 sg13g2_and2_1 _11013_ (.A(net212),
    .B(_04556_),
    .X(_01190_));
 sg13g2_mux2_1 _11014_ (.A0(\shift_storage.storage[53] ),
    .A1(\shift_storage.storage[52] ),
    .S(net630),
    .X(_04557_));
 sg13g2_and2_1 _11015_ (.A(net323),
    .B(_04557_),
    .X(_01191_));
 sg13g2_mux2_1 _11016_ (.A0(\shift_storage.storage[540] ),
    .A1(\shift_storage.storage[539] ),
    .S(net513),
    .X(_04558_));
 sg13g2_and2_1 _11017_ (.A(net212),
    .B(_04558_),
    .X(_01192_));
 sg13g2_buf_1 fanout122 (.A(\median_processor.input_storage[44] ),
    .X(net122));
 sg13g2_mux2_1 _11019_ (.A0(\shift_storage.storage[541] ),
    .A1(\shift_storage.storage[540] ),
    .S(net516),
    .X(_04560_));
 sg13g2_and2_1 _11020_ (.A(net212),
    .B(_04560_),
    .X(_01193_));
 sg13g2_mux2_1 _11021_ (.A0(\shift_storage.storage[542] ),
    .A1(\shift_storage.storage[541] ),
    .S(net513),
    .X(_04561_));
 sg13g2_and2_1 _11022_ (.A(net211),
    .B(_04561_),
    .X(_01194_));
 sg13g2_mux2_1 _11023_ (.A0(\shift_storage.storage[543] ),
    .A1(\shift_storage.storage[542] ),
    .S(net513),
    .X(_04562_));
 sg13g2_and2_1 _11024_ (.A(net211),
    .B(_04562_),
    .X(_01195_));
 sg13g2_buf_1 fanout121 (.A(net122),
    .X(net121));
 sg13g2_mux2_1 _11026_ (.A0(\shift_storage.storage[544] ),
    .A1(\shift_storage.storage[543] ),
    .S(net513),
    .X(_04564_));
 sg13g2_and2_1 _11027_ (.A(net211),
    .B(_04564_),
    .X(_01196_));
 sg13g2_mux2_1 _11028_ (.A0(\shift_storage.storage[545] ),
    .A1(\shift_storage.storage[544] ),
    .S(net513),
    .X(_04565_));
 sg13g2_and2_1 _11029_ (.A(net211),
    .B(_04565_),
    .X(_01197_));
 sg13g2_mux2_1 _11030_ (.A0(\shift_storage.storage[546] ),
    .A1(\shift_storage.storage[545] ),
    .S(net513),
    .X(_04566_));
 sg13g2_and2_1 _11031_ (.A(net211),
    .B(_04566_),
    .X(_01198_));
 sg13g2_mux2_1 _11032_ (.A0(\shift_storage.storage[547] ),
    .A1(\shift_storage.storage[546] ),
    .S(net513),
    .X(_04567_));
 sg13g2_and2_1 _11033_ (.A(net211),
    .B(_04567_),
    .X(_01199_));
 sg13g2_mux2_1 _11034_ (.A0(\shift_storage.storage[548] ),
    .A1(\shift_storage.storage[547] ),
    .S(net513),
    .X(_04568_));
 sg13g2_and2_1 _11035_ (.A(net211),
    .B(_04568_),
    .X(_01200_));
 sg13g2_mux2_1 _11036_ (.A0(\shift_storage.storage[549] ),
    .A1(\shift_storage.storage[548] ),
    .S(net508),
    .X(_04569_));
 sg13g2_and2_1 _11037_ (.A(net206),
    .B(_04569_),
    .X(_01201_));
 sg13g2_mux2_1 _11038_ (.A0(\shift_storage.storage[54] ),
    .A1(\shift_storage.storage[53] ),
    .S(net630),
    .X(_04570_));
 sg13g2_and2_1 _11039_ (.A(net332),
    .B(_04570_),
    .X(_01202_));
 sg13g2_buf_2 fanout120 (.A(net121),
    .X(net120));
 sg13g2_mux2_1 _11041_ (.A0(\shift_storage.storage[550] ),
    .A1(\shift_storage.storage[549] ),
    .S(net509),
    .X(_04572_));
 sg13g2_and2_1 _11042_ (.A(net206),
    .B(_04572_),
    .X(_01203_));
 sg13g2_mux2_1 _11043_ (.A0(\shift_storage.storage[551] ),
    .A1(\shift_storage.storage[550] ),
    .S(net512),
    .X(_04573_));
 sg13g2_and2_1 _11044_ (.A(net210),
    .B(_04573_),
    .X(_01204_));
 sg13g2_mux2_1 _11045_ (.A0(\shift_storage.storage[552] ),
    .A1(\shift_storage.storage[551] ),
    .S(net512),
    .X(_04574_));
 sg13g2_and2_1 _11046_ (.A(net210),
    .B(_04574_),
    .X(_01205_));
 sg13g2_buf_1 fanout119 (.A(\median_processor.input_storage[45] ),
    .X(net119));
 sg13g2_mux2_1 _11048_ (.A0(\shift_storage.storage[553] ),
    .A1(\shift_storage.storage[552] ),
    .S(net514),
    .X(_04576_));
 sg13g2_and2_1 _11049_ (.A(net213),
    .B(_04576_),
    .X(_01206_));
 sg13g2_mux2_1 _11050_ (.A0(\shift_storage.storage[554] ),
    .A1(\shift_storage.storage[553] ),
    .S(net514),
    .X(_04577_));
 sg13g2_and2_1 _11051_ (.A(net213),
    .B(_04577_),
    .X(_01207_));
 sg13g2_mux2_1 _11052_ (.A0(\shift_storage.storage[555] ),
    .A1(\shift_storage.storage[554] ),
    .S(net514),
    .X(_04578_));
 sg13g2_and2_1 _11053_ (.A(net213),
    .B(_04578_),
    .X(_01208_));
 sg13g2_mux2_1 _11054_ (.A0(\shift_storage.storage[556] ),
    .A1(\shift_storage.storage[555] ),
    .S(net514),
    .X(_04579_));
 sg13g2_and2_1 _11055_ (.A(net213),
    .B(_04579_),
    .X(_01209_));
 sg13g2_mux2_1 _11056_ (.A0(\shift_storage.storage[557] ),
    .A1(\shift_storage.storage[556] ),
    .S(net514),
    .X(_04580_));
 sg13g2_and2_1 _11057_ (.A(net214),
    .B(_04580_),
    .X(_01210_));
 sg13g2_mux2_1 _11058_ (.A0(\shift_storage.storage[558] ),
    .A1(\shift_storage.storage[557] ),
    .S(net515),
    .X(_04581_));
 sg13g2_and2_1 _11059_ (.A(net214),
    .B(_04581_),
    .X(_01211_));
 sg13g2_mux2_1 _11060_ (.A0(\shift_storage.storage[559] ),
    .A1(\shift_storage.storage[558] ),
    .S(net514),
    .X(_04582_));
 sg13g2_and2_1 _11061_ (.A(net214),
    .B(_04582_),
    .X(_01212_));
 sg13g2_buf_2 fanout118 (.A(\median_processor.input_storage[45] ),
    .X(net118));
 sg13g2_mux2_1 _11063_ (.A0(\shift_storage.storage[55] ),
    .A1(\shift_storage.storage[54] ),
    .S(net630),
    .X(_04584_));
 sg13g2_and2_1 _11064_ (.A(net332),
    .B(_04584_),
    .X(_01213_));
 sg13g2_mux2_1 _11065_ (.A0(\shift_storage.storage[560] ),
    .A1(\shift_storage.storage[559] ),
    .S(net522),
    .X(_04585_));
 sg13g2_and2_1 _11066_ (.A(net213),
    .B(_04585_),
    .X(_01214_));
 sg13g2_mux2_1 _11067_ (.A0(\shift_storage.storage[561] ),
    .A1(\shift_storage.storage[560] ),
    .S(net522),
    .X(_04586_));
 sg13g2_and2_1 _11068_ (.A(net221),
    .B(_04586_),
    .X(_01215_));
 sg13g2_buf_2 fanout117 (.A(\median_processor.input_storage[46] ),
    .X(net117));
 sg13g2_mux2_1 _11070_ (.A0(\shift_storage.storage[562] ),
    .A1(\shift_storage.storage[561] ),
    .S(net522),
    .X(_04588_));
 sg13g2_and2_1 _11071_ (.A(net221),
    .B(_04588_),
    .X(_01216_));
 sg13g2_mux2_1 _11072_ (.A0(\shift_storage.storage[563] ),
    .A1(\shift_storage.storage[562] ),
    .S(net522),
    .X(_04589_));
 sg13g2_and2_1 _11073_ (.A(net221),
    .B(_04589_),
    .X(_01217_));
 sg13g2_mux2_1 _11074_ (.A0(\shift_storage.storage[564] ),
    .A1(\shift_storage.storage[563] ),
    .S(net522),
    .X(_04590_));
 sg13g2_and2_1 _11075_ (.A(net221),
    .B(_04590_),
    .X(_01218_));
 sg13g2_mux2_1 _11076_ (.A0(\shift_storage.storage[565] ),
    .A1(\shift_storage.storage[564] ),
    .S(net522),
    .X(_04591_));
 sg13g2_and2_1 _11077_ (.A(net221),
    .B(_04591_),
    .X(_01219_));
 sg13g2_mux2_1 _11078_ (.A0(\shift_storage.storage[566] ),
    .A1(\shift_storage.storage[565] ),
    .S(net522),
    .X(_04592_));
 sg13g2_and2_1 _11079_ (.A(net221),
    .B(_04592_),
    .X(_01220_));
 sg13g2_mux2_1 _11080_ (.A0(\shift_storage.storage[567] ),
    .A1(\shift_storage.storage[566] ),
    .S(net521),
    .X(_04593_));
 sg13g2_and2_1 _11081_ (.A(net218),
    .B(_04593_),
    .X(_01221_));
 sg13g2_mux2_1 _11082_ (.A0(\shift_storage.storage[568] ),
    .A1(\shift_storage.storage[567] ),
    .S(net521),
    .X(_04594_));
 sg13g2_and2_1 _11083_ (.A(net217),
    .B(_04594_),
    .X(_01222_));
 sg13g2_buf_1 fanout116 (.A(\median_processor.input_storage[46] ),
    .X(net116));
 sg13g2_buf_1 fanout115 (.A(net116),
    .X(net115));
 sg13g2_mux2_1 _11086_ (.A0(\shift_storage.storage[569] ),
    .A1(\shift_storage.storage[568] ),
    .S(net518),
    .X(_04597_));
 sg13g2_and2_1 _11087_ (.A(net217),
    .B(_04597_),
    .X(_01223_));
 sg13g2_mux2_1 _11088_ (.A0(\shift_storage.storage[56] ),
    .A1(\shift_storage.storage[55] ),
    .S(net630),
    .X(_04598_));
 sg13g2_and2_1 _11089_ (.A(net332),
    .B(_04598_),
    .X(_01224_));
 sg13g2_mux2_1 _11090_ (.A0(\shift_storage.storage[570] ),
    .A1(\shift_storage.storage[569] ),
    .S(net518),
    .X(_04599_));
 sg13g2_and2_1 _11091_ (.A(net217),
    .B(_04599_),
    .X(_01225_));
 sg13g2_buf_2 fanout114 (.A(net115),
    .X(net114));
 sg13g2_buf_2 fanout113 (.A(\median_processor.input_storage[47] ),
    .X(net113));
 sg13g2_mux2_1 _11094_ (.A0(\shift_storage.storage[571] ),
    .A1(\shift_storage.storage[570] ),
    .S(net518),
    .X(_04602_));
 sg13g2_and2_1 _11095_ (.A(net217),
    .B(_04602_),
    .X(_01226_));
 sg13g2_mux2_1 _11096_ (.A0(\shift_storage.storage[572] ),
    .A1(\shift_storage.storage[571] ),
    .S(net518),
    .X(_04603_));
 sg13g2_and2_1 _11097_ (.A(net217),
    .B(_04603_),
    .X(_01227_));
 sg13g2_mux2_1 _11098_ (.A0(\shift_storage.storage[573] ),
    .A1(\shift_storage.storage[572] ),
    .S(net517),
    .X(_04604_));
 sg13g2_and2_1 _11099_ (.A(net216),
    .B(_04604_),
    .X(_01228_));
 sg13g2_mux2_1 _11100_ (.A0(\shift_storage.storage[574] ),
    .A1(\shift_storage.storage[573] ),
    .S(net517),
    .X(_04605_));
 sg13g2_and2_1 _11101_ (.A(net216),
    .B(_04605_),
    .X(_01229_));
 sg13g2_mux2_1 _11102_ (.A0(\shift_storage.storage[575] ),
    .A1(\shift_storage.storage[574] ),
    .S(net511),
    .X(_04606_));
 sg13g2_and2_1 _11103_ (.A(net209),
    .B(_04606_),
    .X(_01230_));
 sg13g2_mux2_1 _11104_ (.A0(\shift_storage.storage[576] ),
    .A1(\shift_storage.storage[575] ),
    .S(net510),
    .X(_04607_));
 sg13g2_and2_1 _11105_ (.A(net208),
    .B(_04607_),
    .X(_01231_));
 sg13g2_mux2_1 _11106_ (.A0(\shift_storage.storage[577] ),
    .A1(\shift_storage.storage[576] ),
    .S(net511),
    .X(_04608_));
 sg13g2_and2_1 _11107_ (.A(net208),
    .B(_04608_),
    .X(_01232_));
 sg13g2_buf_1 fanout112 (.A(\median_processor.input_storage[48] ),
    .X(net112));
 sg13g2_mux2_1 _11109_ (.A0(\shift_storage.storage[578] ),
    .A1(\shift_storage.storage[577] ),
    .S(net511),
    .X(_04610_));
 sg13g2_and2_1 _11110_ (.A(net209),
    .B(_04610_),
    .X(_01233_));
 sg13g2_mux2_1 _11111_ (.A0(\shift_storage.storage[579] ),
    .A1(\shift_storage.storage[578] ),
    .S(net511),
    .X(_04611_));
 sg13g2_and2_1 _11112_ (.A(net209),
    .B(_04611_),
    .X(_01234_));
 sg13g2_mux2_1 _11113_ (.A0(\shift_storage.storage[57] ),
    .A1(\shift_storage.storage[56] ),
    .S(net631),
    .X(_04612_));
 sg13g2_and2_1 _11114_ (.A(net333),
    .B(_04612_),
    .X(_01235_));
 sg13g2_buf_2 fanout111 (.A(\median_processor.input_storage[48] ),
    .X(net111));
 sg13g2_mux2_1 _11116_ (.A0(\shift_storage.storage[580] ),
    .A1(\shift_storage.storage[579] ),
    .S(net511),
    .X(_04614_));
 sg13g2_and2_1 _11117_ (.A(net209),
    .B(_04614_),
    .X(_01236_));
 sg13g2_mux2_1 _11118_ (.A0(\shift_storage.storage[581] ),
    .A1(\shift_storage.storage[580] ),
    .S(net511),
    .X(_04615_));
 sg13g2_and2_1 _11119_ (.A(net209),
    .B(_04615_),
    .X(_01237_));
 sg13g2_mux2_1 _11120_ (.A0(\shift_storage.storage[582] ),
    .A1(\shift_storage.storage[581] ),
    .S(net511),
    .X(_04616_));
 sg13g2_and2_1 _11121_ (.A(net209),
    .B(_04616_),
    .X(_01238_));
 sg13g2_mux2_1 _11122_ (.A0(\shift_storage.storage[583] ),
    .A1(\shift_storage.storage[582] ),
    .S(net508),
    .X(_04617_));
 sg13g2_and2_1 _11123_ (.A(net207),
    .B(_04617_),
    .X(_01239_));
 sg13g2_mux2_1 _11124_ (.A0(\shift_storage.storage[584] ),
    .A1(\shift_storage.storage[583] ),
    .S(net509),
    .X(_04618_));
 sg13g2_and2_1 _11125_ (.A(net207),
    .B(_04618_),
    .X(_01240_));
 sg13g2_mux2_1 _11126_ (.A0(\shift_storage.storage[585] ),
    .A1(\shift_storage.storage[584] ),
    .S(net508),
    .X(_04619_));
 sg13g2_and2_1 _11127_ (.A(net206),
    .B(_04619_),
    .X(_01241_));
 sg13g2_mux2_1 _11128_ (.A0(\shift_storage.storage[586] ),
    .A1(\shift_storage.storage[585] ),
    .S(net508),
    .X(_04620_));
 sg13g2_and2_1 _11129_ (.A(net206),
    .B(_04620_),
    .X(_01242_));
 sg13g2_buf_2 fanout110 (.A(\median_processor.input_storage[49] ),
    .X(net110));
 sg13g2_mux2_1 _11131_ (.A0(\shift_storage.storage[587] ),
    .A1(\shift_storage.storage[586] ),
    .S(net508),
    .X(_04622_));
 sg13g2_and2_1 _11132_ (.A(net206),
    .B(_04622_),
    .X(_01243_));
 sg13g2_mux2_1 _11133_ (.A0(\shift_storage.storage[588] ),
    .A1(\shift_storage.storage[587] ),
    .S(net508),
    .X(_04623_));
 sg13g2_and2_1 _11134_ (.A(net206),
    .B(_04623_),
    .X(_01244_));
 sg13g2_mux2_1 _11135_ (.A0(\shift_storage.storage[589] ),
    .A1(\shift_storage.storage[588] ),
    .S(net508),
    .X(_04624_));
 sg13g2_and2_1 _11136_ (.A(net206),
    .B(_04624_),
    .X(_01245_));
 sg13g2_buf_2 fanout109 (.A(\median_processor.input_storage[4] ),
    .X(net109));
 sg13g2_mux2_1 _11138_ (.A0(\shift_storage.storage[58] ),
    .A1(\shift_storage.storage[57] ),
    .S(net631),
    .X(_04626_));
 sg13g2_and2_1 _11139_ (.A(net333),
    .B(_04626_),
    .X(_01246_));
 sg13g2_mux2_1 _11140_ (.A0(\shift_storage.storage[590] ),
    .A1(\shift_storage.storage[589] ),
    .S(net508),
    .X(_04627_));
 sg13g2_and2_1 _11141_ (.A(net206),
    .B(_04627_),
    .X(_01247_));
 sg13g2_mux2_1 _11142_ (.A0(\shift_storage.storage[591] ),
    .A1(\shift_storage.storage[590] ),
    .S(net506),
    .X(_04628_));
 sg13g2_and2_1 _11143_ (.A(net204),
    .B(_04628_),
    .X(_01248_));
 sg13g2_mux2_1 _11144_ (.A0(\shift_storage.storage[592] ),
    .A1(\shift_storage.storage[591] ),
    .S(net506),
    .X(_04629_));
 sg13g2_and2_1 _11145_ (.A(net204),
    .B(_04629_),
    .X(_01249_));
 sg13g2_mux2_1 _11146_ (.A0(\shift_storage.storage[593] ),
    .A1(\shift_storage.storage[592] ),
    .S(net506),
    .X(_04630_));
 sg13g2_and2_1 _11147_ (.A(net204),
    .B(_04630_),
    .X(_01250_));
 sg13g2_mux2_1 _11148_ (.A0(\shift_storage.storage[594] ),
    .A1(\shift_storage.storage[593] ),
    .S(net506),
    .X(_04631_));
 sg13g2_and2_1 _11149_ (.A(net204),
    .B(_04631_),
    .X(_01251_));
 sg13g2_mux2_1 _11150_ (.A0(\shift_storage.storage[595] ),
    .A1(\shift_storage.storage[594] ),
    .S(net506),
    .X(_04632_));
 sg13g2_and2_1 _11151_ (.A(net204),
    .B(_04632_),
    .X(_01252_));
 sg13g2_buf_2 fanout108 (.A(\median_processor.input_storage[50] ),
    .X(net108));
 sg13g2_mux2_1 _11153_ (.A0(\shift_storage.storage[596] ),
    .A1(\shift_storage.storage[595] ),
    .S(net506),
    .X(_04634_));
 sg13g2_and2_1 _11154_ (.A(net204),
    .B(_04634_),
    .X(_01253_));
 sg13g2_mux2_1 _11155_ (.A0(\shift_storage.storage[597] ),
    .A1(\shift_storage.storage[596] ),
    .S(net507),
    .X(_04635_));
 sg13g2_and2_1 _11156_ (.A(net205),
    .B(_04635_),
    .X(_01254_));
 sg13g2_mux2_1 _11157_ (.A0(\shift_storage.storage[598] ),
    .A1(\shift_storage.storage[597] ),
    .S(net507),
    .X(_04636_));
 sg13g2_and2_1 _11158_ (.A(net204),
    .B(_04636_),
    .X(_01255_));
 sg13g2_buf_2 fanout107 (.A(\median_processor.input_storage[50] ),
    .X(net107));
 sg13g2_mux2_1 _11160_ (.A0(\shift_storage.storage[599] ),
    .A1(\shift_storage.storage[598] ),
    .S(net506),
    .X(_04638_));
 sg13g2_and2_1 _11161_ (.A(net205),
    .B(_04638_),
    .X(_01256_));
 sg13g2_mux2_1 _11162_ (.A0(\shift_storage.storage[59] ),
    .A1(\shift_storage.storage[58] ),
    .S(net631),
    .X(_04639_));
 sg13g2_and2_1 _11163_ (.A(net333),
    .B(_04639_),
    .X(_01257_));
 sg13g2_mux2_1 _11164_ (.A0(\shift_storage.storage[5] ),
    .A1(\shift_storage.storage[4] ),
    .S(net612),
    .X(_04640_));
 sg13g2_and2_1 _11165_ (.A(net314),
    .B(_04640_),
    .X(_01258_));
 sg13g2_mux2_1 _11166_ (.A0(\shift_storage.storage[600] ),
    .A1(\shift_storage.storage[599] ),
    .S(net507),
    .X(_04641_));
 sg13g2_and2_1 _11167_ (.A(net205),
    .B(_04641_),
    .X(_01259_));
 sg13g2_mux2_1 _11168_ (.A0(\shift_storage.storage[601] ),
    .A1(\shift_storage.storage[600] ),
    .S(net507),
    .X(_04642_));
 sg13g2_and2_1 _11169_ (.A(net205),
    .B(_04642_),
    .X(_01260_));
 sg13g2_mux2_1 _11170_ (.A0(\shift_storage.storage[602] ),
    .A1(\shift_storage.storage[601] ),
    .S(net506),
    .X(_04643_));
 sg13g2_and2_1 _11171_ (.A(net204),
    .B(_04643_),
    .X(_01261_));
 sg13g2_mux2_1 _11172_ (.A0(\shift_storage.storage[603] ),
    .A1(\shift_storage.storage[602] ),
    .S(net510),
    .X(_04644_));
 sg13g2_and2_1 _11173_ (.A(net208),
    .B(_04644_),
    .X(_01262_));
 sg13g2_buf_2 fanout106 (.A(\median_processor.input_storage[51] ),
    .X(net106));
 sg13g2_mux2_1 _11175_ (.A0(\shift_storage.storage[604] ),
    .A1(\shift_storage.storage[603] ),
    .S(net510),
    .X(_04646_));
 sg13g2_and2_1 _11176_ (.A(net208),
    .B(_04646_),
    .X(_01263_));
 sg13g2_mux2_1 _11177_ (.A0(\shift_storage.storage[605] ),
    .A1(\shift_storage.storage[604] ),
    .S(net510),
    .X(_04647_));
 sg13g2_and2_1 _11178_ (.A(net208),
    .B(_04647_),
    .X(_01264_));
 sg13g2_mux2_1 _11179_ (.A0(\shift_storage.storage[606] ),
    .A1(\shift_storage.storage[605] ),
    .S(net510),
    .X(_04648_));
 sg13g2_and2_1 _11180_ (.A(net208),
    .B(_04648_),
    .X(_01265_));
 sg13g2_buf_2 fanout105 (.A(net106),
    .X(net105));
 sg13g2_mux2_1 _11182_ (.A0(\shift_storage.storage[607] ),
    .A1(\shift_storage.storage[606] ),
    .S(net510),
    .X(_04650_));
 sg13g2_and2_1 _11183_ (.A(net208),
    .B(_04650_),
    .X(_01266_));
 sg13g2_mux2_1 _11184_ (.A0(\shift_storage.storage[608] ),
    .A1(\shift_storage.storage[607] ),
    .S(net510),
    .X(_04651_));
 sg13g2_and2_1 _11185_ (.A(net209),
    .B(_04651_),
    .X(_01267_));
 sg13g2_mux2_1 _11186_ (.A0(\shift_storage.storage[609] ),
    .A1(\shift_storage.storage[608] ),
    .S(net510),
    .X(_04652_));
 sg13g2_and2_1 _11187_ (.A(net208),
    .B(_04652_),
    .X(_01268_));
 sg13g2_mux2_1 _11188_ (.A0(\shift_storage.storage[60] ),
    .A1(\shift_storage.storage[59] ),
    .S(net631),
    .X(_04653_));
 sg13g2_and2_1 _11189_ (.A(net333),
    .B(_04653_),
    .X(_01269_));
 sg13g2_mux2_1 _11190_ (.A0(\shift_storage.storage[610] ),
    .A1(\shift_storage.storage[609] ),
    .S(net517),
    .X(_04654_));
 sg13g2_and2_1 _11191_ (.A(net216),
    .B(_04654_),
    .X(_01270_));
 sg13g2_mux2_1 _11192_ (.A0(\shift_storage.storage[611] ),
    .A1(\shift_storage.storage[610] ),
    .S(net517),
    .X(_04655_));
 sg13g2_and2_1 _11193_ (.A(net216),
    .B(_04655_),
    .X(_01271_));
 sg13g2_mux2_1 _11194_ (.A0(\shift_storage.storage[612] ),
    .A1(\shift_storage.storage[611] ),
    .S(net517),
    .X(_04656_));
 sg13g2_and2_1 _11195_ (.A(net216),
    .B(_04656_),
    .X(_01272_));
 sg13g2_buf_1 fanout104 (.A(\median_processor.input_storage[52] ),
    .X(net104));
 sg13g2_mux2_1 _11197_ (.A0(\shift_storage.storage[613] ),
    .A1(\shift_storage.storage[612] ),
    .S(net517),
    .X(_04658_));
 sg13g2_and2_1 _11198_ (.A(net216),
    .B(_04658_),
    .X(_01273_));
 sg13g2_mux2_1 _11199_ (.A0(\shift_storage.storage[614] ),
    .A1(\shift_storage.storage[613] ),
    .S(net518),
    .X(_04659_));
 sg13g2_and2_1 _11200_ (.A(net218),
    .B(_04659_),
    .X(_01274_));
 sg13g2_mux2_1 _11201_ (.A0(\shift_storage.storage[615] ),
    .A1(\shift_storage.storage[614] ),
    .S(net518),
    .X(_04660_));
 sg13g2_and2_1 _11202_ (.A(net218),
    .B(_04660_),
    .X(_01275_));
 sg13g2_buf_2 fanout103 (.A(\median_processor.input_storage[52] ),
    .X(net103));
 sg13g2_mux2_1 _11204_ (.A0(\shift_storage.storage[616] ),
    .A1(\shift_storage.storage[615] ),
    .S(net519),
    .X(_04662_));
 sg13g2_and2_1 _11205_ (.A(net219),
    .B(_04662_),
    .X(_01276_));
 sg13g2_mux2_1 _11206_ (.A0(\shift_storage.storage[617] ),
    .A1(\shift_storage.storage[616] ),
    .S(net519),
    .X(_04663_));
 sg13g2_and2_1 _11207_ (.A(net219),
    .B(_04663_),
    .X(_01277_));
 sg13g2_mux2_1 _11208_ (.A0(\shift_storage.storage[618] ),
    .A1(\shift_storage.storage[617] ),
    .S(net519),
    .X(_04664_));
 sg13g2_and2_1 _11209_ (.A(net219),
    .B(_04664_),
    .X(_01278_));
 sg13g2_mux2_1 _11210_ (.A0(\shift_storage.storage[619] ),
    .A1(\shift_storage.storage[618] ),
    .S(net519),
    .X(_04665_));
 sg13g2_and2_1 _11211_ (.A(net219),
    .B(_04665_),
    .X(_01279_));
 sg13g2_mux2_1 _11212_ (.A0(\shift_storage.storage[61] ),
    .A1(\shift_storage.storage[60] ),
    .S(net631),
    .X(_04666_));
 sg13g2_and2_1 _11213_ (.A(net333),
    .B(_04666_),
    .X(_01280_));
 sg13g2_mux2_1 _11214_ (.A0(\shift_storage.storage[620] ),
    .A1(\shift_storage.storage[619] ),
    .S(net517),
    .X(_04667_));
 sg13g2_and2_1 _11215_ (.A(net216),
    .B(_04667_),
    .X(_01281_));
 sg13g2_mux2_1 _11216_ (.A0(\shift_storage.storage[621] ),
    .A1(\shift_storage.storage[620] ),
    .S(net517),
    .X(_04668_));
 sg13g2_and2_1 _11217_ (.A(net216),
    .B(_04668_),
    .X(_01282_));
 sg13g2_buf_2 fanout102 (.A(\median_processor.input_storage[53] ),
    .X(net102));
 sg13g2_mux2_1 _11219_ (.A0(\shift_storage.storage[622] ),
    .A1(\shift_storage.storage[621] ),
    .S(net518),
    .X(_04670_));
 sg13g2_and2_1 _11220_ (.A(net217),
    .B(_04670_),
    .X(_01283_));
 sg13g2_mux2_1 _11221_ (.A0(\shift_storage.storage[623] ),
    .A1(\shift_storage.storage[622] ),
    .S(net521),
    .X(_04671_));
 sg13g2_and2_1 _11222_ (.A(net217),
    .B(_04671_),
    .X(_01284_));
 sg13g2_mux2_1 _11223_ (.A0(\shift_storage.storage[624] ),
    .A1(\shift_storage.storage[623] ),
    .S(net520),
    .X(_04672_));
 sg13g2_and2_1 _11224_ (.A(net217),
    .B(_04672_),
    .X(_01285_));
 sg13g2_buf_2 fanout101 (.A(\median_processor.input_storage[53] ),
    .X(net101));
 sg13g2_mux2_1 _11226_ (.A0(\shift_storage.storage[625] ),
    .A1(\shift_storage.storage[624] ),
    .S(net521),
    .X(_04674_));
 sg13g2_and2_1 _11227_ (.A(net220),
    .B(_04674_),
    .X(_01286_));
 sg13g2_mux2_1 _11228_ (.A0(\shift_storage.storage[626] ),
    .A1(\shift_storage.storage[625] ),
    .S(net521),
    .X(_04675_));
 sg13g2_and2_1 _11229_ (.A(net220),
    .B(_04675_),
    .X(_01287_));
 sg13g2_mux2_1 _11230_ (.A0(\shift_storage.storage[627] ),
    .A1(\shift_storage.storage[626] ),
    .S(net520),
    .X(_04676_));
 sg13g2_and2_1 _11231_ (.A(net225),
    .B(_04676_),
    .X(_01288_));
 sg13g2_mux2_1 _11232_ (.A0(\shift_storage.storage[628] ),
    .A1(\shift_storage.storage[627] ),
    .S(net520),
    .X(_04677_));
 sg13g2_and2_1 _11233_ (.A(net220),
    .B(_04677_),
    .X(_01289_));
 sg13g2_mux2_1 _11234_ (.A0(\shift_storage.storage[629] ),
    .A1(\shift_storage.storage[628] ),
    .S(net548),
    .X(_04678_));
 sg13g2_and2_1 _11235_ (.A(net247),
    .B(_04678_),
    .X(_01290_));
 sg13g2_mux2_1 _11236_ (.A0(\shift_storage.storage[62] ),
    .A1(\shift_storage.storage[61] ),
    .S(net621),
    .X(_04679_));
 sg13g2_and2_1 _11237_ (.A(net324),
    .B(_04679_),
    .X(_01291_));
 sg13g2_mux2_1 _11238_ (.A0(\shift_storage.storage[630] ),
    .A1(\shift_storage.storage[629] ),
    .S(net548),
    .X(_04680_));
 sg13g2_and2_1 _11239_ (.A(net247),
    .B(_04680_),
    .X(_01292_));
 sg13g2_buf_1 fanout100 (.A(\median_processor.input_storage[54] ),
    .X(net100));
 sg13g2_buf_2 fanout99 (.A(\median_processor.input_storage[54] ),
    .X(net99));
 sg13g2_mux2_1 _11242_ (.A0(\shift_storage.storage[631] ),
    .A1(\shift_storage.storage[630] ),
    .S(net552),
    .X(_04683_));
 sg13g2_and2_1 _11243_ (.A(net251),
    .B(_04683_),
    .X(_01293_));
 sg13g2_mux2_1 _11244_ (.A0(\shift_storage.storage[632] ),
    .A1(\shift_storage.storage[631] ),
    .S(net525),
    .X(_04684_));
 sg13g2_and2_1 _11245_ (.A(net224),
    .B(_04684_),
    .X(_01294_));
 sg13g2_mux2_1 _11246_ (.A0(\shift_storage.storage[633] ),
    .A1(\shift_storage.storage[632] ),
    .S(net524),
    .X(_04685_));
 sg13g2_and2_1 _11247_ (.A(net223),
    .B(_04685_),
    .X(_01295_));
 sg13g2_buf_1 fanout98 (.A(\median_processor.input_storage[55] ),
    .X(net98));
 sg13g2_buf_2 fanout97 (.A(\median_processor.input_storage[55] ),
    .X(net97));
 sg13g2_mux2_1 _11250_ (.A0(\shift_storage.storage[634] ),
    .A1(\shift_storage.storage[633] ),
    .S(net524),
    .X(_04688_));
 sg13g2_and2_1 _11251_ (.A(net223),
    .B(_04688_),
    .X(_01296_));
 sg13g2_mux2_1 _11252_ (.A0(\shift_storage.storage[635] ),
    .A1(\shift_storage.storage[634] ),
    .S(net524),
    .X(_04689_));
 sg13g2_and2_1 _11253_ (.A(net223),
    .B(_04689_),
    .X(_01297_));
 sg13g2_mux2_1 _11254_ (.A0(\shift_storage.storage[636] ),
    .A1(\shift_storage.storage[635] ),
    .S(net524),
    .X(_04690_));
 sg13g2_and2_1 _11255_ (.A(net223),
    .B(_04690_),
    .X(_01298_));
 sg13g2_mux2_1 _11256_ (.A0(\shift_storage.storage[637] ),
    .A1(\shift_storage.storage[636] ),
    .S(net524),
    .X(_04691_));
 sg13g2_and2_1 _11257_ (.A(net223),
    .B(_04691_),
    .X(_01299_));
 sg13g2_mux2_1 _11258_ (.A0(\shift_storage.storage[638] ),
    .A1(\shift_storage.storage[637] ),
    .S(net524),
    .X(_04692_));
 sg13g2_and2_1 _11259_ (.A(net223),
    .B(_04692_),
    .X(_01300_));
 sg13g2_mux2_1 _11260_ (.A0(\shift_storage.storage[639] ),
    .A1(\shift_storage.storage[638] ),
    .S(net524),
    .X(_04693_));
 sg13g2_and2_1 _11261_ (.A(net223),
    .B(_04693_),
    .X(_01301_));
 sg13g2_mux2_1 _11262_ (.A0(\shift_storage.storage[63] ),
    .A1(\shift_storage.storage[62] ),
    .S(net623),
    .X(_04694_));
 sg13g2_and2_1 _11263_ (.A(net324),
    .B(_04694_),
    .X(_01302_));
 sg13g2_buf_1 fanout96 (.A(\median_processor.input_storage[56] ),
    .X(net96));
 sg13g2_mux2_1 _11265_ (.A0(\shift_storage.storage[640] ),
    .A1(\shift_storage.storage[639] ),
    .S(net524),
    .X(_04696_));
 sg13g2_and2_1 _11266_ (.A(net223),
    .B(_04696_),
    .X(_01303_));
 sg13g2_mux2_1 _11267_ (.A0(\shift_storage.storage[641] ),
    .A1(\shift_storage.storage[640] ),
    .S(net552),
    .X(_04697_));
 sg13g2_and2_1 _11268_ (.A(net251),
    .B(_04697_),
    .X(_01304_));
 sg13g2_mux2_1 _11269_ (.A0(\shift_storage.storage[642] ),
    .A1(\shift_storage.storage[641] ),
    .S(net552),
    .X(_04698_));
 sg13g2_and2_1 _11270_ (.A(net251),
    .B(_04698_),
    .X(_01305_));
 sg13g2_buf_2 fanout95 (.A(net96),
    .X(net95));
 sg13g2_mux2_1 _11272_ (.A0(\shift_storage.storage[643] ),
    .A1(\shift_storage.storage[642] ),
    .S(net552),
    .X(_04700_));
 sg13g2_and2_1 _11273_ (.A(net251),
    .B(_04700_),
    .X(_01306_));
 sg13g2_mux2_1 _11274_ (.A0(\shift_storage.storage[644] ),
    .A1(\shift_storage.storage[643] ),
    .S(net552),
    .X(_04701_));
 sg13g2_and2_1 _11275_ (.A(net251),
    .B(_04701_),
    .X(_01307_));
 sg13g2_mux2_1 _11276_ (.A0(\shift_storage.storage[645] ),
    .A1(\shift_storage.storage[644] ),
    .S(net552),
    .X(_04702_));
 sg13g2_and2_1 _11277_ (.A(net251),
    .B(_04702_),
    .X(_01308_));
 sg13g2_mux2_1 _11278_ (.A0(\shift_storage.storage[646] ),
    .A1(\shift_storage.storage[645] ),
    .S(net553),
    .X(_04703_));
 sg13g2_and2_1 _11279_ (.A(net251),
    .B(_04703_),
    .X(_01309_));
 sg13g2_mux2_1 _11280_ (.A0(\shift_storage.storage[647] ),
    .A1(\shift_storage.storage[646] ),
    .S(net553),
    .X(_04704_));
 sg13g2_and2_1 _11281_ (.A(net253),
    .B(_04704_),
    .X(_01310_));
 sg13g2_mux2_1 _11282_ (.A0(\shift_storage.storage[648] ),
    .A1(\shift_storage.storage[647] ),
    .S(net553),
    .X(_04705_));
 sg13g2_and2_1 _11283_ (.A(net253),
    .B(_04705_),
    .X(_01311_));
 sg13g2_mux2_1 _11284_ (.A0(\shift_storage.storage[649] ),
    .A1(\shift_storage.storage[648] ),
    .S(net554),
    .X(_04706_));
 sg13g2_and2_1 _11285_ (.A(net253),
    .B(_04706_),
    .X(_01312_));
 sg13g2_buf_2 fanout94 (.A(\median_processor.input_storage[57] ),
    .X(net94));
 sg13g2_mux2_1 _11287_ (.A0(\shift_storage.storage[64] ),
    .A1(\shift_storage.storage[63] ),
    .S(net623),
    .X(_04708_));
 sg13g2_and2_1 _11288_ (.A(net325),
    .B(_04708_),
    .X(_01313_));
 sg13g2_mux2_1 _11289_ (.A0(\shift_storage.storage[650] ),
    .A1(\shift_storage.storage[649] ),
    .S(net553),
    .X(_04709_));
 sg13g2_and2_1 _11290_ (.A(net253),
    .B(_04709_),
    .X(_01314_));
 sg13g2_mux2_1 _11291_ (.A0(\shift_storage.storage[651] ),
    .A1(\shift_storage.storage[650] ),
    .S(net553),
    .X(_04710_));
 sg13g2_and2_1 _11292_ (.A(net253),
    .B(_04710_),
    .X(_01315_));
 sg13g2_buf_1 fanout93 (.A(\median_processor.input_storage[58] ),
    .X(net93));
 sg13g2_mux2_1 _11294_ (.A0(\shift_storage.storage[652] ),
    .A1(\shift_storage.storage[651] ),
    .S(net553),
    .X(_04712_));
 sg13g2_and2_1 _11295_ (.A(net253),
    .B(_04712_),
    .X(_01316_));
 sg13g2_mux2_1 _11296_ (.A0(\shift_storage.storage[653] ),
    .A1(\shift_storage.storage[652] ),
    .S(net562),
    .X(_04713_));
 sg13g2_and2_1 _11297_ (.A(net262),
    .B(_04713_),
    .X(_01317_));
 sg13g2_mux2_1 _11298_ (.A0(\shift_storage.storage[654] ),
    .A1(\shift_storage.storage[653] ),
    .S(net562),
    .X(_04714_));
 sg13g2_and2_1 _11299_ (.A(net262),
    .B(_04714_),
    .X(_01318_));
 sg13g2_mux2_1 _11300_ (.A0(\shift_storage.storage[655] ),
    .A1(\shift_storage.storage[654] ),
    .S(net562),
    .X(_04715_));
 sg13g2_and2_1 _11301_ (.A(net262),
    .B(_04715_),
    .X(_01319_));
 sg13g2_mux2_1 _11302_ (.A0(\shift_storage.storage[656] ),
    .A1(\shift_storage.storage[655] ),
    .S(net562),
    .X(_04716_));
 sg13g2_and2_1 _11303_ (.A(net262),
    .B(_04716_),
    .X(_01320_));
 sg13g2_mux2_1 _11304_ (.A0(\shift_storage.storage[657] ),
    .A1(\shift_storage.storage[656] ),
    .S(net563),
    .X(_04717_));
 sg13g2_and2_1 _11305_ (.A(net262),
    .B(_04717_),
    .X(_01321_));
 sg13g2_mux2_1 _11306_ (.A0(\shift_storage.storage[658] ),
    .A1(\shift_storage.storage[657] ),
    .S(net562),
    .X(_04718_));
 sg13g2_and2_1 _11307_ (.A(net262),
    .B(_04718_),
    .X(_01322_));
 sg13g2_buf_2 fanout92 (.A(\median_processor.input_storage[58] ),
    .X(net92));
 sg13g2_mux2_1 _11309_ (.A0(\shift_storage.storage[659] ),
    .A1(\shift_storage.storage[658] ),
    .S(net562),
    .X(_04720_));
 sg13g2_and2_1 _11310_ (.A(net262),
    .B(_04720_),
    .X(_01323_));
 sg13g2_mux2_1 _11311_ (.A0(\shift_storage.storage[65] ),
    .A1(\shift_storage.storage[64] ),
    .S(net623),
    .X(_04721_));
 sg13g2_and2_1 _11312_ (.A(net325),
    .B(_04721_),
    .X(_01324_));
 sg13g2_mux2_1 _11313_ (.A0(\shift_storage.storage[660] ),
    .A1(\shift_storage.storage[659] ),
    .S(net565),
    .X(_04722_));
 sg13g2_and2_1 _11314_ (.A(net265),
    .B(_04722_),
    .X(_01325_));
 sg13g2_buf_2 fanout91 (.A(\median_processor.input_storage[59] ),
    .X(net91));
 sg13g2_mux2_1 _11316_ (.A0(\shift_storage.storage[661] ),
    .A1(\shift_storage.storage[660] ),
    .S(net565),
    .X(_04724_));
 sg13g2_and2_1 _11317_ (.A(net265),
    .B(_04724_),
    .X(_01326_));
 sg13g2_mux2_1 _11318_ (.A0(\shift_storage.storage[662] ),
    .A1(\shift_storage.storage[661] ),
    .S(net565),
    .X(_04725_));
 sg13g2_and2_1 _11319_ (.A(net265),
    .B(_04725_),
    .X(_01327_));
 sg13g2_mux2_1 _11320_ (.A0(\shift_storage.storage[663] ),
    .A1(\shift_storage.storage[662] ),
    .S(net565),
    .X(_04726_));
 sg13g2_and2_1 _11321_ (.A(net265),
    .B(_04726_),
    .X(_01328_));
 sg13g2_mux2_1 _11322_ (.A0(\shift_storage.storage[664] ),
    .A1(\shift_storage.storage[663] ),
    .S(net565),
    .X(_04727_));
 sg13g2_and2_1 _11323_ (.A(net265),
    .B(_04727_),
    .X(_01329_));
 sg13g2_mux2_1 _11324_ (.A0(\shift_storage.storage[665] ),
    .A1(\shift_storage.storage[664] ),
    .S(net565),
    .X(_04728_));
 sg13g2_and2_1 _11325_ (.A(net265),
    .B(_04728_),
    .X(_01330_));
 sg13g2_mux2_1 _11326_ (.A0(\shift_storage.storage[666] ),
    .A1(\shift_storage.storage[665] ),
    .S(net562),
    .X(_04729_));
 sg13g2_and2_1 _11327_ (.A(net263),
    .B(_04729_),
    .X(_01331_));
 sg13g2_mux2_1 _11328_ (.A0(\shift_storage.storage[667] ),
    .A1(\shift_storage.storage[666] ),
    .S(net562),
    .X(_04730_));
 sg13g2_and2_1 _11329_ (.A(net262),
    .B(_04730_),
    .X(_01332_));
 sg13g2_buf_2 fanout90 (.A(net91),
    .X(net90));
 sg13g2_mux2_1 _11331_ (.A0(\shift_storage.storage[668] ),
    .A1(\shift_storage.storage[667] ),
    .S(net558),
    .X(_04732_));
 sg13g2_and2_1 _11332_ (.A(net258),
    .B(_04732_),
    .X(_01333_));
 sg13g2_mux2_1 _11333_ (.A0(\shift_storage.storage[669] ),
    .A1(\shift_storage.storage[668] ),
    .S(net558),
    .X(_04733_));
 sg13g2_and2_1 _11334_ (.A(net258),
    .B(_04733_),
    .X(_01334_));
 sg13g2_mux2_1 _11335_ (.A0(\shift_storage.storage[66] ),
    .A1(\shift_storage.storage[65] ),
    .S(net621),
    .X(_04734_));
 sg13g2_and2_1 _11336_ (.A(net324),
    .B(_04734_),
    .X(_01335_));
 sg13g2_buf_2 fanout89 (.A(\median_processor.input_storage[5] ),
    .X(net89));
 sg13g2_mux2_1 _11338_ (.A0(\shift_storage.storage[670] ),
    .A1(\shift_storage.storage[669] ),
    .S(net558),
    .X(_04736_));
 sg13g2_and2_1 _11339_ (.A(net258),
    .B(_04736_),
    .X(_01336_));
 sg13g2_mux2_1 _11340_ (.A0(\shift_storage.storage[671] ),
    .A1(\shift_storage.storage[670] ),
    .S(net558),
    .X(_04737_));
 sg13g2_and2_1 _11341_ (.A(net249),
    .B(_04737_),
    .X(_01337_));
 sg13g2_mux2_1 _11342_ (.A0(\shift_storage.storage[672] ),
    .A1(\shift_storage.storage[671] ),
    .S(net551),
    .X(_04738_));
 sg13g2_and2_1 _11343_ (.A(net250),
    .B(_04738_),
    .X(_01338_));
 sg13g2_mux2_1 _11344_ (.A0(\shift_storage.storage[673] ),
    .A1(\shift_storage.storage[672] ),
    .S(net551),
    .X(_04739_));
 sg13g2_and2_1 _11345_ (.A(net249),
    .B(_04739_),
    .X(_01339_));
 sg13g2_mux2_1 _11346_ (.A0(\shift_storage.storage[674] ),
    .A1(\shift_storage.storage[673] ),
    .S(net550),
    .X(_04740_));
 sg13g2_and2_1 _11347_ (.A(net249),
    .B(_04740_),
    .X(_01340_));
 sg13g2_mux2_1 _11348_ (.A0(\shift_storage.storage[675] ),
    .A1(\shift_storage.storage[674] ),
    .S(net550),
    .X(_04741_));
 sg13g2_and2_1 _11349_ (.A(net253),
    .B(_04741_),
    .X(_01341_));
 sg13g2_mux2_1 _11350_ (.A0(\shift_storage.storage[676] ),
    .A1(\shift_storage.storage[675] ),
    .S(net553),
    .X(_04742_));
 sg13g2_and2_1 _11351_ (.A(net253),
    .B(_04742_),
    .X(_01342_));
 sg13g2_buf_1 fanout88 (.A(\median_processor.input_storage[60] ),
    .X(net88));
 sg13g2_mux2_1 _11353_ (.A0(\shift_storage.storage[677] ),
    .A1(\shift_storage.storage[676] ),
    .S(net553),
    .X(_04744_));
 sg13g2_and2_1 _11354_ (.A(net251),
    .B(_04744_),
    .X(_01343_));
 sg13g2_mux2_1 _11355_ (.A0(\shift_storage.storage[678] ),
    .A1(\shift_storage.storage[677] ),
    .S(net548),
    .X(_04745_));
 sg13g2_and2_1 _11356_ (.A(net247),
    .B(_04745_),
    .X(_01344_));
 sg13g2_mux2_1 _11357_ (.A0(\shift_storage.storage[679] ),
    .A1(\shift_storage.storage[678] ),
    .S(net548),
    .X(_04746_));
 sg13g2_and2_1 _11358_ (.A(net247),
    .B(_04746_),
    .X(_01345_));
 sg13g2_buf_2 fanout87 (.A(\median_processor.input_storage[60] ),
    .X(net87));
 sg13g2_mux2_1 _11360_ (.A0(\shift_storage.storage[67] ),
    .A1(\shift_storage.storage[66] ),
    .S(net631),
    .X(_04748_));
 sg13g2_and2_1 _11361_ (.A(net332),
    .B(_04748_),
    .X(_01346_));
 sg13g2_mux2_1 _11362_ (.A0(\shift_storage.storage[680] ),
    .A1(\shift_storage.storage[679] ),
    .S(net550),
    .X(_04749_));
 sg13g2_and2_1 _11363_ (.A(net249),
    .B(_04749_),
    .X(_01347_));
 sg13g2_mux2_1 _11364_ (.A0(\shift_storage.storage[681] ),
    .A1(\shift_storage.storage[680] ),
    .S(net550),
    .X(_04750_));
 sg13g2_and2_1 _11365_ (.A(net249),
    .B(_04750_),
    .X(_01348_));
 sg13g2_mux2_1 _11366_ (.A0(\shift_storage.storage[682] ),
    .A1(\shift_storage.storage[681] ),
    .S(net550),
    .X(_04751_));
 sg13g2_and2_1 _11367_ (.A(net249),
    .B(_04751_),
    .X(_01349_));
 sg13g2_mux2_1 _11368_ (.A0(\shift_storage.storage[683] ),
    .A1(\shift_storage.storage[682] ),
    .S(net549),
    .X(_04752_));
 sg13g2_and2_1 _11369_ (.A(net246),
    .B(_04752_),
    .X(_01350_));
 sg13g2_mux2_1 _11370_ (.A0(\shift_storage.storage[684] ),
    .A1(\shift_storage.storage[683] ),
    .S(net547),
    .X(_04753_));
 sg13g2_and2_1 _11371_ (.A(net246),
    .B(_04753_),
    .X(_01351_));
 sg13g2_mux2_1 _11372_ (.A0(\shift_storage.storage[685] ),
    .A1(\shift_storage.storage[684] ),
    .S(net547),
    .X(_04754_));
 sg13g2_and2_1 _11373_ (.A(net246),
    .B(_04754_),
    .X(_01352_));
 sg13g2_buf_2 fanout86 (.A(\median_processor.input_storage[61] ),
    .X(net86));
 sg13g2_mux2_1 _11375_ (.A0(\shift_storage.storage[686] ),
    .A1(\shift_storage.storage[685] ),
    .S(net547),
    .X(_04756_));
 sg13g2_and2_1 _11376_ (.A(net246),
    .B(_04756_),
    .X(_01353_));
 sg13g2_mux2_1 _11377_ (.A0(\shift_storage.storage[687] ),
    .A1(\shift_storage.storage[686] ),
    .S(net548),
    .X(_04757_));
 sg13g2_and2_1 _11378_ (.A(net247),
    .B(_04757_),
    .X(_01354_));
 sg13g2_mux2_1 _11379_ (.A0(\shift_storage.storage[688] ),
    .A1(\shift_storage.storage[687] ),
    .S(net548),
    .X(_04758_));
 sg13g2_and2_1 _11380_ (.A(net247),
    .B(_04758_),
    .X(_01355_));
 sg13g2_buf_1 fanout85 (.A(\median_processor.input_storage[62] ),
    .X(net85));
 sg13g2_mux2_1 _11382_ (.A0(\shift_storage.storage[689] ),
    .A1(\shift_storage.storage[688] ),
    .S(net548),
    .X(_04760_));
 sg13g2_and2_1 _11383_ (.A(net256),
    .B(_04760_),
    .X(_01356_));
 sg13g2_mux2_1 _11384_ (.A0(\shift_storage.storage[68] ),
    .A1(\shift_storage.storage[67] ),
    .S(net635),
    .X(_04761_));
 sg13g2_and2_1 _11385_ (.A(net337),
    .B(_04761_),
    .X(_01357_));
 sg13g2_mux2_1 _11386_ (.A0(\shift_storage.storage[690] ),
    .A1(\shift_storage.storage[689] ),
    .S(net520),
    .X(_04762_));
 sg13g2_and2_1 _11387_ (.A(net220),
    .B(_04762_),
    .X(_01358_));
 sg13g2_mux2_1 _11388_ (.A0(\shift_storage.storage[691] ),
    .A1(\shift_storage.storage[690] ),
    .S(net520),
    .X(_04763_));
 sg13g2_and2_1 _11389_ (.A(net220),
    .B(_04763_),
    .X(_01359_));
 sg13g2_mux2_1 _11390_ (.A0(\shift_storage.storage[692] ),
    .A1(\shift_storage.storage[691] ),
    .S(net520),
    .X(_04764_));
 sg13g2_and2_1 _11391_ (.A(net220),
    .B(_04764_),
    .X(_01360_));
 sg13g2_mux2_1 _11392_ (.A0(\shift_storage.storage[693] ),
    .A1(\shift_storage.storage[692] ),
    .S(net519),
    .X(_04765_));
 sg13g2_and2_1 _11393_ (.A(net220),
    .B(_04765_),
    .X(_01361_));
 sg13g2_mux2_1 _11394_ (.A0(\shift_storage.storage[694] ),
    .A1(\shift_storage.storage[693] ),
    .S(net519),
    .X(_04766_));
 sg13g2_and2_1 _11395_ (.A(net219),
    .B(_04766_),
    .X(_01362_));
 sg13g2_buf_2 fanout84 (.A(\median_processor.input_storage[62] ),
    .X(net84));
 sg13g2_buf_2 fanout83 (.A(\median_processor.input_storage[63] ),
    .X(net83));
 sg13g2_mux2_1 _11398_ (.A0(\shift_storage.storage[695] ),
    .A1(\shift_storage.storage[694] ),
    .S(net520),
    .X(_04769_));
 sg13g2_and2_1 _11399_ (.A(net219),
    .B(_04769_),
    .X(_01363_));
 sg13g2_mux2_1 _11400_ (.A0(\shift_storage.storage[696] ),
    .A1(\shift_storage.storage[695] ),
    .S(net519),
    .X(_04770_));
 sg13g2_and2_1 _11401_ (.A(net219),
    .B(_04770_),
    .X(_01364_));
 sg13g2_mux2_1 _11402_ (.A0(\shift_storage.storage[697] ),
    .A1(\shift_storage.storage[696] ),
    .S(net519),
    .X(_04771_));
 sg13g2_and2_1 _11403_ (.A(net219),
    .B(_04771_),
    .X(_01365_));
 sg13g2_buf_2 fanout82 (.A(net83),
    .X(net82));
 sg13g2_buf_2 fanout81 (.A(\median_processor.input_storage[6] ),
    .X(net81));
 sg13g2_mux2_1 _11406_ (.A0(\shift_storage.storage[698] ),
    .A1(\shift_storage.storage[697] ),
    .S(net547),
    .X(_04774_));
 sg13g2_and2_1 _11407_ (.A(net246),
    .B(_04774_),
    .X(_01366_));
 sg13g2_mux2_1 _11408_ (.A0(\shift_storage.storage[699] ),
    .A1(\shift_storage.storage[698] ),
    .S(net547),
    .X(_04775_));
 sg13g2_and2_1 _11409_ (.A(net246),
    .B(_04775_),
    .X(_01367_));
 sg13g2_mux2_1 _11410_ (.A0(\shift_storage.storage[69] ),
    .A1(\shift_storage.storage[68] ),
    .S(net635),
    .X(_04776_));
 sg13g2_and2_1 _11411_ (.A(net337),
    .B(_04776_),
    .X(_01368_));
 sg13g2_mux2_1 _11412_ (.A0(\shift_storage.storage[6] ),
    .A1(\shift_storage.storage[5] ),
    .S(net612),
    .X(_04777_));
 sg13g2_and2_1 _11413_ (.A(net310),
    .B(_04777_),
    .X(_01369_));
 sg13g2_mux2_1 _11414_ (.A0(\shift_storage.storage[700] ),
    .A1(\shift_storage.storage[699] ),
    .S(net547),
    .X(_04778_));
 sg13g2_and2_1 _11415_ (.A(net247),
    .B(_04778_),
    .X(_01370_));
 sg13g2_mux2_1 _11416_ (.A0(\shift_storage.storage[701] ),
    .A1(\shift_storage.storage[700] ),
    .S(net547),
    .X(_04779_));
 sg13g2_and2_1 _11417_ (.A(net246),
    .B(_04779_),
    .X(_01371_));
 sg13g2_mux2_1 _11418_ (.A0(\shift_storage.storage[702] ),
    .A1(\shift_storage.storage[701] ),
    .S(net547),
    .X(_04780_));
 sg13g2_and2_1 _11419_ (.A(net246),
    .B(_04780_),
    .X(_01372_));
 sg13g2_buf_2 fanout80 (.A(net81),
    .X(net80));
 sg13g2_mux2_1 _11421_ (.A0(\shift_storage.storage[703] ),
    .A1(\shift_storage.storage[702] ),
    .S(net549),
    .X(_04782_));
 sg13g2_and2_1 _11422_ (.A(net248),
    .B(_04782_),
    .X(_01373_));
 sg13g2_mux2_1 _11423_ (.A0(\shift_storage.storage[704] ),
    .A1(\shift_storage.storage[703] ),
    .S(net549),
    .X(_04783_));
 sg13g2_and2_1 _11424_ (.A(net248),
    .B(_04783_),
    .X(_01374_));
 sg13g2_mux2_1 _11425_ (.A0(\shift_storage.storage[705] ),
    .A1(\shift_storage.storage[704] ),
    .S(net549),
    .X(_04784_));
 sg13g2_and2_1 _11426_ (.A(net250),
    .B(_04784_),
    .X(_01375_));
 sg13g2_buf_1 fanout79 (.A(\median_processor.input_storage[7] ),
    .X(net79));
 sg13g2_mux2_1 _11428_ (.A0(\shift_storage.storage[706] ),
    .A1(\shift_storage.storage[705] ),
    .S(net549),
    .X(_04786_));
 sg13g2_and2_1 _11429_ (.A(net248),
    .B(_04786_),
    .X(_01376_));
 sg13g2_mux2_1 _11430_ (.A0(\shift_storage.storage[707] ),
    .A1(\shift_storage.storage[706] ),
    .S(net549),
    .X(_04787_));
 sg13g2_and2_1 _11431_ (.A(net248),
    .B(_04787_),
    .X(_01377_));
 sg13g2_mux2_1 _11432_ (.A0(\shift_storage.storage[708] ),
    .A1(\shift_storage.storage[707] ),
    .S(net557),
    .X(_04788_));
 sg13g2_and2_1 _11433_ (.A(net248),
    .B(_04788_),
    .X(_01378_));
 sg13g2_mux2_1 _11434_ (.A0(\shift_storage.storage[709] ),
    .A1(\shift_storage.storage[708] ),
    .S(net549),
    .X(_04789_));
 sg13g2_and2_1 _11435_ (.A(net248),
    .B(_04789_),
    .X(_01379_));
 sg13g2_mux2_1 _11436_ (.A0(\shift_storage.storage[70] ),
    .A1(\shift_storage.storage[69] ),
    .S(net635),
    .X(_04790_));
 sg13g2_and2_1 _11437_ (.A(net337),
    .B(_04790_),
    .X(_01380_));
 sg13g2_mux2_1 _11438_ (.A0(\shift_storage.storage[710] ),
    .A1(\shift_storage.storage[709] ),
    .S(net551),
    .X(_04791_));
 sg13g2_and2_1 _11439_ (.A(net250),
    .B(_04791_),
    .X(_01381_));
 sg13g2_mux2_1 _11440_ (.A0(\shift_storage.storage[711] ),
    .A1(\shift_storage.storage[710] ),
    .S(net551),
    .X(_04792_));
 sg13g2_and2_1 _11441_ (.A(net248),
    .B(_04792_),
    .X(_01382_));
 sg13g2_buf_1 fanout78 (.A(net79),
    .X(net78));
 sg13g2_mux2_1 _11443_ (.A0(\shift_storage.storage[712] ),
    .A1(\shift_storage.storage[711] ),
    .S(net549),
    .X(_04794_));
 sg13g2_and2_1 _11444_ (.A(net248),
    .B(_04794_),
    .X(_01383_));
 sg13g2_mux2_1 _11445_ (.A0(\shift_storage.storage[713] ),
    .A1(\shift_storage.storage[712] ),
    .S(net550),
    .X(_04795_));
 sg13g2_and2_1 _11446_ (.A(net249),
    .B(_04795_),
    .X(_01384_));
 sg13g2_mux2_1 _11447_ (.A0(\shift_storage.storage[714] ),
    .A1(\shift_storage.storage[713] ),
    .S(net550),
    .X(_04796_));
 sg13g2_and2_1 _11448_ (.A(net250),
    .B(_04796_),
    .X(_01385_));
 sg13g2_buf_2 fanout77 (.A(net79),
    .X(net77));
 sg13g2_mux2_1 _11450_ (.A0(\shift_storage.storage[715] ),
    .A1(\shift_storage.storage[714] ),
    .S(net550),
    .X(_04798_));
 sg13g2_and2_1 _11451_ (.A(net249),
    .B(_04798_),
    .X(_01386_));
 sg13g2_mux2_1 _11452_ (.A0(\shift_storage.storage[716] ),
    .A1(\shift_storage.storage[715] ),
    .S(net558),
    .X(_04799_));
 sg13g2_and2_1 _11453_ (.A(net257),
    .B(_04799_),
    .X(_01387_));
 sg13g2_mux2_1 _11454_ (.A0(\shift_storage.storage[717] ),
    .A1(\shift_storage.storage[716] ),
    .S(net558),
    .X(_04800_));
 sg13g2_and2_1 _11455_ (.A(net258),
    .B(_04800_),
    .X(_01388_));
 sg13g2_mux2_1 _11456_ (.A0(\shift_storage.storage[718] ),
    .A1(\shift_storage.storage[717] ),
    .S(net557),
    .X(_04801_));
 sg13g2_and2_1 _11457_ (.A(net257),
    .B(_04801_),
    .X(_01389_));
 sg13g2_mux2_1 _11458_ (.A0(\shift_storage.storage[719] ),
    .A1(\shift_storage.storage[718] ),
    .S(net557),
    .X(_04802_));
 sg13g2_and2_1 _11459_ (.A(net257),
    .B(_04802_),
    .X(_01390_));
 sg13g2_mux2_1 _11460_ (.A0(\shift_storage.storage[71] ),
    .A1(\shift_storage.storage[70] ),
    .S(net627),
    .X(_04803_));
 sg13g2_and2_1 _11461_ (.A(net329),
    .B(_04803_),
    .X(_01391_));
 sg13g2_mux2_1 _11462_ (.A0(\shift_storage.storage[720] ),
    .A1(\shift_storage.storage[719] ),
    .S(net557),
    .X(_04804_));
 sg13g2_and2_1 _11463_ (.A(net257),
    .B(_04804_),
    .X(_01392_));
 sg13g2_buf_2 fanout76 (.A(\median_processor.input_storage[8] ),
    .X(net76));
 sg13g2_mux2_1 _11465_ (.A0(\shift_storage.storage[721] ),
    .A1(\shift_storage.storage[720] ),
    .S(net557),
    .X(_04806_));
 sg13g2_and2_1 _11466_ (.A(net257),
    .B(_04806_),
    .X(_01393_));
 sg13g2_mux2_1 _11467_ (.A0(\shift_storage.storage[722] ),
    .A1(\shift_storage.storage[721] ),
    .S(net557),
    .X(_04807_));
 sg13g2_and2_1 _11468_ (.A(net257),
    .B(_04807_),
    .X(_01394_));
 sg13g2_mux2_1 _11469_ (.A0(\shift_storage.storage[723] ),
    .A1(\shift_storage.storage[722] ),
    .S(net557),
    .X(_04808_));
 sg13g2_and2_1 _11470_ (.A(net257),
    .B(_04808_),
    .X(_01395_));
 sg13g2_buf_2 fanout75 (.A(net76),
    .X(net75));
 sg13g2_mux2_1 _11472_ (.A0(\shift_storage.storage[724] ),
    .A1(\shift_storage.storage[723] ),
    .S(net557),
    .X(_04810_));
 sg13g2_and2_1 _11473_ (.A(net257),
    .B(_04810_),
    .X(_01396_));
 sg13g2_mux2_1 _11474_ (.A0(\shift_storage.storage[725] ),
    .A1(\shift_storage.storage[724] ),
    .S(net559),
    .X(_04811_));
 sg13g2_and2_1 _11475_ (.A(net259),
    .B(_04811_),
    .X(_01397_));
 sg13g2_mux2_1 _11476_ (.A0(\shift_storage.storage[726] ),
    .A1(\shift_storage.storage[725] ),
    .S(net559),
    .X(_04812_));
 sg13g2_and2_1 _11477_ (.A(net259),
    .B(_04812_),
    .X(_01398_));
 sg13g2_mux2_1 _11478_ (.A0(\shift_storage.storage[727] ),
    .A1(\shift_storage.storage[726] ),
    .S(net561),
    .X(_04813_));
 sg13g2_and2_1 _11479_ (.A(net261),
    .B(_04813_),
    .X(_01399_));
 sg13g2_mux2_1 _11480_ (.A0(\shift_storage.storage[728] ),
    .A1(\shift_storage.storage[727] ),
    .S(net559),
    .X(_04814_));
 sg13g2_and2_1 _11481_ (.A(net259),
    .B(_04814_),
    .X(_01400_));
 sg13g2_mux2_1 _11482_ (.A0(\shift_storage.storage[729] ),
    .A1(\shift_storage.storage[728] ),
    .S(net655),
    .X(_04815_));
 sg13g2_and2_1 _11483_ (.A(net357),
    .B(_04815_),
    .X(_01401_));
 sg13g2_mux2_1 _11484_ (.A0(\shift_storage.storage[72] ),
    .A1(\shift_storage.storage[71] ),
    .S(net627),
    .X(_04816_));
 sg13g2_and2_1 _11485_ (.A(net329),
    .B(_04816_),
    .X(_01402_));
 sg13g2_buf_2 fanout74 (.A(\median_processor.input_storage[9] ),
    .X(net74));
 sg13g2_mux2_1 _11487_ (.A0(\shift_storage.storage[730] ),
    .A1(\shift_storage.storage[729] ),
    .S(net655),
    .X(_04818_));
 sg13g2_and2_1 _11488_ (.A(net357),
    .B(_04818_),
    .X(_01403_));
 sg13g2_mux2_1 _11489_ (.A0(\shift_storage.storage[731] ),
    .A1(\shift_storage.storage[730] ),
    .S(net559),
    .X(_04819_));
 sg13g2_and2_1 _11490_ (.A(net259),
    .B(_04819_),
    .X(_01404_));
 sg13g2_mux2_1 _11491_ (.A0(\shift_storage.storage[732] ),
    .A1(\shift_storage.storage[731] ),
    .S(net559),
    .X(_04820_));
 sg13g2_and2_1 _11492_ (.A(net259),
    .B(_04820_),
    .X(_01405_));
 sg13g2_buf_2 fanout73 (.A(_01741_),
    .X(net73));
 sg13g2_mux2_1 _11494_ (.A0(\shift_storage.storage[733] ),
    .A1(\shift_storage.storage[732] ),
    .S(net559),
    .X(_04822_));
 sg13g2_and2_1 _11495_ (.A(net259),
    .B(_04822_),
    .X(_01406_));
 sg13g2_mux2_1 _11496_ (.A0(\shift_storage.storage[734] ),
    .A1(\shift_storage.storage[733] ),
    .S(net559),
    .X(_04823_));
 sg13g2_and2_1 _11497_ (.A(net259),
    .B(_04823_),
    .X(_01407_));
 sg13g2_mux2_1 _11498_ (.A0(\shift_storage.storage[735] ),
    .A1(\shift_storage.storage[734] ),
    .S(net560),
    .X(_04824_));
 sg13g2_and2_1 _11499_ (.A(net260),
    .B(_04824_),
    .X(_01408_));
 sg13g2_mux2_1 _11500_ (.A0(\shift_storage.storage[736] ),
    .A1(\shift_storage.storage[735] ),
    .S(net560),
    .X(_04825_));
 sg13g2_and2_1 _11501_ (.A(net260),
    .B(_04825_),
    .X(_01409_));
 sg13g2_mux2_1 _11502_ (.A0(\shift_storage.storage[737] ),
    .A1(\shift_storage.storage[736] ),
    .S(net560),
    .X(_04826_));
 sg13g2_and2_1 _11503_ (.A(net260),
    .B(_04826_),
    .X(_01410_));
 sg13g2_mux2_1 _11504_ (.A0(\shift_storage.storage[738] ),
    .A1(\shift_storage.storage[737] ),
    .S(net560),
    .X(_04827_));
 sg13g2_and2_1 _11505_ (.A(net260),
    .B(_04827_),
    .X(_01411_));
 sg13g2_mux2_1 _11506_ (.A0(\shift_storage.storage[739] ),
    .A1(\shift_storage.storage[738] ),
    .S(net560),
    .X(_04828_));
 sg13g2_and2_1 _11507_ (.A(net260),
    .B(_04828_),
    .X(_01412_));
 sg13g2_buf_2 fanout72 (.A(_01755_),
    .X(net72));
 sg13g2_mux2_1 _11509_ (.A0(\shift_storage.storage[73] ),
    .A1(\shift_storage.storage[72] ),
    .S(net628),
    .X(_04830_));
 sg13g2_and2_1 _11510_ (.A(net330),
    .B(_04830_),
    .X(_01413_));
 sg13g2_mux2_1 _11511_ (.A0(\shift_storage.storage[740] ),
    .A1(\shift_storage.storage[739] ),
    .S(net560),
    .X(_04831_));
 sg13g2_and2_1 _11512_ (.A(net260),
    .B(_04831_),
    .X(_01414_));
 sg13g2_mux2_1 _11513_ (.A0(\shift_storage.storage[741] ),
    .A1(\shift_storage.storage[740] ),
    .S(net561),
    .X(_04832_));
 sg13g2_and2_1 _11514_ (.A(net261),
    .B(_04832_),
    .X(_01415_));
 sg13g2_buf_2 fanout71 (.A(_01765_),
    .X(net71));
 sg13g2_mux2_1 _11516_ (.A0(\shift_storage.storage[742] ),
    .A1(\shift_storage.storage[741] ),
    .S(net565),
    .X(_04834_));
 sg13g2_and2_1 _11517_ (.A(net265),
    .B(_04834_),
    .X(_01416_));
 sg13g2_mux2_1 _11518_ (.A0(\shift_storage.storage[743] ),
    .A1(\shift_storage.storage[742] ),
    .S(net657),
    .X(_04835_));
 sg13g2_and2_1 _11519_ (.A(net361),
    .B(_04835_),
    .X(_01417_));
 sg13g2_mux2_1 _11520_ (.A0(\shift_storage.storage[744] ),
    .A1(\shift_storage.storage[743] ),
    .S(net657),
    .X(_04836_));
 sg13g2_and2_1 _11521_ (.A(net361),
    .B(_04836_),
    .X(_01418_));
 sg13g2_mux2_1 _11522_ (.A0(\shift_storage.storage[745] ),
    .A1(\shift_storage.storage[744] ),
    .S(net657),
    .X(_04837_));
 sg13g2_and2_1 _11523_ (.A(net361),
    .B(_04837_),
    .X(_01419_));
 sg13g2_mux2_1 _11524_ (.A0(\shift_storage.storage[746] ),
    .A1(\shift_storage.storage[745] ),
    .S(net657),
    .X(_04838_));
 sg13g2_and2_1 _11525_ (.A(net361),
    .B(_04838_),
    .X(_01420_));
 sg13g2_mux2_1 _11526_ (.A0(\shift_storage.storage[747] ),
    .A1(\shift_storage.storage[746] ),
    .S(net657),
    .X(_04839_));
 sg13g2_and2_1 _11527_ (.A(net361),
    .B(_04839_),
    .X(_01421_));
 sg13g2_mux2_1 _11528_ (.A0(\shift_storage.storage[748] ),
    .A1(\shift_storage.storage[747] ),
    .S(net657),
    .X(_04840_));
 sg13g2_and2_1 _11529_ (.A(net362),
    .B(_04840_),
    .X(_01422_));
 sg13g2_buf_2 fanout70 (.A(_01773_),
    .X(net70));
 sg13g2_mux2_1 _11531_ (.A0(\shift_storage.storage[749] ),
    .A1(\shift_storage.storage[748] ),
    .S(net657),
    .X(_04842_));
 sg13g2_and2_1 _11532_ (.A(net362),
    .B(_04842_),
    .X(_01423_));
 sg13g2_mux2_1 _11533_ (.A0(\shift_storage.storage[74] ),
    .A1(\shift_storage.storage[73] ),
    .S(net628),
    .X(_04843_));
 sg13g2_and2_1 _11534_ (.A(net330),
    .B(_04843_),
    .X(_01424_));
 sg13g2_mux2_1 _11535_ (.A0(\shift_storage.storage[750] ),
    .A1(\shift_storage.storage[749] ),
    .S(net657),
    .X(_04844_));
 sg13g2_and2_1 _11536_ (.A(net362),
    .B(_04844_),
    .X(_01425_));
 sg13g2_buf_2 fanout69 (.A(_01781_),
    .X(net69));
 sg13g2_mux2_1 _11538_ (.A0(\shift_storage.storage[751] ),
    .A1(\shift_storage.storage[750] ),
    .S(net659),
    .X(_04846_));
 sg13g2_and2_1 _11539_ (.A(net361),
    .B(_04846_),
    .X(_01426_));
 sg13g2_mux2_1 _11540_ (.A0(\shift_storage.storage[752] ),
    .A1(\shift_storage.storage[751] ),
    .S(net659),
    .X(_04847_));
 sg13g2_and2_1 _11541_ (.A(net361),
    .B(_04847_),
    .X(_01427_));
 sg13g2_mux2_1 _11542_ (.A0(\shift_storage.storage[753] ),
    .A1(\shift_storage.storage[752] ),
    .S(net659),
    .X(_04848_));
 sg13g2_and2_1 _11543_ (.A(net361),
    .B(_04848_),
    .X(_01428_));
 sg13g2_mux2_1 _11544_ (.A0(\shift_storage.storage[754] ),
    .A1(\shift_storage.storage[753] ),
    .S(net656),
    .X(_04849_));
 sg13g2_and2_1 _11545_ (.A(net359),
    .B(_04849_),
    .X(_01429_));
 sg13g2_mux2_1 _11546_ (.A0(\shift_storage.storage[755] ),
    .A1(\shift_storage.storage[754] ),
    .S(net654),
    .X(_04850_));
 sg13g2_and2_1 _11547_ (.A(net357),
    .B(_04850_),
    .X(_01430_));
 sg13g2_mux2_1 _11548_ (.A0(\shift_storage.storage[756] ),
    .A1(\shift_storage.storage[755] ),
    .S(net654),
    .X(_04851_));
 sg13g2_and2_1 _11549_ (.A(net358),
    .B(_04851_),
    .X(_01431_));
 sg13g2_mux2_1 _11550_ (.A0(\shift_storage.storage[757] ),
    .A1(\shift_storage.storage[756] ),
    .S(net655),
    .X(_04852_));
 sg13g2_and2_1 _11551_ (.A(net358),
    .B(_04852_),
    .X(_01432_));
 sg13g2_buf_2 fanout68 (.A(_01796_),
    .X(net68));
 sg13g2_buf_1 fanout67 (.A(_01814_),
    .X(net67));
 sg13g2_mux2_1 _11554_ (.A0(\shift_storage.storage[758] ),
    .A1(\shift_storage.storage[757] ),
    .S(net654),
    .X(_04855_));
 sg13g2_and2_1 _11555_ (.A(net358),
    .B(_04855_),
    .X(_01433_));
 sg13g2_mux2_1 _11556_ (.A0(\shift_storage.storage[759] ),
    .A1(\shift_storage.storage[758] ),
    .S(net654),
    .X(_04856_));
 sg13g2_and2_1 _11557_ (.A(net357),
    .B(_04856_),
    .X(_01434_));
 sg13g2_mux2_1 _11558_ (.A0(\shift_storage.storage[75] ),
    .A1(\shift_storage.storage[74] ),
    .S(net639),
    .X(_04857_));
 sg13g2_and2_1 _11559_ (.A(net338),
    .B(_04857_),
    .X(_01435_));
 sg13g2_buf_2 fanout66 (.A(net67),
    .X(net66));
 sg13g2_buf_1 fanout65 (.A(_01822_),
    .X(net65));
 sg13g2_mux2_1 _11562_ (.A0(\shift_storage.storage[760] ),
    .A1(\shift_storage.storage[759] ),
    .S(net654),
    .X(_04860_));
 sg13g2_and2_1 _11563_ (.A(net260),
    .B(_04860_),
    .X(_01436_));
 sg13g2_mux2_1 _11564_ (.A0(\shift_storage.storage[761] ),
    .A1(\shift_storage.storage[760] ),
    .S(net560),
    .X(_04861_));
 sg13g2_and2_1 _11565_ (.A(net260),
    .B(_04861_),
    .X(_01437_));
 sg13g2_mux2_1 _11566_ (.A0(\shift_storage.storage[762] ),
    .A1(\shift_storage.storage[761] ),
    .S(net560),
    .X(_04862_));
 sg13g2_and2_1 _11567_ (.A(net261),
    .B(_04862_),
    .X(_01438_));
 sg13g2_mux2_1 _11568_ (.A0(\shift_storage.storage[763] ),
    .A1(\shift_storage.storage[762] ),
    .S(net559),
    .X(_04863_));
 sg13g2_and2_1 _11569_ (.A(net259),
    .B(_04863_),
    .X(_01439_));
 sg13g2_mux2_1 _11570_ (.A0(\shift_storage.storage[764] ),
    .A1(\shift_storage.storage[763] ),
    .S(net655),
    .X(_04864_));
 sg13g2_and2_1 _11571_ (.A(net357),
    .B(_04864_),
    .X(_01440_));
 sg13g2_mux2_1 _11572_ (.A0(\shift_storage.storage[765] ),
    .A1(\shift_storage.storage[764] ),
    .S(net655),
    .X(_04865_));
 sg13g2_and2_1 _11573_ (.A(net357),
    .B(_04865_),
    .X(_01441_));
 sg13g2_mux2_1 _11574_ (.A0(\shift_storage.storage[766] ),
    .A1(\shift_storage.storage[765] ),
    .S(net655),
    .X(_04866_));
 sg13g2_and2_1 _11575_ (.A(net357),
    .B(_04866_),
    .X(_01442_));
 sg13g2_buf_2 fanout64 (.A(net65),
    .X(net64));
 sg13g2_mux2_1 _11577_ (.A0(\shift_storage.storage[767] ),
    .A1(\shift_storage.storage[766] ),
    .S(net654),
    .X(_04868_));
 sg13g2_and2_1 _11578_ (.A(net358),
    .B(_04868_),
    .X(_01443_));
 sg13g2_mux2_1 _11579_ (.A0(\shift_storage.storage[768] ),
    .A1(\shift_storage.storage[767] ),
    .S(net654),
    .X(_04869_));
 sg13g2_and2_1 _11580_ (.A(net358),
    .B(_04869_),
    .X(_01444_));
 sg13g2_mux2_1 _11581_ (.A0(\shift_storage.storage[769] ),
    .A1(\shift_storage.storage[768] ),
    .S(net654),
    .X(_04870_));
 sg13g2_and2_1 _11582_ (.A(net357),
    .B(_04870_),
    .X(_01445_));
 sg13g2_buf_2 fanout63 (.A(_01922_),
    .X(net63));
 sg13g2_mux2_1 _11584_ (.A0(\shift_storage.storage[76] ),
    .A1(\shift_storage.storage[75] ),
    .S(net636),
    .X(_04872_));
 sg13g2_and2_1 _11585_ (.A(net338),
    .B(_04872_),
    .X(_01446_));
 sg13g2_mux2_1 _11586_ (.A0(\shift_storage.storage[770] ),
    .A1(\shift_storage.storage[769] ),
    .S(net656),
    .X(_04873_));
 sg13g2_and2_1 _11587_ (.A(net359),
    .B(_04873_),
    .X(_01447_));
 sg13g2_mux2_1 _11588_ (.A0(\shift_storage.storage[771] ),
    .A1(\shift_storage.storage[770] ),
    .S(net656),
    .X(_04874_));
 sg13g2_and2_1 _11589_ (.A(net359),
    .B(_04874_),
    .X(_01448_));
 sg13g2_mux2_1 _11590_ (.A0(\shift_storage.storage[772] ),
    .A1(\shift_storage.storage[771] ),
    .S(net662),
    .X(_04875_));
 sg13g2_and2_1 _11591_ (.A(net359),
    .B(_04875_),
    .X(_01449_));
 sg13g2_mux2_1 _11592_ (.A0(\shift_storage.storage[773] ),
    .A1(\shift_storage.storage[772] ),
    .S(net656),
    .X(_04876_));
 sg13g2_and2_1 _11593_ (.A(net359),
    .B(_04876_),
    .X(_01450_));
 sg13g2_mux2_1 _11594_ (.A0(\shift_storage.storage[774] ),
    .A1(\shift_storage.storage[773] ),
    .S(net656),
    .X(_04877_));
 sg13g2_and2_1 _11595_ (.A(net359),
    .B(_04877_),
    .X(_01451_));
 sg13g2_mux2_1 _11596_ (.A0(\shift_storage.storage[775] ),
    .A1(\shift_storage.storage[774] ),
    .S(net663),
    .X(_04878_));
 sg13g2_and2_1 _11597_ (.A(net367),
    .B(_04878_),
    .X(_01452_));
 sg13g2_buf_2 fanout62 (.A(_01926_),
    .X(net62));
 sg13g2_mux2_1 _11599_ (.A0(\shift_storage.storage[776] ),
    .A1(\shift_storage.storage[775] ),
    .S(net663),
    .X(_04880_));
 sg13g2_and2_1 _11600_ (.A(net367),
    .B(_04880_),
    .X(_01453_));
 sg13g2_mux2_1 _11601_ (.A0(\shift_storage.storage[777] ),
    .A1(\shift_storage.storage[776] ),
    .S(net666),
    .X(_04881_));
 sg13g2_and2_1 _11602_ (.A(net367),
    .B(_04881_),
    .X(_01454_));
 sg13g2_mux2_1 _11603_ (.A0(\shift_storage.storage[778] ),
    .A1(\shift_storage.storage[777] ),
    .S(net666),
    .X(_04882_));
 sg13g2_and2_1 _11604_ (.A(net368),
    .B(_04882_),
    .X(_01455_));
 sg13g2_buf_2 fanout61 (.A(_01945_),
    .X(net61));
 sg13g2_mux2_1 _11606_ (.A0(\shift_storage.storage[779] ),
    .A1(\shift_storage.storage[778] ),
    .S(net663),
    .X(_04884_));
 sg13g2_and2_1 _11607_ (.A(net367),
    .B(_04884_),
    .X(_01456_));
 sg13g2_mux2_1 _11608_ (.A0(\shift_storage.storage[77] ),
    .A1(\shift_storage.storage[76] ),
    .S(net636),
    .X(_04885_));
 sg13g2_and2_1 _11609_ (.A(net338),
    .B(_04885_),
    .X(_01457_));
 sg13g2_mux2_1 _11610_ (.A0(\shift_storage.storage[780] ),
    .A1(\shift_storage.storage[779] ),
    .S(net663),
    .X(_04886_));
 sg13g2_and2_1 _11611_ (.A(net367),
    .B(_04886_),
    .X(_01458_));
 sg13g2_mux2_1 _11612_ (.A0(\shift_storage.storage[781] ),
    .A1(\shift_storage.storage[780] ),
    .S(net667),
    .X(_04887_));
 sg13g2_and2_1 _11613_ (.A(net371),
    .B(_04887_),
    .X(_01459_));
 sg13g2_mux2_1 _11614_ (.A0(\shift_storage.storage[782] ),
    .A1(\shift_storage.storage[781] ),
    .S(net667),
    .X(_04888_));
 sg13g2_and2_1 _11615_ (.A(net371),
    .B(_04888_),
    .X(_01460_));
 sg13g2_mux2_1 _11616_ (.A0(\shift_storage.storage[783] ),
    .A1(\shift_storage.storage[782] ),
    .S(net668),
    .X(_04889_));
 sg13g2_and2_1 _11617_ (.A(net372),
    .B(_04889_),
    .X(_01461_));
 sg13g2_mux2_1 _11618_ (.A0(\shift_storage.storage[784] ),
    .A1(\shift_storage.storage[783] ),
    .S(net667),
    .X(_04890_));
 sg13g2_and2_1 _11619_ (.A(net371),
    .B(_04890_),
    .X(_01462_));
 sg13g2_buf_2 fanout60 (.A(_01982_),
    .X(net60));
 sg13g2_mux2_1 _11621_ (.A0(\shift_storage.storage[785] ),
    .A1(\shift_storage.storage[784] ),
    .S(net667),
    .X(_04892_));
 sg13g2_and2_1 _11622_ (.A(net371),
    .B(_04892_),
    .X(_01463_));
 sg13g2_mux2_1 _11623_ (.A0(\shift_storage.storage[786] ),
    .A1(\shift_storage.storage[785] ),
    .S(net667),
    .X(_04893_));
 sg13g2_and2_1 _11624_ (.A(net371),
    .B(_04893_),
    .X(_01464_));
 sg13g2_mux2_1 _11625_ (.A0(\shift_storage.storage[787] ),
    .A1(\shift_storage.storage[786] ),
    .S(net666),
    .X(_04894_));
 sg13g2_and2_1 _11626_ (.A(net367),
    .B(_04894_),
    .X(_01465_));
 sg13g2_buf_2 fanout59 (.A(_02006_),
    .X(net59));
 sg13g2_mux2_1 _11628_ (.A0(\shift_storage.storage[788] ),
    .A1(\shift_storage.storage[787] ),
    .S(net656),
    .X(_04896_));
 sg13g2_and2_1 _11629_ (.A(net360),
    .B(_04896_),
    .X(_01466_));
 sg13g2_mux2_1 _11630_ (.A0(\shift_storage.storage[789] ),
    .A1(\shift_storage.storage[788] ),
    .S(net656),
    .X(_04897_));
 sg13g2_and2_1 _11631_ (.A(net359),
    .B(_04897_),
    .X(_01467_));
 sg13g2_mux2_1 _11632_ (.A0(\shift_storage.storage[78] ),
    .A1(\shift_storage.storage[77] ),
    .S(net639),
    .X(_04898_));
 sg13g2_and2_1 _11633_ (.A(net338),
    .B(_04898_),
    .X(_01468_));
 sg13g2_mux2_1 _11634_ (.A0(\shift_storage.storage[790] ),
    .A1(\shift_storage.storage[789] ),
    .S(net656),
    .X(_04899_));
 sg13g2_and2_1 _11635_ (.A(net359),
    .B(_04899_),
    .X(_01469_));
 sg13g2_mux2_1 _11636_ (.A0(\shift_storage.storage[791] ),
    .A1(\shift_storage.storage[790] ),
    .S(net659),
    .X(_04900_));
 sg13g2_and2_1 _11637_ (.A(net364),
    .B(_04900_),
    .X(_01470_));
 sg13g2_mux2_1 _11638_ (.A0(\shift_storage.storage[792] ),
    .A1(\shift_storage.storage[791] ),
    .S(net659),
    .X(_04901_));
 sg13g2_and2_1 _11639_ (.A(net364),
    .B(_04901_),
    .X(_01471_));
 sg13g2_mux2_1 _11640_ (.A0(\shift_storage.storage[793] ),
    .A1(\shift_storage.storage[792] ),
    .S(net659),
    .X(_04902_));
 sg13g2_and2_1 _11641_ (.A(net364),
    .B(_04902_),
    .X(_01472_));
 sg13g2_buf_2 fanout58 (.A(_02042_),
    .X(net58));
 sg13g2_mux2_1 _11643_ (.A0(\shift_storage.storage[794] ),
    .A1(\shift_storage.storage[793] ),
    .S(net659),
    .X(_04904_));
 sg13g2_and2_1 _11644_ (.A(net364),
    .B(_04904_),
    .X(_01473_));
 sg13g2_mux2_1 _11645_ (.A0(\shift_storage.storage[795] ),
    .A1(\shift_storage.storage[794] ),
    .S(net659),
    .X(_04905_));
 sg13g2_and2_1 _11646_ (.A(net364),
    .B(_04905_),
    .X(_01474_));
 sg13g2_mux2_1 _11647_ (.A0(\shift_storage.storage[796] ),
    .A1(\shift_storage.storage[795] ),
    .S(net660),
    .X(_04906_));
 sg13g2_and2_1 _11648_ (.A(net365),
    .B(_04906_),
    .X(_01475_));
 sg13g2_buf_2 fanout57 (.A(_02058_),
    .X(net57));
 sg13g2_mux2_1 _11650_ (.A0(\shift_storage.storage[797] ),
    .A1(\shift_storage.storage[796] ),
    .S(net660),
    .X(_04908_));
 sg13g2_and2_1 _11651_ (.A(net365),
    .B(_04908_),
    .X(_01476_));
 sg13g2_mux2_1 _11652_ (.A0(\shift_storage.storage[798] ),
    .A1(\shift_storage.storage[797] ),
    .S(net660),
    .X(_04909_));
 sg13g2_and2_1 _11653_ (.A(net365),
    .B(_04909_),
    .X(_01477_));
 sg13g2_mux2_1 _11654_ (.A0(\shift_storage.storage[799] ),
    .A1(\shift_storage.storage[798] ),
    .S(net660),
    .X(_04910_));
 sg13g2_and2_1 _11655_ (.A(net364),
    .B(_04910_),
    .X(_01478_));
 sg13g2_mux2_1 _11656_ (.A0(\shift_storage.storage[79] ),
    .A1(\shift_storage.storage[78] ),
    .S(net647),
    .X(_04911_));
 sg13g2_and2_1 _11657_ (.A(net345),
    .B(_04911_),
    .X(_01479_));
 sg13g2_mux2_1 _11658_ (.A0(\shift_storage.storage[7] ),
    .A1(\shift_storage.storage[6] ),
    .S(net608),
    .X(_04912_));
 sg13g2_and2_1 _11659_ (.A(net313),
    .B(_04912_),
    .X(_01480_));
 sg13g2_mux2_1 _11660_ (.A0(\shift_storage.storage[800] ),
    .A1(\shift_storage.storage[799] ),
    .S(net658),
    .X(_04913_));
 sg13g2_and2_1 _11661_ (.A(net363),
    .B(_04913_),
    .X(_01481_));
 sg13g2_mux2_1 _11662_ (.A0(\shift_storage.storage[801] ),
    .A1(\shift_storage.storage[800] ),
    .S(net658),
    .X(_04914_));
 sg13g2_and2_1 _11663_ (.A(net363),
    .B(_04914_),
    .X(_01482_));
 sg13g2_buf_2 fanout56 (.A(_02185_),
    .X(net56));
 sg13g2_mux2_1 _11665_ (.A0(\shift_storage.storage[802] ),
    .A1(\shift_storage.storage[801] ),
    .S(net658),
    .X(_04916_));
 sg13g2_and2_1 _11666_ (.A(net363),
    .B(_04916_),
    .X(_01483_));
 sg13g2_mux2_1 _11667_ (.A0(\shift_storage.storage[803] ),
    .A1(\shift_storage.storage[802] ),
    .S(net658),
    .X(_04917_));
 sg13g2_and2_1 _11668_ (.A(net363),
    .B(_04917_),
    .X(_01484_));
 sg13g2_mux2_1 _11669_ (.A0(\shift_storage.storage[804] ),
    .A1(\shift_storage.storage[803] ),
    .S(net658),
    .X(_04918_));
 sg13g2_and2_1 _11670_ (.A(net362),
    .B(_04918_),
    .X(_01485_));
 sg13g2_buf_2 fanout55 (.A(_02250_),
    .X(net55));
 sg13g2_mux2_1 _11672_ (.A0(\shift_storage.storage[805] ),
    .A1(\shift_storage.storage[804] ),
    .S(net658),
    .X(_04920_));
 sg13g2_and2_1 _11673_ (.A(net362),
    .B(_04920_),
    .X(_01486_));
 sg13g2_mux2_1 _11674_ (.A0(\shift_storage.storage[806] ),
    .A1(\shift_storage.storage[805] ),
    .S(net564),
    .X(_04921_));
 sg13g2_and2_1 _11675_ (.A(net264),
    .B(_04921_),
    .X(_01487_));
 sg13g2_mux2_1 _11676_ (.A0(\shift_storage.storage[807] ),
    .A1(\shift_storage.storage[806] ),
    .S(net564),
    .X(_04922_));
 sg13g2_and2_1 _11677_ (.A(net264),
    .B(_04922_),
    .X(_01488_));
 sg13g2_mux2_1 _11678_ (.A0(\shift_storage.storage[808] ),
    .A1(\shift_storage.storage[807] ),
    .S(net564),
    .X(_04923_));
 sg13g2_and2_1 _11679_ (.A(net264),
    .B(_04923_),
    .X(_01489_));
 sg13g2_mux2_1 _11680_ (.A0(\shift_storage.storage[809] ),
    .A1(\shift_storage.storage[808] ),
    .S(net564),
    .X(_04924_));
 sg13g2_and2_1 _11681_ (.A(net264),
    .B(_04924_),
    .X(_01490_));
 sg13g2_mux2_1 _11682_ (.A0(\shift_storage.storage[80] ),
    .A1(\shift_storage.storage[79] ),
    .S(net642),
    .X(_04925_));
 sg13g2_and2_1 _11683_ (.A(net345),
    .B(_04925_),
    .X(_01491_));
 sg13g2_mux2_1 _11684_ (.A0(\shift_storage.storage[810] ),
    .A1(\shift_storage.storage[809] ),
    .S(net564),
    .X(_04926_));
 sg13g2_and2_1 _11685_ (.A(net264),
    .B(_04926_),
    .X(_01492_));
 sg13g2_buf_2 fanout54 (.A(_02375_),
    .X(net54));
 sg13g2_mux2_1 _11687_ (.A0(\shift_storage.storage[811] ),
    .A1(\shift_storage.storage[810] ),
    .S(net564),
    .X(_04928_));
 sg13g2_and2_1 _11688_ (.A(net264),
    .B(_04928_),
    .X(_01493_));
 sg13g2_mux2_1 _11689_ (.A0(\shift_storage.storage[812] ),
    .A1(\shift_storage.storage[811] ),
    .S(net564),
    .X(_04929_));
 sg13g2_and2_1 _11690_ (.A(net264),
    .B(_04929_),
    .X(_01494_));
 sg13g2_mux2_1 _11691_ (.A0(\shift_storage.storage[813] ),
    .A1(\shift_storage.storage[812] ),
    .S(net564),
    .X(_04930_));
 sg13g2_and2_1 _11692_ (.A(net264),
    .B(_04930_),
    .X(_01495_));
 sg13g2_buf_2 fanout53 (.A(net54),
    .X(net53));
 sg13g2_mux2_1 _11694_ (.A0(\shift_storage.storage[814] ),
    .A1(\shift_storage.storage[813] ),
    .S(net566),
    .X(_04932_));
 sg13g2_and2_1 _11695_ (.A(net266),
    .B(_04932_),
    .X(_01496_));
 sg13g2_mux2_1 _11696_ (.A0(\shift_storage.storage[815] ),
    .A1(\shift_storage.storage[814] ),
    .S(net566),
    .X(_04933_));
 sg13g2_and2_1 _11697_ (.A(net266),
    .B(_04933_),
    .X(_01497_));
 sg13g2_mux2_1 _11698_ (.A0(\shift_storage.storage[816] ),
    .A1(\shift_storage.storage[815] ),
    .S(net658),
    .X(_04934_));
 sg13g2_and2_1 _11699_ (.A(net362),
    .B(_04934_),
    .X(_01498_));
 sg13g2_mux2_1 _11700_ (.A0(\shift_storage.storage[817] ),
    .A1(\shift_storage.storage[816] ),
    .S(net658),
    .X(_04935_));
 sg13g2_and2_1 _11701_ (.A(net362),
    .B(_04935_),
    .X(_01499_));
 sg13g2_mux2_1 _11702_ (.A0(\shift_storage.storage[818] ),
    .A1(\shift_storage.storage[817] ),
    .S(net672),
    .X(_04936_));
 sg13g2_and2_1 _11703_ (.A(net377),
    .B(_04936_),
    .X(_01500_));
 sg13g2_mux2_1 _11704_ (.A0(\shift_storage.storage[819] ),
    .A1(\shift_storage.storage[818] ),
    .S(net672),
    .X(_04937_));
 sg13g2_and2_1 _11705_ (.A(net377),
    .B(_04937_),
    .X(_01501_));
 sg13g2_mux2_1 _11706_ (.A0(\shift_storage.storage[81] ),
    .A1(\shift_storage.storage[80] ),
    .S(net642),
    .X(_04938_));
 sg13g2_and2_1 _11707_ (.A(net345),
    .B(_04938_),
    .X(_01502_));
 sg13g2_buf_1 fanout52 (.A(_03041_),
    .X(net52));
 sg13g2_buf_2 fanout51 (.A(_03041_),
    .X(net51));
 sg13g2_mux2_1 _11710_ (.A0(\shift_storage.storage[820] ),
    .A1(\shift_storage.storage[819] ),
    .S(net672),
    .X(_04941_));
 sg13g2_and2_1 _11711_ (.A(net377),
    .B(_04941_),
    .X(_01503_));
 sg13g2_mux2_1 _11712_ (.A0(\shift_storage.storage[821] ),
    .A1(\shift_storage.storage[820] ),
    .S(net672),
    .X(_04942_));
 sg13g2_and2_1 _11713_ (.A(net377),
    .B(_04942_),
    .X(_01504_));
 sg13g2_mux2_1 _11714_ (.A0(\shift_storage.storage[822] ),
    .A1(\shift_storage.storage[821] ),
    .S(net672),
    .X(_04943_));
 sg13g2_and2_1 _11715_ (.A(net378),
    .B(_04943_),
    .X(_01505_));
 sg13g2_buf_1 fanout50 (.A(_03046_),
    .X(net50));
 sg13g2_buf_2 fanout49 (.A(_03046_),
    .X(net49));
 sg13g2_mux2_1 _11718_ (.A0(\shift_storage.storage[823] ),
    .A1(\shift_storage.storage[822] ),
    .S(net673),
    .X(_04946_));
 sg13g2_and2_1 _11719_ (.A(net377),
    .B(_04946_),
    .X(_01506_));
 sg13g2_mux2_1 _11720_ (.A0(\shift_storage.storage[824] ),
    .A1(\shift_storage.storage[823] ),
    .S(net673),
    .X(_04947_));
 sg13g2_and2_1 _11721_ (.A(net377),
    .B(_04947_),
    .X(_01507_));
 sg13g2_mux2_1 _11722_ (.A0(\shift_storage.storage[825] ),
    .A1(\shift_storage.storage[824] ),
    .S(net672),
    .X(_04948_));
 sg13g2_and2_1 _11723_ (.A(net378),
    .B(_04948_),
    .X(_01508_));
 sg13g2_mux2_1 _11724_ (.A0(\shift_storage.storage[826] ),
    .A1(\shift_storage.storage[825] ),
    .S(net672),
    .X(_04949_));
 sg13g2_and2_1 _11725_ (.A(net377),
    .B(_04949_),
    .X(_01509_));
 sg13g2_mux2_1 _11726_ (.A0(\shift_storage.storage[827] ),
    .A1(\shift_storage.storage[826] ),
    .S(net672),
    .X(_04950_));
 sg13g2_and2_1 _11727_ (.A(net377),
    .B(_04950_),
    .X(_01510_));
 sg13g2_mux2_1 _11728_ (.A0(\shift_storage.storage[828] ),
    .A1(\shift_storage.storage[827] ),
    .S(net674),
    .X(_04951_));
 sg13g2_and2_1 _11729_ (.A(net379),
    .B(_04951_),
    .X(_01511_));
 sg13g2_mux2_1 _11730_ (.A0(\shift_storage.storage[829] ),
    .A1(\shift_storage.storage[828] ),
    .S(net674),
    .X(_04952_));
 sg13g2_and2_1 _11731_ (.A(net379),
    .B(_04952_),
    .X(_01512_));
 sg13g2_buf_2 fanout48 (.A(_03075_),
    .X(net48));
 sg13g2_mux2_1 _11733_ (.A0(\shift_storage.storage[82] ),
    .A1(\shift_storage.storage[81] ),
    .S(net628),
    .X(_04954_));
 sg13g2_and2_1 _11734_ (.A(net330),
    .B(_04954_),
    .X(_01513_));
 sg13g2_mux2_1 _11735_ (.A0(\shift_storage.storage[830] ),
    .A1(\shift_storage.storage[829] ),
    .S(net674),
    .X(_04955_));
 sg13g2_and2_1 _11736_ (.A(net379),
    .B(_04955_),
    .X(_01514_));
 sg13g2_mux2_1 _11737_ (.A0(\shift_storage.storage[831] ),
    .A1(\shift_storage.storage[830] ),
    .S(net674),
    .X(_04956_));
 sg13g2_and2_1 _11738_ (.A(net379),
    .B(_04956_),
    .X(_01515_));
 sg13g2_buf_1 fanout47 (.A(net48),
    .X(net47));
 sg13g2_mux2_1 _11740_ (.A0(\shift_storage.storage[832] ),
    .A1(\shift_storage.storage[831] ),
    .S(net674),
    .X(_04958_));
 sg13g2_and2_1 _11741_ (.A(net379),
    .B(_04958_),
    .X(_01516_));
 sg13g2_mux2_1 _11742_ (.A0(\shift_storage.storage[833] ),
    .A1(\shift_storage.storage[832] ),
    .S(net674),
    .X(_04959_));
 sg13g2_and2_1 _11743_ (.A(net380),
    .B(_04959_),
    .X(_01517_));
 sg13g2_mux2_1 _11744_ (.A0(\shift_storage.storage[834] ),
    .A1(\shift_storage.storage[833] ),
    .S(net682),
    .X(_04960_));
 sg13g2_and2_1 _11745_ (.A(net387),
    .B(_04960_),
    .X(_01518_));
 sg13g2_mux2_1 _11746_ (.A0(\shift_storage.storage[835] ),
    .A1(\shift_storage.storage[834] ),
    .S(net682),
    .X(_04961_));
 sg13g2_and2_1 _11747_ (.A(net387),
    .B(_04961_),
    .X(_01519_));
 sg13g2_mux2_1 _11748_ (.A0(\shift_storage.storage[836] ),
    .A1(\shift_storage.storage[835] ),
    .S(net682),
    .X(_04962_));
 sg13g2_and2_1 _11749_ (.A(net387),
    .B(_04962_),
    .X(_01520_));
 sg13g2_mux2_1 _11750_ (.A0(\shift_storage.storage[837] ),
    .A1(\shift_storage.storage[836] ),
    .S(net682),
    .X(_04963_));
 sg13g2_and2_1 _11751_ (.A(net387),
    .B(_04963_),
    .X(_01521_));
 sg13g2_mux2_1 _11752_ (.A0(\shift_storage.storage[838] ),
    .A1(\shift_storage.storage[837] ),
    .S(net668),
    .X(_04964_));
 sg13g2_and2_1 _11753_ (.A(net372),
    .B(_04964_),
    .X(_01522_));
 sg13g2_buf_2 fanout46 (.A(net48),
    .X(net46));
 sg13g2_mux2_1 _11755_ (.A0(\shift_storage.storage[839] ),
    .A1(\shift_storage.storage[838] ),
    .S(net671),
    .X(_04966_));
 sg13g2_and2_1 _11756_ (.A(net372),
    .B(_04966_),
    .X(_01523_));
 sg13g2_mux2_1 _11757_ (.A0(\shift_storage.storage[83] ),
    .A1(\shift_storage.storage[82] ),
    .S(net628),
    .X(_04967_));
 sg13g2_and2_1 _11758_ (.A(net330),
    .B(_04967_),
    .X(_01524_));
 sg13g2_mux2_1 _11759_ (.A0(\shift_storage.storage[840] ),
    .A1(\shift_storage.storage[839] ),
    .S(net668),
    .X(_04968_));
 sg13g2_and2_1 _11760_ (.A(net372),
    .B(_04968_),
    .X(_01525_));
 sg13g2_buf_1 fanout45 (.A(_03099_),
    .X(net45));
 sg13g2_mux2_1 _11762_ (.A0(\shift_storage.storage[841] ),
    .A1(\shift_storage.storage[840] ),
    .S(net668),
    .X(_04970_));
 sg13g2_and2_1 _11763_ (.A(net372),
    .B(_04970_),
    .X(_01526_));
 sg13g2_mux2_1 _11764_ (.A0(\shift_storage.storage[842] ),
    .A1(\shift_storage.storage[841] ),
    .S(net660),
    .X(_04971_));
 sg13g2_and2_1 _11765_ (.A(net364),
    .B(_04971_),
    .X(_01527_));
 sg13g2_mux2_1 _11766_ (.A0(\shift_storage.storage[843] ),
    .A1(\shift_storage.storage[842] ),
    .S(net660),
    .X(_04972_));
 sg13g2_and2_1 _11767_ (.A(net365),
    .B(_04972_),
    .X(_01528_));
 sg13g2_mux2_1 _11768_ (.A0(\shift_storage.storage[844] ),
    .A1(\shift_storage.storage[843] ),
    .S(net660),
    .X(_04973_));
 sg13g2_and2_1 _11769_ (.A(net365),
    .B(_04973_),
    .X(_01529_));
 sg13g2_mux2_1 _11770_ (.A0(\shift_storage.storage[845] ),
    .A1(\shift_storage.storage[844] ),
    .S(net660),
    .X(_04974_));
 sg13g2_and2_1 _11771_ (.A(net365),
    .B(_04974_),
    .X(_01530_));
 sg13g2_mux2_1 _11772_ (.A0(\shift_storage.storage[846] ),
    .A1(\shift_storage.storage[845] ),
    .S(net667),
    .X(_04975_));
 sg13g2_and2_1 _11773_ (.A(net364),
    .B(_04975_),
    .X(_01531_));
 sg13g2_mux2_1 _11774_ (.A0(\shift_storage.storage[847] ),
    .A1(\shift_storage.storage[846] ),
    .S(net667),
    .X(_04976_));
 sg13g2_and2_1 _11775_ (.A(net371),
    .B(_04976_),
    .X(_01532_));
 sg13g2_buf_2 fanout44 (.A(_03099_),
    .X(net44));
 sg13g2_mux2_1 _11777_ (.A0(\shift_storage.storage[848] ),
    .A1(\shift_storage.storage[847] ),
    .S(net667),
    .X(_04978_));
 sg13g2_and2_1 _11778_ (.A(net372),
    .B(_04978_),
    .X(_01533_));
 sg13g2_mux2_1 _11779_ (.A0(\shift_storage.storage[849] ),
    .A1(\shift_storage.storage[848] ),
    .S(net671),
    .X(_04979_));
 sg13g2_and2_1 _11780_ (.A(net375),
    .B(_04979_),
    .X(_01534_));
 sg13g2_mux2_1 _11781_ (.A0(\shift_storage.storage[84] ),
    .A1(\shift_storage.storage[83] ),
    .S(net642),
    .X(_04980_));
 sg13g2_and2_1 _11782_ (.A(net343),
    .B(_04980_),
    .X(_01535_));
 sg13g2_buf_2 fanout43 (.A(_03118_),
    .X(net43));
 sg13g2_mux2_1 _11784_ (.A0(\shift_storage.storage[850] ),
    .A1(\shift_storage.storage[849] ),
    .S(net668),
    .X(_04982_));
 sg13g2_and2_1 _11785_ (.A(net371),
    .B(_04982_),
    .X(_01536_));
 sg13g2_mux2_1 _11786_ (.A0(\shift_storage.storage[851] ),
    .A1(\shift_storage.storage[850] ),
    .S(net668),
    .X(_04983_));
 sg13g2_and2_1 _11787_ (.A(net371),
    .B(_04983_),
    .X(_01537_));
 sg13g2_mux2_1 _11788_ (.A0(\shift_storage.storage[852] ),
    .A1(\shift_storage.storage[851] ),
    .S(net669),
    .X(_04984_));
 sg13g2_and2_1 _11789_ (.A(net373),
    .B(_04984_),
    .X(_01538_));
 sg13g2_mux2_1 _11790_ (.A0(\shift_storage.storage[853] ),
    .A1(\shift_storage.storage[852] ),
    .S(net669),
    .X(_04985_));
 sg13g2_and2_1 _11791_ (.A(net373),
    .B(_04985_),
    .X(_01539_));
 sg13g2_mux2_1 _11792_ (.A0(\shift_storage.storage[854] ),
    .A1(\shift_storage.storage[853] ),
    .S(net669),
    .X(_04986_));
 sg13g2_and2_1 _11793_ (.A(net373),
    .B(_04986_),
    .X(_01540_));
 sg13g2_mux2_1 _11794_ (.A0(\shift_storage.storage[855] ),
    .A1(\shift_storage.storage[854] ),
    .S(net669),
    .X(_04987_));
 sg13g2_and2_1 _11795_ (.A(net373),
    .B(_04987_),
    .X(_01541_));
 sg13g2_mux2_1 _11796_ (.A0(\shift_storage.storage[856] ),
    .A1(\shift_storage.storage[855] ),
    .S(net669),
    .X(_04988_));
 sg13g2_and2_1 _11797_ (.A(net373),
    .B(_04988_),
    .X(_01542_));
 sg13g2_buf_2 fanout42 (.A(net43),
    .X(net42));
 sg13g2_mux2_1 _11799_ (.A0(\shift_storage.storage[857] ),
    .A1(\shift_storage.storage[856] ),
    .S(net669),
    .X(_04990_));
 sg13g2_and2_1 _11800_ (.A(net373),
    .B(_04990_),
    .X(_01543_));
 sg13g2_mux2_1 _11801_ (.A0(\shift_storage.storage[858] ),
    .A1(\shift_storage.storage[857] ),
    .S(net696),
    .X(_04991_));
 sg13g2_and2_1 _11802_ (.A(net401),
    .B(_04991_),
    .X(_01544_));
 sg13g2_mux2_1 _11803_ (.A0(\shift_storage.storage[859] ),
    .A1(\shift_storage.storage[858] ),
    .S(net696),
    .X(_04992_));
 sg13g2_and2_1 _11804_ (.A(net401),
    .B(_04992_),
    .X(_01545_));
 sg13g2_buf_2 fanout41 (.A(_03137_),
    .X(net41));
 sg13g2_mux2_1 _11806_ (.A0(\shift_storage.storage[85] ),
    .A1(\shift_storage.storage[84] ),
    .S(net641),
    .X(_04994_));
 sg13g2_and2_1 _11807_ (.A(net343),
    .B(_04994_),
    .X(_01546_));
 sg13g2_mux2_1 _11808_ (.A0(\shift_storage.storage[860] ),
    .A1(\shift_storage.storage[859] ),
    .S(net696),
    .X(_04995_));
 sg13g2_and2_1 _11809_ (.A(net401),
    .B(_04995_),
    .X(_01547_));
 sg13g2_mux2_1 _11810_ (.A0(\shift_storage.storage[861] ),
    .A1(\shift_storage.storage[860] ),
    .S(net696),
    .X(_04996_));
 sg13g2_and2_1 _11811_ (.A(net401),
    .B(_04996_),
    .X(_01548_));
 sg13g2_mux2_1 _11812_ (.A0(\shift_storage.storage[862] ),
    .A1(\shift_storage.storage[861] ),
    .S(net696),
    .X(_04997_));
 sg13g2_and2_1 _11813_ (.A(net402),
    .B(_04997_),
    .X(_01549_));
 sg13g2_mux2_1 _11814_ (.A0(\shift_storage.storage[863] ),
    .A1(\shift_storage.storage[862] ),
    .S(net697),
    .X(_04998_));
 sg13g2_and2_1 _11815_ (.A(net402),
    .B(_04998_),
    .X(_01550_));
 sg13g2_mux2_1 _11816_ (.A0(\shift_storage.storage[864] ),
    .A1(\shift_storage.storage[863] ),
    .S(net700),
    .X(_04999_));
 sg13g2_and2_1 _11817_ (.A(net404),
    .B(_04999_),
    .X(_01551_));
 sg13g2_mux2_1 _11818_ (.A0(\shift_storage.storage[865] ),
    .A1(\shift_storage.storage[864] ),
    .S(net698),
    .X(_05000_));
 sg13g2_and2_1 _11819_ (.A(net403),
    .B(_05000_),
    .X(_01552_));
 sg13g2_buf_2 fanout40 (.A(_03137_),
    .X(net40));
 sg13g2_mux2_1 _11821_ (.A0(\shift_storage.storage[866] ),
    .A1(\shift_storage.storage[865] ),
    .S(net698),
    .X(_05002_));
 sg13g2_and2_1 _11822_ (.A(net403),
    .B(_05002_),
    .X(_01553_));
 sg13g2_mux2_1 _11823_ (.A0(\shift_storage.storage[867] ),
    .A1(\shift_storage.storage[866] ),
    .S(net698),
    .X(_05003_));
 sg13g2_and2_1 _11824_ (.A(net403),
    .B(_05003_),
    .X(_01554_));
 sg13g2_mux2_1 _11825_ (.A0(\shift_storage.storage[868] ),
    .A1(\shift_storage.storage[867] ),
    .S(net697),
    .X(_05004_));
 sg13g2_and2_1 _11826_ (.A(net402),
    .B(_05004_),
    .X(_01555_));
 sg13g2_buf_2 fanout39 (.A(_03157_),
    .X(net39));
 sg13g2_mux2_1 _11828_ (.A0(\shift_storage.storage[869] ),
    .A1(\shift_storage.storage[868] ),
    .S(net695),
    .X(_05006_));
 sg13g2_and2_1 _11829_ (.A(net400),
    .B(_05006_),
    .X(_01556_));
 sg13g2_mux2_1 _11830_ (.A0(\shift_storage.storage[86] ),
    .A1(\shift_storage.storage[85] ),
    .S(net641),
    .X(_05007_));
 sg13g2_and2_1 _11831_ (.A(net343),
    .B(_05007_),
    .X(_01557_));
 sg13g2_mux2_1 _11832_ (.A0(\shift_storage.storage[870] ),
    .A1(\shift_storage.storage[869] ),
    .S(net695),
    .X(_05008_));
 sg13g2_and2_1 _11833_ (.A(net400),
    .B(_05008_),
    .X(_01558_));
 sg13g2_mux2_1 _11834_ (.A0(\shift_storage.storage[871] ),
    .A1(\shift_storage.storage[870] ),
    .S(net695),
    .X(_05009_));
 sg13g2_and2_1 _11835_ (.A(net400),
    .B(_05009_),
    .X(_01559_));
 sg13g2_mux2_1 _11836_ (.A0(\shift_storage.storage[872] ),
    .A1(\shift_storage.storage[871] ),
    .S(net695),
    .X(_05010_));
 sg13g2_and2_1 _11837_ (.A(net400),
    .B(_05010_),
    .X(_01560_));
 sg13g2_mux2_1 _11838_ (.A0(\shift_storage.storage[873] ),
    .A1(\shift_storage.storage[872] ),
    .S(net695),
    .X(_05011_));
 sg13g2_and2_1 _11839_ (.A(net400),
    .B(_05011_),
    .X(_01561_));
 sg13g2_mux2_1 _11840_ (.A0(\shift_storage.storage[874] ),
    .A1(\shift_storage.storage[873] ),
    .S(net695),
    .X(_05012_));
 sg13g2_and2_1 _11841_ (.A(net400),
    .B(_05012_),
    .X(_01562_));
 sg13g2_buf_2 fanout38 (.A(_03157_),
    .X(net38));
 sg13g2_mux2_1 _11843_ (.A0(\shift_storage.storage[875] ),
    .A1(\shift_storage.storage[874] ),
    .S(net665),
    .X(_05014_));
 sg13g2_and2_1 _11844_ (.A(net370),
    .B(_05014_),
    .X(_01563_));
 sg13g2_mux2_1 _11845_ (.A0(\shift_storage.storage[876] ),
    .A1(\shift_storage.storage[875] ),
    .S(net664),
    .X(_05015_));
 sg13g2_and2_1 _11846_ (.A(net369),
    .B(_05015_),
    .X(_01564_));
 sg13g2_mux2_1 _11847_ (.A0(\shift_storage.storage[877] ),
    .A1(\shift_storage.storage[876] ),
    .S(net664),
    .X(_05016_));
 sg13g2_and2_1 _11848_ (.A(net369),
    .B(_05016_),
    .X(_01565_));
 sg13g2_buf_1 fanout37 (.A(_03178_),
    .X(net37));
 sg13g2_mux2_1 _11850_ (.A0(\shift_storage.storage[878] ),
    .A1(\shift_storage.storage[877] ),
    .S(net665),
    .X(_05018_));
 sg13g2_and2_1 _11851_ (.A(net370),
    .B(_05018_),
    .X(_01566_));
 sg13g2_mux2_1 _11852_ (.A0(\shift_storage.storage[879] ),
    .A1(\shift_storage.storage[878] ),
    .S(net665),
    .X(_05019_));
 sg13g2_and2_1 _11853_ (.A(net370),
    .B(_05019_),
    .X(_01567_));
 sg13g2_mux2_1 _11854_ (.A0(\shift_storage.storage[87] ),
    .A1(\shift_storage.storage[86] ),
    .S(net641),
    .X(_05020_));
 sg13g2_and2_1 _11855_ (.A(net343),
    .B(_05020_),
    .X(_01568_));
 sg13g2_mux2_1 _11856_ (.A0(\shift_storage.storage[880] ),
    .A1(\shift_storage.storage[879] ),
    .S(net665),
    .X(_05021_));
 sg13g2_and2_1 _11857_ (.A(net370),
    .B(_05021_),
    .X(_01569_));
 sg13g2_mux2_1 _11858_ (.A0(\shift_storage.storage[881] ),
    .A1(\shift_storage.storage[880] ),
    .S(net665),
    .X(_05022_));
 sg13g2_and2_1 _11859_ (.A(net370),
    .B(_05022_),
    .X(_01570_));
 sg13g2_mux2_1 _11860_ (.A0(\shift_storage.storage[882] ),
    .A1(\shift_storage.storage[881] ),
    .S(net665),
    .X(_05023_));
 sg13g2_and2_1 _11861_ (.A(net370),
    .B(_05023_),
    .X(_01571_));
 sg13g2_mux2_1 _11862_ (.A0(\shift_storage.storage[883] ),
    .A1(\shift_storage.storage[882] ),
    .S(net663),
    .X(_05024_));
 sg13g2_and2_1 _11863_ (.A(net368),
    .B(_05024_),
    .X(_01572_));
 sg13g2_buf_2 fanout36 (.A(_03178_),
    .X(net36));
 sg13g2_buf_2 fanout35 (.A(_02544_),
    .X(net35));
 sg13g2_mux2_1 _11866_ (.A0(\shift_storage.storage[884] ),
    .A1(\shift_storage.storage[883] ),
    .S(net663),
    .X(_05027_));
 sg13g2_and2_1 _11867_ (.A(net368),
    .B(_05027_),
    .X(_01573_));
 sg13g2_mux2_1 _11868_ (.A0(\shift_storage.storage[885] ),
    .A1(\shift_storage.storage[884] ),
    .S(net663),
    .X(_05028_));
 sg13g2_and2_1 _11869_ (.A(net367),
    .B(_05028_),
    .X(_01574_));
 sg13g2_mux2_1 _11870_ (.A0(\shift_storage.storage[886] ),
    .A1(\shift_storage.storage[885] ),
    .S(net663),
    .X(_05029_));
 sg13g2_and2_1 _11871_ (.A(net367),
    .B(_05029_),
    .X(_01575_));
 sg13g2_buf_8 wire34 (.A(net34),
    .X(net4050));
 sg13g2_buf_8 wire33 (.A(net33),
    .X(net4049));
 sg13g2_mux2_1 _11874_ (.A0(\shift_storage.storage[887] ),
    .A1(\shift_storage.storage[886] ),
    .S(net664),
    .X(_05032_));
 sg13g2_and2_1 _11875_ (.A(net369),
    .B(_05032_),
    .X(_01576_));
 sg13g2_mux2_1 _11876_ (.A0(\shift_storage.storage[888] ),
    .A1(\shift_storage.storage[887] ),
    .S(net664),
    .X(_05033_));
 sg13g2_and2_1 _11877_ (.A(net369),
    .B(_05033_),
    .X(_01577_));
 sg13g2_mux2_1 _11878_ (.A0(\shift_storage.storage[889] ),
    .A1(\shift_storage.storage[888] ),
    .S(net664),
    .X(_05034_));
 sg13g2_and2_1 _11879_ (.A(net369),
    .B(_05034_),
    .X(_01578_));
 sg13g2_mux2_1 _11880_ (.A0(\shift_storage.storage[88] ),
    .A1(\shift_storage.storage[87] ),
    .S(net626),
    .X(_05035_));
 sg13g2_and2_1 _11881_ (.A(net328),
    .B(_05035_),
    .X(_01579_));
 sg13g2_mux2_1 _11882_ (.A0(\shift_storage.storage[890] ),
    .A1(\shift_storage.storage[889] ),
    .S(net664),
    .X(_05036_));
 sg13g2_and2_1 _11883_ (.A(net369),
    .B(_05036_),
    .X(_01580_));
 sg13g2_mux2_1 _11884_ (.A0(\shift_storage.storage[891] ),
    .A1(\shift_storage.storage[890] ),
    .S(net664),
    .X(_05037_));
 sg13g2_and2_1 _11885_ (.A(net369),
    .B(_05037_),
    .X(_01581_));
 sg13g2_mux2_1 _11886_ (.A0(\shift_storage.storage[892] ),
    .A1(\shift_storage.storage[891] ),
    .S(net665),
    .X(_05038_));
 sg13g2_and2_1 _11887_ (.A(net370),
    .B(_05038_),
    .X(_01582_));
 sg13g2_buf_2 fanout32 (.A(_01761_),
    .X(net32));
 sg13g2_mux2_1 _11889_ (.A0(\shift_storage.storage[893] ),
    .A1(\shift_storage.storage[892] ),
    .S(net664),
    .X(_05040_));
 sg13g2_and2_1 _11890_ (.A(net369),
    .B(_05040_),
    .X(_01583_));
 sg13g2_mux2_1 _11891_ (.A0(\shift_storage.storage[894] ),
    .A1(\shift_storage.storage[893] ),
    .S(net696),
    .X(_05041_));
 sg13g2_and2_1 _11892_ (.A(net401),
    .B(_05041_),
    .X(_01584_));
 sg13g2_mux2_1 _11893_ (.A0(\shift_storage.storage[895] ),
    .A1(\shift_storage.storage[894] ),
    .S(net696),
    .X(_05042_));
 sg13g2_and2_1 _11894_ (.A(net401),
    .B(_05042_),
    .X(_01585_));
 sg13g2_buf_2 fanout31 (.A(_01861_),
    .X(net31));
 sg13g2_mux2_1 _11896_ (.A0(\shift_storage.storage[896] ),
    .A1(\shift_storage.storage[895] ),
    .S(net696),
    .X(_05044_));
 sg13g2_and2_1 _11897_ (.A(net401),
    .B(_05044_),
    .X(_01586_));
 sg13g2_mux2_1 _11898_ (.A0(\shift_storage.storage[897] ),
    .A1(\shift_storage.storage[896] ),
    .S(net697),
    .X(_05045_));
 sg13g2_and2_1 _11899_ (.A(net401),
    .B(_05045_),
    .X(_01587_));
 sg13g2_mux2_1 _11900_ (.A0(\shift_storage.storage[898] ),
    .A1(\shift_storage.storage[897] ),
    .S(net697),
    .X(_05046_));
 sg13g2_and2_1 _11901_ (.A(net402),
    .B(_05046_),
    .X(_01588_));
 sg13g2_mux2_1 _11902_ (.A0(\shift_storage.storage[899] ),
    .A1(\shift_storage.storage[898] ),
    .S(net698),
    .X(_05047_));
 sg13g2_and2_1 _11903_ (.A(net403),
    .B(_05047_),
    .X(_01589_));
 sg13g2_mux2_1 _11904_ (.A0(\shift_storage.storage[89] ),
    .A1(\shift_storage.storage[88] ),
    .S(net626),
    .X(_05048_));
 sg13g2_and2_1 _11905_ (.A(net328),
    .B(_05048_),
    .X(_01590_));
 sg13g2_mux2_1 _11906_ (.A0(\shift_storage.storage[8] ),
    .A1(\shift_storage.storage[7] ),
    .S(net608),
    .X(_05049_));
 sg13g2_and2_1 _11907_ (.A(net310),
    .B(_05049_),
    .X(_01591_));
 sg13g2_mux2_1 _11908_ (.A0(\shift_storage.storage[900] ),
    .A1(\shift_storage.storage[899] ),
    .S(net698),
    .X(_05050_));
 sg13g2_and2_1 _11909_ (.A(net403),
    .B(_05050_),
    .X(_01592_));
 sg13g2_buf_2 fanout30 (.A(_01913_),
    .X(net30));
 sg13g2_mux2_1 _11911_ (.A0(\shift_storage.storage[901] ),
    .A1(\shift_storage.storage[900] ),
    .S(net698),
    .X(_05052_));
 sg13g2_and2_1 _11912_ (.A(net403),
    .B(_05052_),
    .X(_01593_));
 sg13g2_mux2_1 _11913_ (.A0(\shift_storage.storage[902] ),
    .A1(\shift_storage.storage[901] ),
    .S(net694),
    .X(_05053_));
 sg13g2_and2_1 _11914_ (.A(net399),
    .B(_05053_),
    .X(_01594_));
 sg13g2_mux2_1 _11915_ (.A0(\shift_storage.storage[903] ),
    .A1(\shift_storage.storage[902] ),
    .S(net694),
    .X(_05054_));
 sg13g2_and2_1 _11916_ (.A(net399),
    .B(_05054_),
    .X(_01595_));
 sg13g2_buf_2 fanout29 (.A(_01913_),
    .X(net29));
 sg13g2_mux2_1 _11918_ (.A0(\shift_storage.storage[904] ),
    .A1(\shift_storage.storage[903] ),
    .S(net694),
    .X(_05056_));
 sg13g2_and2_1 _11919_ (.A(net399),
    .B(_05056_),
    .X(_01596_));
 sg13g2_mux2_1 _11920_ (.A0(\shift_storage.storage[905] ),
    .A1(\shift_storage.storage[904] ),
    .S(net694),
    .X(_05057_));
 sg13g2_and2_1 _11921_ (.A(net399),
    .B(_05057_),
    .X(_01597_));
 sg13g2_mux2_1 _11922_ (.A0(\shift_storage.storage[906] ),
    .A1(\shift_storage.storage[905] ),
    .S(net694),
    .X(_05058_));
 sg13g2_and2_1 _11923_ (.A(net399),
    .B(_05058_),
    .X(_01598_));
 sg13g2_mux2_1 _11924_ (.A0(\shift_storage.storage[907] ),
    .A1(\shift_storage.storage[906] ),
    .S(net694),
    .X(_05059_));
 sg13g2_and2_1 _11925_ (.A(net399),
    .B(_05059_),
    .X(_01599_));
 sg13g2_mux2_1 _11926_ (.A0(\shift_storage.storage[908] ),
    .A1(\shift_storage.storage[907] ),
    .S(net695),
    .X(_05060_));
 sg13g2_and2_1 _11927_ (.A(net400),
    .B(_05060_),
    .X(_01600_));
 sg13g2_mux2_1 _11928_ (.A0(\shift_storage.storage[909] ),
    .A1(\shift_storage.storage[908] ),
    .S(net712),
    .X(_05061_));
 sg13g2_and2_1 _11929_ (.A(net418),
    .B(_05061_),
    .X(_01601_));
 sg13g2_mux2_1 _11930_ (.A0(\shift_storage.storage[90] ),
    .A1(\shift_storage.storage[89] ),
    .S(net626),
    .X(_05062_));
 sg13g2_and2_1 _11931_ (.A(net328),
    .B(_05062_),
    .X(_01602_));
 sg13g2_buf_1 fanout28 (.A(_01963_),
    .X(net28));
 sg13g2_mux2_1 _11933_ (.A0(\shift_storage.storage[910] ),
    .A1(\shift_storage.storage[909] ),
    .S(net694),
    .X(_05064_));
 sg13g2_and2_1 _11934_ (.A(net399),
    .B(_05064_),
    .X(_01603_));
 sg13g2_mux2_1 _11935_ (.A0(\shift_storage.storage[911] ),
    .A1(\shift_storage.storage[910] ),
    .S(net694),
    .X(_05065_));
 sg13g2_and2_1 _11936_ (.A(net399),
    .B(_05065_),
    .X(_01604_));
 sg13g2_mux2_1 _11937_ (.A0(\shift_storage.storage[912] ),
    .A1(\shift_storage.storage[911] ),
    .S(net701),
    .X(_05066_));
 sg13g2_and2_1 _11938_ (.A(net406),
    .B(_05066_),
    .X(_01605_));
 sg13g2_buf_2 fanout27 (.A(_01963_),
    .X(net27));
 sg13g2_mux2_1 _11940_ (.A0(\shift_storage.storage[913] ),
    .A1(\shift_storage.storage[912] ),
    .S(net701),
    .X(_05068_));
 sg13g2_and2_1 _11941_ (.A(net406),
    .B(_05068_),
    .X(_01606_));
 sg13g2_mux2_1 _11942_ (.A0(\shift_storage.storage[914] ),
    .A1(\shift_storage.storage[913] ),
    .S(net701),
    .X(_05069_));
 sg13g2_and2_1 _11943_ (.A(net406),
    .B(_05069_),
    .X(_01607_));
 sg13g2_mux2_1 _11944_ (.A0(\shift_storage.storage[915] ),
    .A1(\shift_storage.storage[914] ),
    .S(net701),
    .X(_05070_));
 sg13g2_and2_1 _11945_ (.A(net407),
    .B(_05070_),
    .X(_01608_));
 sg13g2_mux2_1 _11946_ (.A0(\shift_storage.storage[916] ),
    .A1(\shift_storage.storage[915] ),
    .S(net701),
    .X(_05071_));
 sg13g2_and2_1 _11947_ (.A(net406),
    .B(_05071_),
    .X(_01609_));
 sg13g2_mux2_1 _11948_ (.A0(\shift_storage.storage[917] ),
    .A1(\shift_storage.storage[916] ),
    .S(net702),
    .X(_05072_));
 sg13g2_and2_1 _11949_ (.A(net406),
    .B(_05072_),
    .X(_01610_));
 sg13g2_mux2_1 _11950_ (.A0(\shift_storage.storage[918] ),
    .A1(\shift_storage.storage[917] ),
    .S(net702),
    .X(_05073_));
 sg13g2_and2_1 _11951_ (.A(net406),
    .B(_05073_),
    .X(_01611_));
 sg13g2_mux2_1 _11952_ (.A0(\shift_storage.storage[919] ),
    .A1(\shift_storage.storage[918] ),
    .S(net701),
    .X(_05074_));
 sg13g2_and2_1 _11953_ (.A(net407),
    .B(_05074_),
    .X(_01612_));
 sg13g2_buf_1 fanout26 (.A(_02022_),
    .X(net26));
 sg13g2_mux2_1 _11955_ (.A0(\shift_storage.storage[91] ),
    .A1(\shift_storage.storage[90] ),
    .S(net625),
    .X(_05076_));
 sg13g2_and2_1 _11956_ (.A(net327),
    .B(_05076_),
    .X(_01613_));
 sg13g2_mux2_1 _11957_ (.A0(\shift_storage.storage[920] ),
    .A1(\shift_storage.storage[919] ),
    .S(net702),
    .X(_05077_));
 sg13g2_and2_1 _11958_ (.A(net407),
    .B(_05077_),
    .X(_01614_));
 sg13g2_mux2_1 _11959_ (.A0(\shift_storage.storage[921] ),
    .A1(\shift_storage.storage[920] ),
    .S(net704),
    .X(_05078_));
 sg13g2_and2_1 _11960_ (.A(net409),
    .B(_05078_),
    .X(_01615_));
 sg13g2_buf_2 fanout25 (.A(net26),
    .X(net25));
 sg13g2_mux2_1 _11962_ (.A0(\shift_storage.storage[922] ),
    .A1(\shift_storage.storage[921] ),
    .S(net704),
    .X(_05080_));
 sg13g2_and2_1 _11963_ (.A(net409),
    .B(_05080_),
    .X(_01616_));
 sg13g2_mux2_1 _11964_ (.A0(\shift_storage.storage[923] ),
    .A1(\shift_storage.storage[922] ),
    .S(net704),
    .X(_05081_));
 sg13g2_and2_1 _11965_ (.A(net409),
    .B(_05081_),
    .X(_01617_));
 sg13g2_mux2_1 _11966_ (.A0(\shift_storage.storage[924] ),
    .A1(\shift_storage.storage[923] ),
    .S(net704),
    .X(_05082_));
 sg13g2_and2_1 _11967_ (.A(net409),
    .B(_05082_),
    .X(_01618_));
 sg13g2_mux2_1 _11968_ (.A0(\shift_storage.storage[925] ),
    .A1(\shift_storage.storage[924] ),
    .S(net708),
    .X(_05083_));
 sg13g2_and2_1 _11969_ (.A(net413),
    .B(_05083_),
    .X(_01619_));
 sg13g2_mux2_1 _11970_ (.A0(\shift_storage.storage[926] ),
    .A1(\shift_storage.storage[925] ),
    .S(net709),
    .X(_05084_));
 sg13g2_and2_1 _11971_ (.A(net414),
    .B(_05084_),
    .X(_01620_));
 sg13g2_mux2_1 _11972_ (.A0(\shift_storage.storage[927] ),
    .A1(\shift_storage.storage[926] ),
    .S(net708),
    .X(_05085_));
 sg13g2_and2_1 _11973_ (.A(net413),
    .B(_05085_),
    .X(_01621_));
 sg13g2_mux2_1 _11974_ (.A0(\shift_storage.storage[928] ),
    .A1(\shift_storage.storage[927] ),
    .S(net709),
    .X(_05086_));
 sg13g2_and2_1 _11975_ (.A(net414),
    .B(_05086_),
    .X(_01622_));
 sg13g2_buf_2 fanout24 (.A(_02062_),
    .X(net24));
 sg13g2_mux2_1 _11977_ (.A0(\shift_storage.storage[929] ),
    .A1(\shift_storage.storage[928] ),
    .S(net704),
    .X(_05088_));
 sg13g2_and2_1 _11978_ (.A(net409),
    .B(_05088_),
    .X(_01623_));
 sg13g2_mux2_1 _11979_ (.A0(\shift_storage.storage[92] ),
    .A1(\shift_storage.storage[91] ),
    .S(net626),
    .X(_05089_));
 sg13g2_and2_1 _11980_ (.A(net328),
    .B(_05089_),
    .X(_01624_));
 sg13g2_mux2_1 _11981_ (.A0(\shift_storage.storage[930] ),
    .A1(\shift_storage.storage[929] ),
    .S(net704),
    .X(_05090_));
 sg13g2_and2_1 _11982_ (.A(net409),
    .B(_05090_),
    .X(_01625_));
 sg13g2_buf_2 fanout23 (.A(_02522_),
    .X(net23));
 sg13g2_mux2_1 _11984_ (.A0(\shift_storage.storage[931] ),
    .A1(\shift_storage.storage[930] ),
    .S(net704),
    .X(_05092_));
 sg13g2_and2_1 _11985_ (.A(net409),
    .B(_05092_),
    .X(_01626_));
 sg13g2_mux2_1 _11986_ (.A0(\shift_storage.storage[932] ),
    .A1(\shift_storage.storage[931] ),
    .S(net704),
    .X(_05093_));
 sg13g2_and2_1 _11987_ (.A(net409),
    .B(_05093_),
    .X(_01627_));
 sg13g2_mux2_1 _11988_ (.A0(\shift_storage.storage[933] ),
    .A1(\shift_storage.storage[932] ),
    .S(net705),
    .X(_05094_));
 sg13g2_and2_1 _11989_ (.A(net410),
    .B(_05094_),
    .X(_01628_));
 sg13g2_mux2_1 _11990_ (.A0(\shift_storage.storage[934] ),
    .A1(\shift_storage.storage[933] ),
    .S(net703),
    .X(_05095_));
 sg13g2_and2_1 _11991_ (.A(net410),
    .B(_05095_),
    .X(_01629_));
 sg13g2_mux2_1 _11992_ (.A0(\shift_storage.storage[935] ),
    .A1(\shift_storage.storage[934] ),
    .S(net703),
    .X(_05096_));
 sg13g2_and2_1 _11993_ (.A(net408),
    .B(_05096_),
    .X(_01630_));
 sg13g2_mux2_1 _11994_ (.A0(\shift_storage.storage[936] ),
    .A1(\shift_storage.storage[935] ),
    .S(net705),
    .X(_05097_));
 sg13g2_and2_1 _11995_ (.A(net408),
    .B(_05097_),
    .X(_01631_));
 sg13g2_mux2_1 _11996_ (.A0(\shift_storage.storage[937] ),
    .A1(\shift_storage.storage[936] ),
    .S(net703),
    .X(_05098_));
 sg13g2_and2_1 _11997_ (.A(net408),
    .B(_05098_),
    .X(_01632_));
 sg13g2_buf_2 fanout22 (.A(_02663_),
    .X(net22));
 sg13g2_mux2_1 _11999_ (.A0(\shift_storage.storage[938] ),
    .A1(\shift_storage.storage[937] ),
    .S(net705),
    .X(_05100_));
 sg13g2_and2_1 _12000_ (.A(net410),
    .B(_05100_),
    .X(_01633_));
 sg13g2_mux2_1 _12001_ (.A0(\shift_storage.storage[939] ),
    .A1(\shift_storage.storage[938] ),
    .S(net703),
    .X(_05101_));
 sg13g2_and2_1 _12002_ (.A(net408),
    .B(_05101_),
    .X(_01634_));
 sg13g2_mux2_1 _12003_ (.A0(\shift_storage.storage[93] ),
    .A1(\shift_storage.storage[92] ),
    .S(net625),
    .X(_05102_));
 sg13g2_and2_1 _12004_ (.A(net327),
    .B(_05102_),
    .X(_01635_));
 sg13g2_buf_8 wire21 (.A(net21),
    .X(net4037));
 sg13g2_mux2_1 _12006_ (.A0(\shift_storage.storage[940] ),
    .A1(\shift_storage.storage[939] ),
    .S(net703),
    .X(_05104_));
 sg13g2_and2_1 _12007_ (.A(net408),
    .B(_05104_),
    .X(_01636_));
 sg13g2_mux2_1 _12008_ (.A0(\shift_storage.storage[941] ),
    .A1(\shift_storage.storage[940] ),
    .S(net703),
    .X(_05105_));
 sg13g2_and2_1 _12009_ (.A(net408),
    .B(_05105_),
    .X(_01637_));
 sg13g2_mux2_1 _12010_ (.A0(\shift_storage.storage[942] ),
    .A1(\shift_storage.storage[941] ),
    .S(net703),
    .X(_05106_));
 sg13g2_and2_1 _12011_ (.A(net408),
    .B(_05106_),
    .X(_01638_));
 sg13g2_mux2_1 _12012_ (.A0(\shift_storage.storage[943] ),
    .A1(\shift_storage.storage[942] ),
    .S(net703),
    .X(_05107_));
 sg13g2_and2_1 _12013_ (.A(net408),
    .B(_05107_),
    .X(_01639_));
 sg13g2_mux2_1 _12014_ (.A0(\shift_storage.storage[944] ),
    .A1(\shift_storage.storage[943] ),
    .S(net701),
    .X(_05108_));
 sg13g2_and2_1 _12015_ (.A(net406),
    .B(_05108_),
    .X(_01640_));
 sg13g2_mux2_1 _12016_ (.A0(\shift_storage.storage[945] ),
    .A1(\shift_storage.storage[944] ),
    .S(net701),
    .X(_05109_));
 sg13g2_and2_1 _12017_ (.A(net406),
    .B(_05109_),
    .X(_01641_));
 sg13g2_mux2_1 _12018_ (.A0(\shift_storage.storage[946] ),
    .A1(\shift_storage.storage[945] ),
    .S(net702),
    .X(_05110_));
 sg13g2_and2_1 _12019_ (.A(net407),
    .B(_05110_),
    .X(_01642_));
 sg13g2_buf_2 fanout20 (.A(_02193_),
    .X(net20));
 sg13g2_mux2_1 _12021_ (.A0(\shift_storage.storage[947] ),
    .A1(\shift_storage.storage[946] ),
    .S(net702),
    .X(_05112_));
 sg13g2_and2_1 _12022_ (.A(net407),
    .B(_05112_),
    .X(_01643_));
 sg13g2_mux2_1 _12023_ (.A0(\shift_storage.storage[948] ),
    .A1(\shift_storage.storage[947] ),
    .S(net711),
    .X(_05113_));
 sg13g2_and2_1 _12024_ (.A(net407),
    .B(_05113_),
    .X(_01644_));
 sg13g2_mux2_1 _12025_ (.A0(\shift_storage.storage[949] ),
    .A1(\shift_storage.storage[948] ),
    .S(net702),
    .X(_05114_));
 sg13g2_and2_1 _12026_ (.A(net417),
    .B(_05114_),
    .X(_01645_));
 sg13g2_buf_2 fanout19 (.A(_02258_),
    .X(net19));
 sg13g2_mux2_1 _12028_ (.A0(\shift_storage.storage[94] ),
    .A1(\shift_storage.storage[93] ),
    .S(net625),
    .X(_05116_));
 sg13g2_and2_1 _12029_ (.A(net327),
    .B(_05116_),
    .X(_01646_));
 sg13g2_mux2_1 _12030_ (.A0(\shift_storage.storage[950] ),
    .A1(\shift_storage.storage[949] ),
    .S(net702),
    .X(_05117_));
 sg13g2_and2_1 _12031_ (.A(net407),
    .B(_05117_),
    .X(_01647_));
 sg13g2_mux2_1 _12032_ (.A0(\shift_storage.storage[951] ),
    .A1(\shift_storage.storage[950] ),
    .S(net706),
    .X(_05118_));
 sg13g2_and2_1 _12033_ (.A(net411),
    .B(_05118_),
    .X(_01648_));
 sg13g2_mux2_1 _12034_ (.A0(\shift_storage.storage[952] ),
    .A1(\shift_storage.storage[951] ),
    .S(net706),
    .X(_05119_));
 sg13g2_and2_1 _12035_ (.A(net411),
    .B(_05119_),
    .X(_01649_));
 sg13g2_mux2_1 _12036_ (.A0(\shift_storage.storage[953] ),
    .A1(\shift_storage.storage[952] ),
    .S(net706),
    .X(_05120_));
 sg13g2_and2_1 _12037_ (.A(net411),
    .B(_05120_),
    .X(_01650_));
 sg13g2_mux2_1 _12038_ (.A0(\shift_storage.storage[954] ),
    .A1(\shift_storage.storage[953] ),
    .S(net698),
    .X(_05121_));
 sg13g2_and2_1 _12039_ (.A(net404),
    .B(_05121_),
    .X(_01651_));
 sg13g2_mux2_1 _12040_ (.A0(\shift_storage.storage[955] ),
    .A1(\shift_storage.storage[954] ),
    .S(net698),
    .X(_05122_));
 sg13g2_and2_1 _12041_ (.A(net404),
    .B(_05122_),
    .X(_01652_));
 sg13g2_buf_2 fanout18 (.A(_02403_),
    .X(net18));
 sg13g2_mux2_1 _12043_ (.A0(\shift_storage.storage[956] ),
    .A1(\shift_storage.storage[955] ),
    .S(net699),
    .X(_05124_));
 sg13g2_and2_1 _12044_ (.A(net403),
    .B(_05124_),
    .X(_01653_));
 sg13g2_mux2_1 _12045_ (.A0(\shift_storage.storage[957] ),
    .A1(\shift_storage.storage[956] ),
    .S(net699),
    .X(_05125_));
 sg13g2_and2_1 _12046_ (.A(net404),
    .B(_05125_),
    .X(_01654_));
 sg13g2_mux2_1 _12047_ (.A0(\shift_storage.storage[958] ),
    .A1(\shift_storage.storage[957] ),
    .S(net699),
    .X(_05126_));
 sg13g2_and2_1 _12048_ (.A(net403),
    .B(_05126_),
    .X(_01655_));
 sg13g2_buf_2 fanout17 (.A(_02382_),
    .X(net17));
 sg13g2_mux2_1 _12050_ (.A0(\shift_storage.storage[959] ),
    .A1(\shift_storage.storage[958] ),
    .S(net699),
    .X(_05128_));
 sg13g2_and2_1 _12051_ (.A(net404),
    .B(_05128_),
    .X(_01656_));
 sg13g2_mux2_1 _12052_ (.A0(\shift_storage.storage[95] ),
    .A1(\shift_storage.storage[94] ),
    .S(net625),
    .X(_05129_));
 sg13g2_and2_1 _12053_ (.A(net327),
    .B(_05129_),
    .X(_01657_));
 sg13g2_mux2_1 _12054_ (.A0(\shift_storage.storage[960] ),
    .A1(\shift_storage.storage[959] ),
    .S(net699),
    .X(_05130_));
 sg13g2_and2_1 _12055_ (.A(net404),
    .B(_05130_),
    .X(_01658_));
 sg13g2_mux2_1 _12056_ (.A0(\shift_storage.storage[961] ),
    .A1(\shift_storage.storage[960] ),
    .S(net699),
    .X(_05131_));
 sg13g2_and2_1 _12057_ (.A(net412),
    .B(_05131_),
    .X(_01659_));
 sg13g2_mux2_1 _12058_ (.A0(\shift_storage.storage[962] ),
    .A1(\shift_storage.storage[961] ),
    .S(net699),
    .X(_05132_));
 sg13g2_and2_1 _12059_ (.A(net404),
    .B(_05132_),
    .X(_01660_));
 sg13g2_mux2_1 _12060_ (.A0(\shift_storage.storage[963] ),
    .A1(\shift_storage.storage[962] ),
    .S(net716),
    .X(_05133_));
 sg13g2_and2_1 _12061_ (.A(net423),
    .B(_05133_),
    .X(_01661_));
 sg13g2_mux2_1 _12062_ (.A0(\shift_storage.storage[964] ),
    .A1(\shift_storage.storage[963] ),
    .S(net716),
    .X(_05134_));
 sg13g2_and2_1 _12063_ (.A(net422),
    .B(_05134_),
    .X(_01662_));
 sg13g2_buf_8 wire16 (.A(net16),
    .X(net4032));
 sg13g2_mux2_1 _12065_ (.A0(\shift_storage.storage[965] ),
    .A1(\shift_storage.storage[964] ),
    .S(net723),
    .X(_05136_));
 sg13g2_and2_1 _12066_ (.A(net429),
    .B(_05136_),
    .X(_01663_));
 sg13g2_mux2_1 _12067_ (.A0(\shift_storage.storage[966] ),
    .A1(\shift_storage.storage[965] ),
    .S(net723),
    .X(_05137_));
 sg13g2_and2_1 _12068_ (.A(net429),
    .B(_05137_),
    .X(_01664_));
 sg13g2_mux2_1 _12069_ (.A0(\shift_storage.storage[967] ),
    .A1(\shift_storage.storage[966] ),
    .S(net707),
    .X(_05138_));
 sg13g2_and2_1 _12070_ (.A(net412),
    .B(_05138_),
    .X(_01665_));
 sg13g2_buf_8 wire15 (.A(net15),
    .X(net4031));
 sg13g2_mux2_1 _12072_ (.A0(\shift_storage.storage[968] ),
    .A1(\shift_storage.storage[967] ),
    .S(net707),
    .X(_05140_));
 sg13g2_and2_1 _12073_ (.A(net412),
    .B(_05140_),
    .X(_01666_));
 sg13g2_mux2_1 _12074_ (.A0(\shift_storage.storage[969] ),
    .A1(\shift_storage.storage[968] ),
    .S(net707),
    .X(_05141_));
 sg13g2_and2_1 _12075_ (.A(net412),
    .B(_05141_),
    .X(_01667_));
 sg13g2_mux2_1 _12076_ (.A0(\shift_storage.storage[96] ),
    .A1(\shift_storage.storage[95] ),
    .S(net625),
    .X(_05142_));
 sg13g2_and2_1 _12077_ (.A(net327),
    .B(_05142_),
    .X(_01668_));
 sg13g2_mux2_1 _12078_ (.A0(\shift_storage.storage[970] ),
    .A1(\shift_storage.storage[969] ),
    .S(net707),
    .X(_05143_));
 sg13g2_and2_1 _12079_ (.A(net415),
    .B(_05143_),
    .X(_01669_));
 sg13g2_mux2_1 _12080_ (.A0(\shift_storage.storage[971] ),
    .A1(\shift_storage.storage[970] ),
    .S(net707),
    .X(_05144_));
 sg13g2_and2_1 _12081_ (.A(net415),
    .B(_05144_),
    .X(_01670_));
 sg13g2_mux2_1 _12082_ (.A0(\shift_storage.storage[972] ),
    .A1(\shift_storage.storage[971] ),
    .S(net707),
    .X(_05145_));
 sg13g2_and2_1 _12083_ (.A(net412),
    .B(_05145_),
    .X(_01671_));
 sg13g2_mux2_1 _12084_ (.A0(\shift_storage.storage[973] ),
    .A1(\shift_storage.storage[972] ),
    .S(net707),
    .X(_05146_));
 sg13g2_and2_1 _12085_ (.A(net411),
    .B(_05146_),
    .X(_01672_));
 sg13g2_buf_1 fanout14 (.A(_02089_),
    .X(net14));
 sg13g2_mux2_1 _12087_ (.A0(\shift_storage.storage[974] ),
    .A1(\shift_storage.storage[973] ),
    .S(net706),
    .X(_05148_));
 sg13g2_and2_1 _12088_ (.A(net411),
    .B(_05148_),
    .X(_01673_));
 sg13g2_mux2_1 _12089_ (.A0(\shift_storage.storage[975] ),
    .A1(\shift_storage.storage[974] ),
    .S(net706),
    .X(_05149_));
 sg13g2_and2_1 _12090_ (.A(net411),
    .B(_05149_),
    .X(_01674_));
 sg13g2_mux2_1 _12091_ (.A0(\shift_storage.storage[976] ),
    .A1(\shift_storage.storage[975] ),
    .S(net706),
    .X(_05150_));
 sg13g2_and2_1 _12092_ (.A(net411),
    .B(_05150_),
    .X(_01675_));
 sg13g2_buf_1 fanout13 (.A(net14),
    .X(net13));
 sg13g2_mux2_1 _12094_ (.A0(\shift_storage.storage[977] ),
    .A1(\shift_storage.storage[976] ),
    .S(net706),
    .X(_05152_));
 sg13g2_and2_1 _12095_ (.A(net411),
    .B(_05152_),
    .X(_01676_));
 sg13g2_mux2_1 _12096_ (.A0(\shift_storage.storage[978] ),
    .A1(\shift_storage.storage[977] ),
    .S(net706),
    .X(_05153_));
 sg13g2_and2_1 _12097_ (.A(net413),
    .B(_05153_),
    .X(_01677_));
 sg13g2_mux2_1 _12098_ (.A0(\shift_storage.storage[979] ),
    .A1(\shift_storage.storage[978] ),
    .S(net708),
    .X(_05154_));
 sg13g2_and2_1 _12099_ (.A(net413),
    .B(_05154_),
    .X(_01678_));
 sg13g2_mux2_1 _12100_ (.A0(\shift_storage.storage[97] ),
    .A1(\shift_storage.storage[96] ),
    .S(net620),
    .X(_05155_));
 sg13g2_and2_1 _12101_ (.A(net322),
    .B(_05155_),
    .X(_01679_));
 sg13g2_mux2_1 _12102_ (.A0(\shift_storage.storage[980] ),
    .A1(\shift_storage.storage[979] ),
    .S(net708),
    .X(_05156_));
 sg13g2_and2_1 _12103_ (.A(net413),
    .B(_05156_),
    .X(_01680_));
 sg13g2_mux2_1 _12104_ (.A0(\shift_storage.storage[981] ),
    .A1(\shift_storage.storage[980] ),
    .S(net708),
    .X(_05157_));
 sg13g2_and2_1 _12105_ (.A(net413),
    .B(_05157_),
    .X(_01681_));
 sg13g2_mux2_1 _12106_ (.A0(\shift_storage.storage[982] ),
    .A1(\shift_storage.storage[981] ),
    .S(net708),
    .X(_05158_));
 sg13g2_and2_1 _12107_ (.A(net414),
    .B(_05158_),
    .X(_01682_));
 sg13g2_buf_2 fanout12 (.A(net13),
    .X(net12));
 sg13g2_mux2_1 _12109_ (.A0(\shift_storage.storage[983] ),
    .A1(\shift_storage.storage[982] ),
    .S(net708),
    .X(_05160_));
 sg13g2_and2_1 _12110_ (.A(net413),
    .B(_05160_),
    .X(_01683_));
 sg13g2_mux2_1 _12111_ (.A0(\shift_storage.storage[984] ),
    .A1(\shift_storage.storage[983] ),
    .S(net708),
    .X(_05161_));
 sg13g2_and2_1 _12112_ (.A(net413),
    .B(_05161_),
    .X(_01684_));
 sg13g2_mux2_1 _12113_ (.A0(\shift_storage.storage[985] ),
    .A1(\shift_storage.storage[984] ),
    .S(net709),
    .X(_05162_));
 sg13g2_and2_1 _12114_ (.A(net414),
    .B(_05162_),
    .X(_01685_));
 sg13g2_buf_2 fanout11 (.A(_02277_),
    .X(net11));
 sg13g2_mux2_1 _12116_ (.A0(\shift_storage.storage[986] ),
    .A1(\shift_storage.storage[985] ),
    .S(net709),
    .X(_05164_));
 sg13g2_and2_1 _12117_ (.A(net414),
    .B(_05164_),
    .X(_01686_));
 sg13g2_mux2_1 _12118_ (.A0(\shift_storage.storage[987] ),
    .A1(\shift_storage.storage[986] ),
    .S(net709),
    .X(_05165_));
 sg13g2_and2_1 _12119_ (.A(net415),
    .B(_05165_),
    .X(_01687_));
 sg13g2_mux2_1 _12120_ (.A0(\shift_storage.storage[988] ),
    .A1(\shift_storage.storage[987] ),
    .S(net709),
    .X(_05166_));
 sg13g2_and2_1 _12121_ (.A(net414),
    .B(_05166_),
    .X(_01688_));
 sg13g2_mux2_1 _12122_ (.A0(\shift_storage.storage[989] ),
    .A1(\shift_storage.storage[988] ),
    .S(net710),
    .X(_05167_));
 sg13g2_and2_1 _12123_ (.A(net414),
    .B(_05167_),
    .X(_01689_));
 sg13g2_mux2_1 _12124_ (.A0(\shift_storage.storage[98] ),
    .A1(\shift_storage.storage[97] ),
    .S(net620),
    .X(_05168_));
 sg13g2_and2_1 _12125_ (.A(net322),
    .B(_05168_),
    .X(_01690_));
 sg13g2_mux2_1 _12126_ (.A0(\shift_storage.storage[990] ),
    .A1(\shift_storage.storage[989] ),
    .S(net725),
    .X(_05169_));
 sg13g2_and2_1 _12127_ (.A(net431),
    .B(_05169_),
    .X(_01691_));
 sg13g2_mux2_1 _12128_ (.A0(\shift_storage.storage[991] ),
    .A1(\shift_storage.storage[990] ),
    .S(net726),
    .X(_05170_));
 sg13g2_and2_1 _12129_ (.A(net432),
    .B(_05170_),
    .X(_01692_));
 sg13g2_buf_2 fanout10 (.A(_02569_),
    .X(net10));
 sg13g2_mux2_1 _12131_ (.A0(\shift_storage.storage[992] ),
    .A1(\shift_storage.storage[991] ),
    .S(net726),
    .X(_05172_));
 sg13g2_and2_1 _12132_ (.A(net432),
    .B(_05172_),
    .X(_01693_));
 sg13g2_mux2_1 _12133_ (.A0(\shift_storage.storage[993] ),
    .A1(\shift_storage.storage[992] ),
    .S(net725),
    .X(_05173_));
 sg13g2_and2_1 _12134_ (.A(net431),
    .B(_05173_),
    .X(_01694_));
 sg13g2_mux2_1 _12135_ (.A0(\shift_storage.storage[994] ),
    .A1(\shift_storage.storage[993] ),
    .S(net725),
    .X(_05174_));
 sg13g2_and2_1 _12136_ (.A(net431),
    .B(_05174_),
    .X(_01695_));
 sg13g2_mux2_1 _12137_ (.A0(\shift_storage.storage[995] ),
    .A1(\shift_storage.storage[994] ),
    .S(net725),
    .X(_05175_));
 sg13g2_and2_1 _12138_ (.A(net431),
    .B(_05175_),
    .X(_01696_));
 sg13g2_mux2_1 _12139_ (.A0(\shift_storage.storage[996] ),
    .A1(\shift_storage.storage[995] ),
    .S(net725),
    .X(_05176_));
 sg13g2_and2_1 _12140_ (.A(net431),
    .B(_05176_),
    .X(_01697_));
 sg13g2_mux2_1 _12141_ (.A0(\shift_storage.storage[997] ),
    .A1(\shift_storage.storage[996] ),
    .S(net725),
    .X(_05177_));
 sg13g2_and2_1 _12142_ (.A(net431),
    .B(_05177_),
    .X(_01698_));
 sg13g2_mux2_1 _12143_ (.A0(\shift_storage.storage[998] ),
    .A1(\shift_storage.storage[997] ),
    .S(net725),
    .X(_05178_));
 sg13g2_and2_1 _12144_ (.A(net431),
    .B(_05178_),
    .X(_01699_));
 sg13g2_mux2_1 _12145_ (.A0(\shift_storage.storage[999] ),
    .A1(\shift_storage.storage[998] ),
    .S(net725),
    .X(_05179_));
 sg13g2_and2_1 _12146_ (.A(net431),
    .B(_05179_),
    .X(_01700_));
 sg13g2_mux2_1 _12147_ (.A0(\shift_storage.storage[99] ),
    .A1(\shift_storage.storage[98] ),
    .S(net620),
    .X(_05180_));
 sg13g2_and2_1 _12148_ (.A(net322),
    .B(_05180_),
    .X(_01701_));
 sg13g2_mux2_1 _12149_ (.A0(\shift_storage.storage[9] ),
    .A1(\shift_storage.storage[8] ),
    .S(net609),
    .X(_05181_));
 sg13g2_and2_1 _12150_ (.A(net311),
    .B(_05181_),
    .X(_01702_));
 sg13g2_buf_2 fanout9 (.A(_02684_),
    .X(net9));
 sg13g2_inv_1 _12152_ (.Y(_05183_),
    .A(net496));
 sg13g2_buf_4 fanout8 (.X(net8),
    .A(_02881_));
 sg13g2_mux2_1 _12154_ (.A0(_02938_),
    .A1(_03038_),
    .S(net198),
    .X(_05185_));
 sg13g2_buf_8 wire7 (.A(net7),
    .X(net4023));
 sg13g2_buf_2 fanout6 (.A(_02789_),
    .X(net6));
 sg13g2_buf_2 fanout5 (.A(_02898_),
    .X(net5));
 sg13g2_nand3_1 _12158_ (.B(\median_processor.median_processor.median_out[0] ),
    .C(data_in_p2c_1),
    .A(net496),
    .Y(_05189_));
 sg13g2_nand2_1 _12159_ (.Y(_05190_),
    .A(net198),
    .B(_02938_));
 sg13g2_a21oi_1 _12160_ (.A1(_05189_),
    .A2(_05190_),
    .Y(_05191_),
    .B1(net494));
 sg13g2_a221oi_1 _12161_ (.B2(net494),
    .C1(_05191_),
    .B1(_05185_),
    .A1(_02938_),
    .Y(net34),
    .A2(_03038_));
 sg13g2_nor2b_2 _12162_ (.A(data_in_p2c_1),
    .B_N(\median_processor.median_processor.median_out[0] ),
    .Y(_05192_));
 sg13g2_o21ai_1 _12163_ (.B1(net496),
    .Y(_05193_),
    .A1(net504),
    .A2(_05192_));
 sg13g2_xor2_1 _12164_ (.B(_05192_),
    .A(net504),
    .X(_05194_));
 sg13g2_nor2_1 _12165_ (.A(net198),
    .B(\median_processor.median_processor.median_out[1] ),
    .Y(_05195_));
 sg13g2_a22oi_1 _12166_ (.Y(_05196_),
    .B1(_05194_),
    .B2(_05195_),
    .A2(_05193_),
    .A1(\median_processor.median_processor.median_out[1] ));
 sg13g2_and2_1 _12167_ (.A(\median_processor.median_processor.median_out[1] ),
    .B(net504),
    .X(_05197_));
 sg13g2_mux2_1 _12168_ (.A0(net504),
    .A1(\median_processor.median_processor.median_out[1] ),
    .S(net496),
    .X(_05198_));
 sg13g2_a22oi_1 _12169_ (.Y(_05199_),
    .B1(_05198_),
    .B2(net494),
    .A2(_05197_),
    .A1(_05192_));
 sg13g2_o21ai_1 _12170_ (.B1(_05199_),
    .Y(net33),
    .A1(net494),
    .A2(_05196_));
 sg13g2_nand2b_1 _12171_ (.Y(_05200_),
    .B(net504),
    .A_N(\median_processor.median_processor.median_out[1] ));
 sg13g2_nor2b_1 _12172_ (.A(net504),
    .B_N(\median_processor.median_processor.median_out[1] ),
    .Y(_05201_));
 sg13g2_a21o_2 _12173_ (.A2(_05200_),
    .A1(_05192_),
    .B1(_05201_),
    .X(_05202_));
 sg13g2_buf_2 fanout4 (.A(_02934_),
    .X(net4));
 sg13g2_o21ai_1 _12175_ (.B1(net496),
    .Y(_05204_),
    .A1(data_in_p2c_3),
    .A2(_05202_));
 sg13g2_nor2_1 _12176_ (.A(net198),
    .B(\median_processor.median_processor.median_out[2] ),
    .Y(_05205_));
 sg13g2_xnor2_1 _12177_ (.Y(_05206_),
    .A(_03050_),
    .B(_05202_));
 sg13g2_a22oi_1 _12178_ (.Y(_05207_),
    .B1(_05205_),
    .B2(_05206_),
    .A2(_05204_),
    .A1(\median_processor.median_processor.median_out[2] ));
 sg13g2_nand2_1 _12179_ (.Y(_05208_),
    .A(net496),
    .B(\median_processor.median_processor.median_out[2] ));
 sg13g2_o21ai_1 _12180_ (.B1(_05208_),
    .Y(_05209_),
    .A1(net496),
    .A2(_03050_));
 sg13g2_nor2_1 _12181_ (.A(_02966_),
    .B(_03050_),
    .Y(_05210_));
 sg13g2_a22oi_1 _12182_ (.Y(_05211_),
    .B1(_05210_),
    .B2(_05202_),
    .A2(_05209_),
    .A1(net494));
 sg13g2_o21ai_1 _12183_ (.B1(_05211_),
    .Y(net21),
    .A1(net494),
    .A2(_05207_));
 sg13g2_nor2_1 _12184_ (.A(_03050_),
    .B(_05202_),
    .Y(_05212_));
 sg13g2_a21oi_1 _12185_ (.A1(_03050_),
    .A2(_05202_),
    .Y(_05213_),
    .B1(\median_processor.median_processor.median_out[2] ));
 sg13g2_or2_1 _12186_ (.X(_05214_),
    .B(_05213_),
    .A(_05212_));
 sg13g2_buf_2 fanout3 (.A(net4),
    .X(net3));
 sg13g2_nor2_1 _12188_ (.A(\median_processor.median_processor.median_out[3] ),
    .B(net503),
    .Y(_05216_));
 sg13g2_nor2_1 _12189_ (.A(net198),
    .B(_02979_),
    .Y(_05217_));
 sg13g2_a21oi_1 _12190_ (.A1(net198),
    .A2(net503),
    .Y(_05218_),
    .B1(_05217_));
 sg13g2_o21ai_1 _12191_ (.B1(net496),
    .Y(_05219_),
    .A1(_03056_),
    .A2(_05214_));
 sg13g2_xnor2_1 _12192_ (.Y(_05220_),
    .A(net503),
    .B(_05214_));
 sg13g2_a22oi_1 _12193_ (.Y(_05221_),
    .B1(_05220_),
    .B2(_05217_),
    .A2(_05219_),
    .A1(_02979_));
 sg13g2_nor2_1 _12194_ (.A(net494),
    .B(_05221_),
    .Y(_05222_));
 sg13g2_a221oi_1 _12195_ (.B2(net494),
    .C1(_05222_),
    .B1(_05218_),
    .A1(_05214_),
    .Y(net16),
    .A2(_05216_));
 sg13g2_o21ai_1 _12196_ (.B1(net503),
    .Y(_05223_),
    .A1(_05212_),
    .A2(_05213_));
 sg13g2_nor3_1 _12197_ (.A(net503),
    .B(_05212_),
    .C(_05213_),
    .Y(_05224_));
 sg13g2_a21o_1 _12198_ (.A2(_05223_),
    .A1(\median_processor.median_processor.median_out[3] ),
    .B1(_05224_),
    .X(_05225_));
 sg13g2_buf_8 wire2 (.A(net2),
    .X(net4017));
 sg13g2_o21ai_1 _12200_ (.B1(net497),
    .Y(_05227_),
    .A1(net501),
    .A2(_05225_));
 sg13g2_nor2_1 _12201_ (.A(net198),
    .B(\median_processor.median_processor.median_out[4] ),
    .Y(_05228_));
 sg13g2_xor2_1 _12202_ (.B(_05225_),
    .A(net501),
    .X(_05229_));
 sg13g2_a22oi_1 _12203_ (.Y(_05230_),
    .B1(_05228_),
    .B2(_05229_),
    .A2(_05227_),
    .A1(\median_processor.median_processor.median_out[4] ));
 sg13g2_mux2_1 _12204_ (.A0(net501),
    .A1(\median_processor.median_processor.median_out[4] ),
    .S(net497),
    .X(_05231_));
 sg13g2_and2_1 _12205_ (.A(\median_processor.median_processor.median_out[4] ),
    .B(net501),
    .X(_05232_));
 sg13g2_a22oi_1 _12206_ (.Y(_05233_),
    .B1(_05232_),
    .B2(_05225_),
    .A2(_05231_),
    .A1(net495));
 sg13g2_o21ai_1 _12207_ (.B1(_05233_),
    .Y(net15),
    .A1(net495),
    .A2(_05230_));
 sg13g2_nor2b_1 _12208_ (.A(net501),
    .B_N(_05225_),
    .Y(_05234_));
 sg13g2_nand2b_1 _12209_ (.Y(_05235_),
    .B(net501),
    .A_N(_05225_));
 sg13g2_o21ai_1 _12210_ (.B1(_05235_),
    .Y(_05236_),
    .A1(\median_processor.median_processor.median_out[4] ),
    .A2(_05234_));
 sg13g2_buf_8 wire1 (.A(net1),
    .X(net4016));
 sg13g2_nor2_1 _12212_ (.A(\median_processor.median_processor.median_out[5] ),
    .B(net500),
    .Y(_05238_));
 sg13g2_mux2_1 _12213_ (.A0(_03006_),
    .A1(_03063_),
    .S(_05183_),
    .X(_05239_));
 sg13g2_o21ai_1 _12214_ (.B1(net497),
    .Y(_05240_),
    .A1(_03063_),
    .A2(_05236_));
 sg13g2_nand2_1 _12215_ (.Y(_05241_),
    .A(_03006_),
    .B(_05240_));
 sg13g2_xnor2_1 _12216_ (.Y(_05242_),
    .A(net500),
    .B(_05236_));
 sg13g2_nand3_1 _12217_ (.B(\median_processor.median_processor.median_out[5] ),
    .C(_05242_),
    .A(net497),
    .Y(_05243_));
 sg13g2_a21oi_1 _12218_ (.A1(_05241_),
    .A2(_05243_),
    .Y(_05244_),
    .B1(out_select_p2c_2));
 sg13g2_a221oi_1 _12219_ (.B2(net495),
    .C1(_05244_),
    .B1(_05239_),
    .A1(_05236_),
    .Y(net7),
    .A2(_05238_));
 sg13g2_nand2_1 _12220_ (.Y(_05245_),
    .A(net500),
    .B(_05236_));
 sg13g2_o21ai_1 _12221_ (.B1(_03006_),
    .Y(_05246_),
    .A1(net500),
    .A2(_05236_));
 sg13g2_nand2_2 _12222_ (.Y(_05247_),
    .A(_05245_),
    .B(_05246_));
 sg13g2_nor2_1 _12223_ (.A(\median_processor.median_processor.median_out[6] ),
    .B(net498),
    .Y(_05248_));
 sg13g2_nor2_1 _12224_ (.A(_05183_),
    .B(_03019_),
    .Y(_05249_));
 sg13g2_a21oi_1 _12225_ (.A1(net198),
    .A2(net498),
    .Y(_05250_),
    .B1(_05249_));
 sg13g2_o21ai_1 _12226_ (.B1(net497),
    .Y(_05251_),
    .A1(_03067_),
    .A2(_05247_));
 sg13g2_xnor2_1 _12227_ (.Y(_05252_),
    .A(net498),
    .B(_05247_));
 sg13g2_a22oi_1 _12228_ (.Y(_05253_),
    .B1(_05252_),
    .B2(_05249_),
    .A2(_05251_),
    .A1(_03019_));
 sg13g2_nor2_1 _12229_ (.A(net495),
    .B(_05253_),
    .Y(_05254_));
 sg13g2_a221oi_1 _12230_ (.B2(net495),
    .C1(_05254_),
    .B1(_05250_),
    .A1(_05247_),
    .Y(net2),
    .A2(_05248_));
 sg13g2_nor2_1 _12231_ (.A(net498),
    .B(_05247_),
    .Y(_05255_));
 sg13g2_a21oi_1 _12232_ (.A1(net498),
    .A2(_05247_),
    .Y(_05256_),
    .B1(_03019_));
 sg13g2_nor2_1 _12233_ (.A(_05255_),
    .B(_05256_),
    .Y(_05257_));
 sg13g2_nor2_1 _12234_ (.A(\median_processor.median_processor.median_out[7] ),
    .B(data_in_p2c_8),
    .Y(_05258_));
 sg13g2_mux2_1 _12235_ (.A0(_03032_),
    .A1(_03071_),
    .S(_05183_),
    .X(_05259_));
 sg13g2_o21ai_1 _12236_ (.B1(net497),
    .Y(_05260_),
    .A1(_03071_),
    .A2(_05257_));
 sg13g2_nand2_1 _12237_ (.Y(_05261_),
    .A(_03032_),
    .B(_05260_));
 sg13g2_xnor2_1 _12238_ (.Y(_05262_),
    .A(data_in_p2c_8),
    .B(_05257_));
 sg13g2_nand3_1 _12239_ (.B(\median_processor.median_processor.median_out[7] ),
    .C(_05262_),
    .A(net497),
    .Y(_05263_));
 sg13g2_a21oi_1 _12240_ (.A1(_05261_),
    .A2(_05263_),
    .Y(_05264_),
    .B1(net495));
 sg13g2_a221oi_1 _12241_ (.B2(net495),
    .C1(_05264_),
    .B1(_05259_),
    .A1(_05257_),
    .Y(net1),
    .A2(_05258_));
 sg13g2_buf_4 clkbuf_leaf_0_clk_p2c (.X(clknet_leaf_0_clk_p2c),
    .A(clknet_5_0__leaf_clk_p2c));
 sg13g2_dfrbp_1 \median_processor.input_storage[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_117_clk_p2c),
    .RESET_B(net776),
    .D(_00000_),
    .Q_N(_06967_),
    .Q(\median_processor.input_storage[0] ));
 sg13g2_dfrbp_1 \median_processor.input_storage[10]$_SDFFE_PN0P_  (.CLK(clknet_leaf_118_clk_p2c),
    .RESET_B(net777),
    .D(_00001_),
    .Q_N(_06966_),
    .Q(\median_processor.input_storage[10] ));
 sg13g2_dfrbp_1 \median_processor.input_storage[11]$_SDFFE_PN0P_  (.CLK(clknet_leaf_159_clk_p2c),
    .RESET_B(net778),
    .D(_00002_),
    .Q_N(_06965_),
    .Q(\median_processor.input_storage[11] ));
 sg13g2_dfrbp_1 \median_processor.input_storage[12]$_SDFFE_PN0P_  (.CLK(clknet_leaf_157_clk_p2c),
    .RESET_B(net779),
    .D(_00003_),
    .Q_N(_06964_),
    .Q(\median_processor.input_storage[12] ));
 sg13g2_dfrbp_1 \median_processor.input_storage[13]$_SDFFE_PN0P_  (.CLK(clknet_leaf_155_clk_p2c),
    .RESET_B(net780),
    .D(_00004_),
    .Q_N(_06963_),
    .Q(\median_processor.input_storage[13] ));
 sg13g2_dfrbp_1 \median_processor.input_storage[14]$_SDFFE_PN0P_  (.CLK(clknet_leaf_155_clk_p2c),
    .RESET_B(net781),
    .D(_00005_),
    .Q_N(_06962_),
    .Q(\median_processor.input_storage[14] ));
 sg13g2_dfrbp_1 \median_processor.input_storage[15]$_SDFFE_PN0P_  (.CLK(clknet_leaf_144_clk_p2c),
    .RESET_B(net782),
    .D(_00006_),
    .Q_N(_06961_),
    .Q(\median_processor.input_storage[15] ));
 sg13g2_dfrbp_1 \median_processor.input_storage[16]$_SDFFE_PN0P_  (.CLK(clknet_leaf_118_clk_p2c),
    .RESET_B(net783),
    .D(_00007_),
    .Q_N(_06960_),
    .Q(\median_processor.input_storage[16] ));
 sg13g2_dfrbp_1 \median_processor.input_storage[17]$_SDFFE_PN0P_  (.CLK(clknet_leaf_128_clk_p2c),
    .RESET_B(net784),
    .D(_00008_),
    .Q_N(_06959_),
    .Q(\median_processor.input_storage[17] ));
 sg13g2_dfrbp_1 \median_processor.input_storage[18]$_SDFFE_PN0P_  (.CLK(clknet_leaf_132_clk_p2c),
    .RESET_B(net785),
    .D(_00009_),
    .Q_N(_06958_),
    .Q(\median_processor.input_storage[18] ));
 sg13g2_dfrbp_1 \median_processor.input_storage[19]$_SDFFE_PN0P_  (.CLK(clknet_leaf_132_clk_p2c),
    .RESET_B(net786),
    .D(_00010_),
    .Q_N(_06957_),
    .Q(\median_processor.input_storage[19] ));
 sg13g2_dfrbp_1 \median_processor.input_storage[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_118_clk_p2c),
    .RESET_B(net787),
    .D(_00011_),
    .Q_N(_06956_),
    .Q(\median_processor.input_storage[1] ));
 sg13g2_dfrbp_1 \median_processor.input_storage[20]$_SDFFE_PN0P_  (.CLK(clknet_leaf_134_clk_p2c),
    .RESET_B(net788),
    .D(_00012_),
    .Q_N(_06955_),
    .Q(\median_processor.input_storage[20] ));
 sg13g2_dfrbp_1 \median_processor.input_storage[21]$_SDFFE_PN0P_  (.CLK(clknet_leaf_157_clk_p2c),
    .RESET_B(net789),
    .D(_00013_),
    .Q_N(_06954_),
    .Q(\median_processor.input_storage[21] ));
 sg13g2_dfrbp_1 \median_processor.input_storage[22]$_SDFFE_PN0P_  (.CLK(clknet_leaf_143_clk_p2c),
    .RESET_B(net790),
    .D(_00014_),
    .Q_N(_06953_),
    .Q(\median_processor.input_storage[22] ));
 sg13g2_dfrbp_1 \median_processor.input_storage[23]$_SDFFE_PN0P_  (.CLK(clknet_leaf_142_clk_p2c),
    .RESET_B(net791),
    .D(_00015_),
    .Q_N(_06952_),
    .Q(\median_processor.input_storage[23] ));
 sg13g2_dfrbp_1 \median_processor.input_storage[24]$_SDFFE_PN0P_  (.CLK(clknet_leaf_133_clk_p2c),
    .RESET_B(net792),
    .D(_00016_),
    .Q_N(_06951_),
    .Q(\median_processor.input_storage[24] ));
 sg13g2_dfrbp_1 \median_processor.input_storage[25]$_SDFFE_PN0P_  (.CLK(clknet_leaf_133_clk_p2c),
    .RESET_B(net793),
    .D(_00017_),
    .Q_N(_06950_),
    .Q(\median_processor.input_storage[25] ));
 sg13g2_dfrbp_1 \median_processor.input_storage[26]$_SDFFE_PN0P_  (.CLK(clknet_leaf_130_clk_p2c),
    .RESET_B(net794),
    .D(_00018_),
    .Q_N(_06949_),
    .Q(\median_processor.input_storage[26] ));
 sg13g2_dfrbp_1 \median_processor.input_storage[27]$_SDFFE_PN0P_  (.CLK(clknet_leaf_131_clk_p2c),
    .RESET_B(net795),
    .D(_00019_),
    .Q_N(_06948_),
    .Q(\median_processor.input_storage[27] ));
 sg13g2_dfrbp_1 \median_processor.input_storage[28]$_SDFFE_PN0P_  (.CLK(clknet_leaf_135_clk_p2c),
    .RESET_B(net796),
    .D(_00020_),
    .Q_N(_06947_),
    .Q(\median_processor.input_storage[28] ));
 sg13g2_dfrbp_1 \median_processor.input_storage[29]$_SDFFE_PN0P_  (.CLK(clknet_leaf_156_clk_p2c),
    .RESET_B(net797),
    .D(_00021_),
    .Q_N(_06946_),
    .Q(\median_processor.input_storage[29] ));
 sg13g2_dfrbp_1 \median_processor.input_storage[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_157_clk_p2c),
    .RESET_B(net798),
    .D(_00022_),
    .Q_N(_06945_),
    .Q(\median_processor.input_storage[2] ));
 sg13g2_dfrbp_1 \median_processor.input_storage[30]$_SDFFE_PN0P_  (.CLK(clknet_leaf_144_clk_p2c),
    .RESET_B(net799),
    .D(_00023_),
    .Q_N(_06944_),
    .Q(\median_processor.input_storage[30] ));
 sg13g2_dfrbp_1 \median_processor.input_storage[31]$_SDFFE_PN0P_  (.CLK(clknet_leaf_144_clk_p2c),
    .RESET_B(net800),
    .D(_00024_),
    .Q_N(_06943_),
    .Q(\median_processor.input_storage[31] ));
 sg13g2_dfrbp_1 \median_processor.input_storage[32]$_SDFFE_PN0P_  (.CLK(clknet_leaf_129_clk_p2c),
    .RESET_B(net801),
    .D(_00025_),
    .Q_N(_06942_),
    .Q(\median_processor.input_storage[32] ));
 sg13g2_dfrbp_1 \median_processor.input_storage[33]$_SDFFE_PN0P_  (.CLK(clknet_leaf_129_clk_p2c),
    .RESET_B(net802),
    .D(_00026_),
    .Q_N(_06941_),
    .Q(\median_processor.input_storage[33] ));
 sg13g2_dfrbp_1 \median_processor.input_storage[34]$_SDFFE_PN0P_  (.CLK(clknet_leaf_129_clk_p2c),
    .RESET_B(net803),
    .D(_00027_),
    .Q_N(_06940_),
    .Q(\median_processor.input_storage[34] ));
 sg13g2_dfrbp_1 \median_processor.input_storage[35]$_SDFFE_PN0P_  (.CLK(clknet_leaf_132_clk_p2c),
    .RESET_B(net804),
    .D(_00028_),
    .Q_N(_06939_),
    .Q(\median_processor.input_storage[35] ));
 sg13g2_dfrbp_1 \median_processor.input_storage[36]$_SDFFE_PN0P_  (.CLK(clknet_leaf_134_clk_p2c),
    .RESET_B(net805),
    .D(_00029_),
    .Q_N(_06938_),
    .Q(\median_processor.input_storage[36] ));
 sg13g2_dfrbp_1 \median_processor.input_storage[37]$_SDFFE_PN0P_  (.CLK(clknet_leaf_156_clk_p2c),
    .RESET_B(net806),
    .D(_00030_),
    .Q_N(_06937_),
    .Q(\median_processor.input_storage[37] ));
 sg13g2_dfrbp_1 \median_processor.input_storage[38]$_SDFFE_PN0P_  (.CLK(clknet_leaf_144_clk_p2c),
    .RESET_B(net807),
    .D(_00031_),
    .Q_N(_06936_),
    .Q(\median_processor.input_storage[38] ));
 sg13g2_dfrbp_1 \median_processor.input_storage[39]$_SDFFE_PN0P_  (.CLK(clknet_leaf_136_clk_p2c),
    .RESET_B(net808),
    .D(_00032_),
    .Q_N(_06935_),
    .Q(\median_processor.input_storage[39] ));
 sg13g2_dfrbp_1 \median_processor.input_storage[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_159_clk_p2c),
    .RESET_B(net809),
    .D(_00033_),
    .Q_N(_06934_),
    .Q(\median_processor.input_storage[3] ));
 sg13g2_dfrbp_1 \median_processor.input_storage[40]$_SDFFE_PN0P_  (.CLK(clknet_leaf_119_clk_p2c),
    .RESET_B(net810),
    .D(_00034_),
    .Q_N(_06933_),
    .Q(\median_processor.input_storage[40] ));
 sg13g2_dfrbp_1 \median_processor.input_storage[41]$_SDFFE_PN0P_  (.CLK(clknet_leaf_118_clk_p2c),
    .RESET_B(net811),
    .D(_00035_),
    .Q_N(_06932_),
    .Q(\median_processor.input_storage[41] ));
 sg13g2_dfrbp_1 \median_processor.input_storage[42]$_SDFFE_PN0P_  (.CLK(clknet_leaf_119_clk_p2c),
    .RESET_B(net812),
    .D(_00036_),
    .Q_N(_06931_),
    .Q(\median_processor.input_storage[42] ));
 sg13g2_dfrbp_1 \median_processor.input_storage[43]$_SDFFE_PN0P_  (.CLK(clknet_leaf_118_clk_p2c),
    .RESET_B(net813),
    .D(_00037_),
    .Q_N(_06930_),
    .Q(\median_processor.input_storage[43] ));
 sg13g2_dfrbp_1 \median_processor.input_storage[44]$_SDFFE_PN0P_  (.CLK(clknet_leaf_157_clk_p2c),
    .RESET_B(net814),
    .D(_00038_),
    .Q_N(_06929_),
    .Q(\median_processor.input_storage[44] ));
 sg13g2_dfrbp_1 \median_processor.input_storage[45]$_SDFFE_PN0P_  (.CLK(clknet_leaf_143_clk_p2c),
    .RESET_B(net815),
    .D(_00039_),
    .Q_N(_06928_),
    .Q(\median_processor.input_storage[45] ));
 sg13g2_dfrbp_1 \median_processor.input_storage[46]$_SDFFE_PN0P_  (.CLK(clknet_leaf_143_clk_p2c),
    .RESET_B(net816),
    .D(_00040_),
    .Q_N(_06927_),
    .Q(\median_processor.input_storage[46] ));
 sg13g2_dfrbp_1 \median_processor.input_storage[47]$_SDFFE_PN0P_  (.CLK(clknet_leaf_134_clk_p2c),
    .RESET_B(net817),
    .D(_00041_),
    .Q_N(_06926_),
    .Q(\median_processor.input_storage[47] ));
 sg13g2_dfrbp_1 \median_processor.input_storage[48]$_SDFFE_PN0P_  (.CLK(clknet_leaf_128_clk_p2c),
    .RESET_B(net818),
    .D(_00042_),
    .Q_N(_06925_),
    .Q(\median_processor.input_storage[48] ));
 sg13g2_dfrbp_1 \median_processor.input_storage[49]$_SDFFE_PN0P_  (.CLK(clknet_leaf_128_clk_p2c),
    .RESET_B(net819),
    .D(_00043_),
    .Q_N(_06924_),
    .Q(\median_processor.input_storage[49] ));
 sg13g2_dfrbp_1 \median_processor.input_storage[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_157_clk_p2c),
    .RESET_B(net820),
    .D(_00044_),
    .Q_N(_06923_),
    .Q(\median_processor.input_storage[4] ));
 sg13g2_dfrbp_1 \median_processor.input_storage[50]$_SDFFE_PN0P_  (.CLK(clknet_leaf_129_clk_p2c),
    .RESET_B(net821),
    .D(_00045_),
    .Q_N(_06922_),
    .Q(\median_processor.input_storage[50] ));
 sg13g2_dfrbp_1 \median_processor.input_storage[51]$_SDFFE_PN0P_  (.CLK(clknet_leaf_131_clk_p2c),
    .RESET_B(net822),
    .D(_00046_),
    .Q_N(_06921_),
    .Q(\median_processor.input_storage[51] ));
 sg13g2_dfrbp_1 \median_processor.input_storage[52]$_SDFFE_PN0P_  (.CLK(clknet_leaf_134_clk_p2c),
    .RESET_B(net823),
    .D(_00047_),
    .Q_N(_06920_),
    .Q(\median_processor.input_storage[52] ));
 sg13g2_dfrbp_1 \median_processor.input_storage[53]$_SDFFE_PN0P_  (.CLK(clknet_leaf_143_clk_p2c),
    .RESET_B(net824),
    .D(_00048_),
    .Q_N(_06919_),
    .Q(\median_processor.input_storage[53] ));
 sg13g2_dfrbp_1 \median_processor.input_storage[54]$_SDFFE_PN0P_  (.CLK(clknet_leaf_136_clk_p2c),
    .RESET_B(net825),
    .D(_00049_),
    .Q_N(_06918_),
    .Q(\median_processor.input_storage[54] ));
 sg13g2_dfrbp_1 \median_processor.input_storage[55]$_SDFFE_PN0P_  (.CLK(clknet_leaf_137_clk_p2c),
    .RESET_B(net826),
    .D(_00050_),
    .Q_N(_06917_),
    .Q(\median_processor.input_storage[55] ));
 sg13g2_dfrbp_1 \median_processor.input_storage[56]$_SDFFE_PN0P_  (.CLK(clknet_leaf_117_clk_p2c),
    .RESET_B(net827),
    .D(_00051_),
    .Q_N(_06916_),
    .Q(\median_processor.input_storage[56] ));
 sg13g2_dfrbp_1 \median_processor.input_storage[57]$_SDFFE_PN0P_  (.CLK(clknet_leaf_117_clk_p2c),
    .RESET_B(net828),
    .D(_00052_),
    .Q_N(_06915_),
    .Q(\median_processor.input_storage[57] ));
 sg13g2_dfrbp_1 \median_processor.input_storage[58]$_SDFFE_PN0P_  (.CLK(clknet_leaf_157_clk_p2c),
    .RESET_B(net829),
    .D(_00053_),
    .Q_N(_06914_),
    .Q(\median_processor.input_storage[58] ));
 sg13g2_dfrbp_1 \median_processor.input_storage[59]$_SDFFE_PN0P_  (.CLK(clknet_leaf_159_clk_p2c),
    .RESET_B(net830),
    .D(_00054_),
    .Q_N(_06913_),
    .Q(\median_processor.input_storage[59] ));
 sg13g2_dfrbp_1 \median_processor.input_storage[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_155_clk_p2c),
    .RESET_B(net831),
    .D(_00055_),
    .Q_N(_06912_),
    .Q(\median_processor.input_storage[5] ));
 sg13g2_dfrbp_1 \median_processor.input_storage[60]$_SDFFE_PN0P_  (.CLK(clknet_leaf_158_clk_p2c),
    .RESET_B(net832),
    .D(_00056_),
    .Q_N(_06911_),
    .Q(\median_processor.input_storage[60] ));
 sg13g2_dfrbp_1 \median_processor.input_storage[61]$_SDFFE_PN0P_  (.CLK(clknet_leaf_156_clk_p2c),
    .RESET_B(net833),
    .D(_00057_),
    .Q_N(_06910_),
    .Q(\median_processor.input_storage[61] ));
 sg13g2_dfrbp_1 \median_processor.input_storage[62]$_SDFFE_PN0P_  (.CLK(clknet_leaf_155_clk_p2c),
    .RESET_B(net834),
    .D(_00058_),
    .Q_N(_06909_),
    .Q(\median_processor.input_storage[62] ));
 sg13g2_dfrbp_1 \median_processor.input_storage[63]$_SDFFE_PN0P_  (.CLK(clknet_leaf_144_clk_p2c),
    .RESET_B(net835),
    .D(_00059_),
    .Q_N(_06908_),
    .Q(\median_processor.input_storage[63] ));
 sg13g2_dfrbp_1 \median_processor.input_storage[6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_145_clk_p2c),
    .RESET_B(net836),
    .D(_00060_),
    .Q_N(_06907_),
    .Q(\median_processor.input_storage[6] ));
 sg13g2_dfrbp_1 \median_processor.input_storage[7]$_SDFFE_PN0P_  (.CLK(clknet_leaf_144_clk_p2c),
    .RESET_B(net837),
    .D(_00061_),
    .Q_N(_06906_),
    .Q(\median_processor.input_storage[7] ));
 sg13g2_dfrbp_1 \median_processor.input_storage[8]$_SDFFE_PN0P_  (.CLK(clknet_leaf_117_clk_p2c),
    .RESET_B(net838),
    .D(_00062_),
    .Q_N(_06905_),
    .Q(\median_processor.input_storage[8] ));
 sg13g2_dfrbp_1 \median_processor.input_storage[9]$_SDFFE_PN0P_  (.CLK(clknet_leaf_117_clk_p2c),
    .RESET_B(net839),
    .D(_00063_),
    .Q_N(_06904_),
    .Q(\median_processor.input_storage[9] ));
 sg13g2_dfrbp_1 \median_processor.median_processor.median_out[0]$_DFFE_PP_  (.CLK(clknet_leaf_117_clk_p2c),
    .RESET_B(net840),
    .D(_00064_),
    .Q_N(_06903_),
    .Q(\median_processor.median_processor.median_out[0] ));
 sg13g2_dfrbp_1 \median_processor.median_processor.median_out[1]$_DFFE_PP_  (.CLK(clknet_leaf_120_clk_p2c),
    .RESET_B(net841),
    .D(_00065_),
    .Q_N(_06902_),
    .Q(\median_processor.median_processor.median_out[1] ));
 sg13g2_dfrbp_1 \median_processor.median_processor.median_out[2]$_DFFE_PP_  (.CLK(clknet_leaf_116_clk_p2c),
    .RESET_B(net842),
    .D(_00066_),
    .Q_N(_06901_),
    .Q(\median_processor.median_processor.median_out[2] ));
 sg13g2_dfrbp_1 \median_processor.median_processor.median_out[3]$_DFFE_PP_  (.CLK(clknet_leaf_116_clk_p2c),
    .RESET_B(net843),
    .D(_00067_),
    .Q_N(_06900_),
    .Q(\median_processor.median_processor.median_out[3] ));
 sg13g2_dfrbp_1 \median_processor.median_processor.median_out[4]$_DFFE_PP_  (.CLK(clknet_leaf_158_clk_p2c),
    .RESET_B(net844),
    .D(_00068_),
    .Q_N(_06899_),
    .Q(\median_processor.median_processor.median_out[4] ));
 sg13g2_dfrbp_1 \median_processor.median_processor.median_out[5]$_DFFE_PP_  (.CLK(clknet_leaf_156_clk_p2c),
    .RESET_B(net845),
    .D(_00069_),
    .Q_N(_06898_),
    .Q(\median_processor.median_processor.median_out[5] ));
 sg13g2_dfrbp_1 \median_processor.median_processor.median_out[6]$_DFFE_PP_  (.CLK(clknet_leaf_145_clk_p2c),
    .RESET_B(net846),
    .D(_00070_),
    .Q_N(_06897_),
    .Q(\median_processor.median_processor.median_out[6] ));
 sg13g2_dfrbp_1 \median_processor.median_processor.median_out[7]$_DFFE_PP_  (.CLK(clknet_leaf_145_clk_p2c),
    .RESET_B(net847),
    .D(_00071_),
    .Q_N(_06896_),
    .Q(\median_processor.median_processor.median_out[7] ));
 sg13g2_IOPadIn port_aux_enable_cell (.p2c(aux_enable_p2c),
    .pad(aux_enable_pad));
 sg13g2_IOPadIn port_clk_cell (.p2c(clk_p2c),
    .pad(clk_pad));
 sg13g2_IOPadIn port_data_in1_cell (.p2c(data_in_p2c_1),
    .pad(data_in_pad[0]));
 sg13g2_IOPadIn port_data_in2_cell (.p2c(data_in_p2c_2),
    .pad(data_in_pad[1]));
 sg13g2_IOPadIn port_data_in3_cell (.p2c(data_in_p2c_3),
    .pad(data_in_pad[2]));
 sg13g2_IOPadIn port_data_in4_cell (.p2c(data_in_p2c_4),
    .pad(data_in_pad[3]));
 sg13g2_IOPadIn port_data_in5_cell (.p2c(data_in_p2c_5),
    .pad(data_in_pad[4]));
 sg13g2_IOPadIn port_data_in6_cell (.p2c(data_in_p2c_6),
    .pad(data_in_pad[5]));
 sg13g2_IOPadIn port_data_in7_cell (.p2c(data_in_p2c_7),
    .pad(data_in_pad[6]));
 sg13g2_IOPadIn port_data_in8_cell (.p2c(data_in_p2c_8),
    .pad(data_in_pad[7]));
 sg13g2_IOPadOut16mA port_data_out1_cell (.c2p(net4050),
    .pad(data_out_pad[0]));
 sg13g2_IOPadOut16mA port_data_out2_cell (.c2p(net4049),
    .pad(data_out_pad[1]));
 sg13g2_IOPadOut16mA port_data_out3_cell (.c2p(net4037),
    .pad(data_out_pad[2]));
 sg13g2_IOPadOut16mA port_data_out4_cell (.c2p(net4032),
    .pad(data_out_pad[3]));
 sg13g2_IOPadOut16mA port_data_out5_cell (.c2p(net4031),
    .pad(data_out_pad[4]));
 sg13g2_IOPadOut16mA port_data_out6_cell (.c2p(net4023),
    .pad(data_out_pad[5]));
 sg13g2_IOPadOut16mA port_data_out7_cell (.c2p(net4017),
    .pad(data_out_pad[6]));
 sg13g2_IOPadOut16mA port_data_out8_cell (.c2p(net4016),
    .pad(data_out_pad[7]));
 sg13g2_IOPadOut16mA port_lfsr_out_cell (.c2p(lfsr_out_c2p),
    .pad(lfsr_out_pad));
 sg13g2_IOPadIn port_out_select1_cell (.p2c(out_select_p2c_1),
    .pad(out_select_pad[0]));
 sg13g2_IOPadIn port_out_select2_cell (.p2c(out_select_p2c_2),
    .pad(out_select_pad[1]));
 sg13g2_IOPadIn port_reg_addr1_cell (.p2c(reg_addr_p2c_1),
    .pad(reg_addr_pad[0]));
 sg13g2_IOPadIn port_reg_addr2_cell (.p2c(reg_addr_p2c_2),
    .pad(reg_addr_pad[1]));
 sg13g2_IOPadIn port_reg_addr3_cell (.p2c(reg_addr_p2c_3),
    .pad(reg_addr_pad[2]));
 sg13g2_IOPadIn port_rst_cell (.p2c(\median_processor.rst ),
    .pad(rst_pad));
 sg13g2_IOPadIn port_shreg_in_cell (.p2c(\shift_storage.shreg_in ),
    .pad(shreg_in_pad));
 sg13g2_IOPadOut16mA port_shreg_out_cell (.c2p(\shift_storage.shreg_out ),
    .pad(shreg_out_pad));
 sg13g2_IOPadIn port_wr_enable_cell (.p2c(\median_processor.wr_enable ),
    .pad(wr_enable_pad));
 sg13g2_dfrbp_1 \rando_generator.lfsr_reg[0]$_SDFF_PN0_  (.CLK(clknet_leaf_78_clk_p2c),
    .RESET_B(net848),
    .D(_00072_),
    .Q_N(_06895_),
    .Q(lfsr_out_c2p));
 sg13g2_dfrbp_1 \rando_generator.lfsr_reg[10]$_SDFF_PN0_  (.CLK(clknet_leaf_75_clk_p2c),
    .RESET_B(net849),
    .D(_00073_),
    .Q_N(_06894_),
    .Q(\rando_generator.lfsr_reg[10] ));
 sg13g2_dfrbp_1 \rando_generator.lfsr_reg[11]$_SDFF_PN0_  (.CLK(clknet_leaf_75_clk_p2c),
    .RESET_B(net850),
    .D(_00074_),
    .Q_N(_06893_),
    .Q(\rando_generator.lfsr_reg[11] ));
 sg13g2_dfrbp_1 \rando_generator.lfsr_reg[12]$_SDFF_PN0_  (.CLK(clknet_leaf_75_clk_p2c),
    .RESET_B(net851),
    .D(_00075_),
    .Q_N(_06892_),
    .Q(\rando_generator.lfsr_reg[12] ));
 sg13g2_dfrbp_1 \rando_generator.lfsr_reg[13]$_SDFF_PN0_  (.CLK(clknet_leaf_74_clk_p2c),
    .RESET_B(net852),
    .D(_00076_),
    .Q_N(_06891_),
    .Q(\rando_generator.lfsr_reg[13] ));
 sg13g2_dfrbp_1 \rando_generator.lfsr_reg[14]$_SDFF_PN0_  (.CLK(clknet_leaf_75_clk_p2c),
    .RESET_B(net853),
    .D(_00077_),
    .Q_N(_06890_),
    .Q(\rando_generator.lfsr_reg[14] ));
 sg13g2_dfrbp_1 \rando_generator.lfsr_reg[15]$_SDFF_PN0_  (.CLK(clknet_leaf_80_clk_p2c),
    .RESET_B(net854),
    .D(_00078_),
    .Q_N(_06889_),
    .Q(\rando_generator.lfsr_reg[15] ));
 sg13g2_dfrbp_1 \rando_generator.lfsr_reg[16]$_SDFF_PN0_  (.CLK(clknet_leaf_80_clk_p2c),
    .RESET_B(net855),
    .D(_00079_),
    .Q_N(_06888_),
    .Q(\rando_generator.lfsr_reg[16] ));
 sg13g2_dfrbp_1 \rando_generator.lfsr_reg[17]$_SDFF_PN0_  (.CLK(clknet_leaf_80_clk_p2c),
    .RESET_B(net856),
    .D(_00080_),
    .Q_N(_06887_),
    .Q(\rando_generator.lfsr_reg[17] ));
 sg13g2_dfrbp_1 \rando_generator.lfsr_reg[18]$_SDFF_PN0_  (.CLK(clknet_leaf_80_clk_p2c),
    .RESET_B(net857),
    .D(_00081_),
    .Q_N(_06886_),
    .Q(\rando_generator.lfsr_reg[18] ));
 sg13g2_dfrbp_1 \rando_generator.lfsr_reg[19]$_SDFF_PN0_  (.CLK(clknet_leaf_80_clk_p2c),
    .RESET_B(net858),
    .D(_00082_),
    .Q_N(_06885_),
    .Q(\rando_generator.lfsr_reg[19] ));
 sg13g2_dfrbp_1 \rando_generator.lfsr_reg[1]$_SDFF_PN0_  (.CLK(clknet_leaf_77_clk_p2c),
    .RESET_B(net859),
    .D(_00083_),
    .Q_N(_06884_),
    .Q(\rando_generator.lfsr_reg[1] ));
 sg13g2_dfrbp_1 \rando_generator.lfsr_reg[20]$_SDFF_PN0_  (.CLK(clknet_leaf_79_clk_p2c),
    .RESET_B(net860),
    .D(_00084_),
    .Q_N(_06883_),
    .Q(\rando_generator.lfsr_reg[20] ));
 sg13g2_dfrbp_1 \rando_generator.lfsr_reg[21]$_SDFF_PN0_  (.CLK(clknet_leaf_79_clk_p2c),
    .RESET_B(net861),
    .D(_00085_),
    .Q_N(_06882_),
    .Q(\rando_generator.lfsr_reg[21] ));
 sg13g2_dfrbp_1 \rando_generator.lfsr_reg[22]$_SDFF_PN0_  (.CLK(clknet_leaf_79_clk_p2c),
    .RESET_B(net862),
    .D(_00086_),
    .Q_N(_06881_),
    .Q(\rando_generator.lfsr_reg[22] ));
 sg13g2_dfrbp_1 \rando_generator.lfsr_reg[23]$_SDFF_PN0_  (.CLK(clknet_leaf_79_clk_p2c),
    .RESET_B(net863),
    .D(_00087_),
    .Q_N(_06880_),
    .Q(\rando_generator.lfsr_reg[23] ));
 sg13g2_dfrbp_1 \rando_generator.lfsr_reg[24]$_SDFF_PN0_  (.CLK(clknet_leaf_79_clk_p2c),
    .RESET_B(net864),
    .D(_00088_),
    .Q_N(_06879_),
    .Q(\rando_generator.lfsr_reg[24] ));
 sg13g2_dfrbp_1 \rando_generator.lfsr_reg[25]$_SDFF_PN0_  (.CLK(clknet_leaf_79_clk_p2c),
    .RESET_B(net865),
    .D(_00089_),
    .Q_N(_06878_),
    .Q(\rando_generator.lfsr_reg[25] ));
 sg13g2_dfrbp_1 \rando_generator.lfsr_reg[26]$_SDFF_PN0_  (.CLK(clknet_leaf_78_clk_p2c),
    .RESET_B(net866),
    .D(_00090_),
    .Q_N(_06877_),
    .Q(\rando_generator.lfsr_reg[26] ));
 sg13g2_dfrbp_1 \rando_generator.lfsr_reg[27]$_SDFF_PN0_  (.CLK(clknet_leaf_78_clk_p2c),
    .RESET_B(net867),
    .D(_00091_),
    .Q_N(_06876_),
    .Q(\rando_generator.lfsr_reg[27] ));
 sg13g2_dfrbp_1 \rando_generator.lfsr_reg[28]$_SDFF_PN0_  (.CLK(clknet_leaf_78_clk_p2c),
    .RESET_B(net868),
    .D(_00092_),
    .Q_N(_06875_),
    .Q(\rando_generator.lfsr_reg[28] ));
 sg13g2_dfrbp_1 \rando_generator.lfsr_reg[29]$_SDFF_PN0_  (.CLK(clknet_leaf_78_clk_p2c),
    .RESET_B(net869),
    .D(_00093_),
    .Q_N(_06874_),
    .Q(\rando_generator.lfsr_reg[29] ));
 sg13g2_dfrbp_1 \rando_generator.lfsr_reg[2]$_SDFF_PN0_  (.CLK(clknet_leaf_77_clk_p2c),
    .RESET_B(net870),
    .D(_00094_),
    .Q_N(_06873_),
    .Q(\rando_generator.lfsr_reg[2] ));
 sg13g2_dfrbp_1 \rando_generator.lfsr_reg[30]$_SDFF_PN0_  (.CLK(clknet_leaf_78_clk_p2c),
    .RESET_B(net871),
    .D(_00095_),
    .Q_N(_06872_),
    .Q(\rando_generator.lfsr_reg[30] ));
 sg13g2_dfrbp_1 \rando_generator.lfsr_reg[3]$_SDFF_PN0_  (.CLK(clknet_leaf_77_clk_p2c),
    .RESET_B(net872),
    .D(_00096_),
    .Q_N(_06871_),
    .Q(\rando_generator.lfsr_reg[3] ));
 sg13g2_dfrbp_1 \rando_generator.lfsr_reg[4]$_SDFF_PN0_  (.CLK(clknet_leaf_77_clk_p2c),
    .RESET_B(net873),
    .D(_00097_),
    .Q_N(_06870_),
    .Q(\rando_generator.lfsr_reg[4] ));
 sg13g2_dfrbp_1 \rando_generator.lfsr_reg[5]$_SDFF_PN0_  (.CLK(clknet_leaf_76_clk_p2c),
    .RESET_B(net874),
    .D(_00098_),
    .Q_N(_06869_),
    .Q(\rando_generator.lfsr_reg[5] ));
 sg13g2_dfrbp_1 \rando_generator.lfsr_reg[6]$_SDFF_PN0_  (.CLK(clknet_leaf_77_clk_p2c),
    .RESET_B(net875),
    .D(_00099_),
    .Q_N(_06868_),
    .Q(\rando_generator.lfsr_reg[6] ));
 sg13g2_dfrbp_1 \rando_generator.lfsr_reg[7]$_SDFF_PN0_  (.CLK(clknet_leaf_78_clk_p2c),
    .RESET_B(net876),
    .D(_00100_),
    .Q_N(_06867_),
    .Q(\rando_generator.lfsr_reg[7] ));
 sg13g2_dfrbp_1 \rando_generator.lfsr_reg[8]$_SDFF_PN0_  (.CLK(clknet_leaf_76_clk_p2c),
    .RESET_B(net877),
    .D(_00101_),
    .Q_N(_06866_),
    .Q(\rando_generator.lfsr_reg[8] ));
 sg13g2_dfrbp_1 \rando_generator.lfsr_reg[9]$_SDFF_PN0_  (.CLK(clknet_leaf_80_clk_p2c),
    .RESET_B(net878),
    .D(_00102_),
    .Q_N(_06865_),
    .Q(\rando_generator.lfsr_reg[9] ));
 sg13g2_dfrbp_1 \shift_storage.storage[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_77_clk_p2c),
    .RESET_B(net879),
    .D(_00103_),
    .Q_N(_06864_),
    .Q(\shift_storage.storage[0] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1000]$_SDFFE_PN0P_  (.CLK(clknet_leaf_197_clk_p2c),
    .RESET_B(net880),
    .D(_00104_),
    .Q_N(_06863_),
    .Q(\shift_storage.storage[1000] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1001]$_SDFFE_PN0P_  (.CLK(clknet_leaf_190_clk_p2c),
    .RESET_B(net881),
    .D(_00105_),
    .Q_N(_06862_),
    .Q(\shift_storage.storage[1001] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1002]$_SDFFE_PN0P_  (.CLK(clknet_leaf_190_clk_p2c),
    .RESET_B(net882),
    .D(_00106_),
    .Q_N(_06861_),
    .Q(\shift_storage.storage[1002] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1003]$_SDFFE_PN0P_  (.CLK(clknet_leaf_190_clk_p2c),
    .RESET_B(net883),
    .D(_00107_),
    .Q_N(_06860_),
    .Q(\shift_storage.storage[1003] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1004]$_SDFFE_PN0P_  (.CLK(clknet_leaf_191_clk_p2c),
    .RESET_B(net884),
    .D(_00108_),
    .Q_N(_06859_),
    .Q(\shift_storage.storage[1004] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1005]$_SDFFE_PN0P_  (.CLK(clknet_leaf_190_clk_p2c),
    .RESET_B(net885),
    .D(_00109_),
    .Q_N(_06858_),
    .Q(\shift_storage.storage[1005] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1006]$_SDFFE_PN0P_  (.CLK(clknet_leaf_190_clk_p2c),
    .RESET_B(net886),
    .D(_00110_),
    .Q_N(_06857_),
    .Q(\shift_storage.storage[1006] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1007]$_SDFFE_PN0P_  (.CLK(clknet_leaf_192_clk_p2c),
    .RESET_B(net887),
    .D(_00111_),
    .Q_N(_06856_),
    .Q(\shift_storage.storage[1007] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1008]$_SDFFE_PN0P_  (.CLK(clknet_leaf_192_clk_p2c),
    .RESET_B(net888),
    .D(_00112_),
    .Q_N(_06855_),
    .Q(\shift_storage.storage[1008] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1009]$_SDFFE_PN0P_  (.CLK(clknet_leaf_191_clk_p2c),
    .RESET_B(net889),
    .D(_00113_),
    .Q_N(_06854_),
    .Q(\shift_storage.storage[1009] ));
 sg13g2_dfrbp_1 \shift_storage.storage[100]$_SDFFE_PN0P_  (.CLK(clknet_leaf_43_clk_p2c),
    .RESET_B(net890),
    .D(_00114_),
    .Q_N(_06853_),
    .Q(\shift_storage.storage[100] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1010]$_SDFFE_PN0P_  (.CLK(clknet_leaf_191_clk_p2c),
    .RESET_B(net891),
    .D(_00115_),
    .Q_N(_06852_),
    .Q(\shift_storage.storage[1010] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1011]$_SDFFE_PN0P_  (.CLK(clknet_leaf_182_clk_p2c),
    .RESET_B(net892),
    .D(_00116_),
    .Q_N(_06851_),
    .Q(\shift_storage.storage[1011] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1012]$_SDFFE_PN0P_  (.CLK(clknet_leaf_182_clk_p2c),
    .RESET_B(net893),
    .D(_00117_),
    .Q_N(_06850_),
    .Q(\shift_storage.storage[1012] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1013]$_SDFFE_PN0P_  (.CLK(clknet_leaf_182_clk_p2c),
    .RESET_B(net894),
    .D(_00118_),
    .Q_N(_06849_),
    .Q(\shift_storage.storage[1013] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1014]$_SDFFE_PN0P_  (.CLK(clknet_leaf_182_clk_p2c),
    .RESET_B(net895),
    .D(_00119_),
    .Q_N(_06848_),
    .Q(\shift_storage.storage[1014] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1015]$_SDFFE_PN0P_  (.CLK(clknet_leaf_180_clk_p2c),
    .RESET_B(net896),
    .D(_00120_),
    .Q_N(_06847_),
    .Q(\shift_storage.storage[1015] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1016]$_SDFFE_PN0P_  (.CLK(clknet_leaf_193_clk_p2c),
    .RESET_B(net897),
    .D(_00121_),
    .Q_N(_06846_),
    .Q(\shift_storage.storage[1016] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1017]$_SDFFE_PN0P_  (.CLK(clknet_leaf_193_clk_p2c),
    .RESET_B(net898),
    .D(_00122_),
    .Q_N(_06845_),
    .Q(\shift_storage.storage[1017] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1018]$_SDFFE_PN0P_  (.CLK(clknet_leaf_192_clk_p2c),
    .RESET_B(net899),
    .D(_00123_),
    .Q_N(_06844_),
    .Q(\shift_storage.storage[1018] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1019]$_SDFFE_PN0P_  (.CLK(clknet_leaf_192_clk_p2c),
    .RESET_B(net900),
    .D(_00124_),
    .Q_N(_06843_),
    .Q(\shift_storage.storage[1019] ));
 sg13g2_dfrbp_1 \shift_storage.storage[101]$_SDFFE_PN0P_  (.CLK(clknet_leaf_43_clk_p2c),
    .RESET_B(net901),
    .D(_00125_),
    .Q_N(_06842_),
    .Q(\shift_storage.storage[101] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1020]$_SDFFE_PN0P_  (.CLK(clknet_leaf_193_clk_p2c),
    .RESET_B(net902),
    .D(_00126_),
    .Q_N(_06841_),
    .Q(\shift_storage.storage[1020] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1021]$_SDFFE_PN0P_  (.CLK(clknet_leaf_194_clk_p2c),
    .RESET_B(net903),
    .D(_00127_),
    .Q_N(_06840_),
    .Q(\shift_storage.storage[1021] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1022]$_SDFFE_PN0P_  (.CLK(clknet_leaf_194_clk_p2c),
    .RESET_B(net904),
    .D(_00128_),
    .Q_N(_06839_),
    .Q(\shift_storage.storage[1022] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1023]$_SDFFE_PN0P_  (.CLK(clknet_leaf_212_clk_p2c),
    .RESET_B(net905),
    .D(_00129_),
    .Q_N(_06838_),
    .Q(\shift_storage.storage[1023] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1024]$_SDFFE_PN0P_  (.CLK(clknet_leaf_213_clk_p2c),
    .RESET_B(net906),
    .D(_00130_),
    .Q_N(_06837_),
    .Q(\shift_storage.storage[1024] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1025]$_SDFFE_PN0P_  (.CLK(clknet_leaf_213_clk_p2c),
    .RESET_B(net907),
    .D(_00131_),
    .Q_N(_06836_),
    .Q(\shift_storage.storage[1025] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1026]$_SDFFE_PN0P_  (.CLK(clknet_leaf_213_clk_p2c),
    .RESET_B(net908),
    .D(_00132_),
    .Q_N(_06835_),
    .Q(\shift_storage.storage[1026] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1027]$_SDFFE_PN0P_  (.CLK(clknet_leaf_231_clk_p2c),
    .RESET_B(net909),
    .D(_00133_),
    .Q_N(_06834_),
    .Q(\shift_storage.storage[1027] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1028]$_SDFFE_PN0P_  (.CLK(clknet_leaf_231_clk_p2c),
    .RESET_B(net910),
    .D(_00134_),
    .Q_N(_06833_),
    .Q(\shift_storage.storage[1028] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1029]$_SDFFE_PN0P_  (.CLK(clknet_leaf_213_clk_p2c),
    .RESET_B(net911),
    .D(_00135_),
    .Q_N(_06832_),
    .Q(\shift_storage.storage[1029] ));
 sg13g2_dfrbp_1 \shift_storage.storage[102]$_SDFFE_PN0P_  (.CLK(clknet_leaf_41_clk_p2c),
    .RESET_B(net912),
    .D(_00136_),
    .Q_N(_06831_),
    .Q(\shift_storage.storage[102] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1030]$_SDFFE_PN0P_  (.CLK(clknet_leaf_213_clk_p2c),
    .RESET_B(net913),
    .D(_00137_),
    .Q_N(_06830_),
    .Q(\shift_storage.storage[1030] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1031]$_SDFFE_PN0P_  (.CLK(clknet_leaf_231_clk_p2c),
    .RESET_B(net914),
    .D(_00138_),
    .Q_N(_06829_),
    .Q(\shift_storage.storage[1031] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1032]$_SDFFE_PN0P_  (.CLK(clknet_leaf_230_clk_p2c),
    .RESET_B(net915),
    .D(_00139_),
    .Q_N(_06828_),
    .Q(\shift_storage.storage[1032] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1033]$_SDFFE_PN0P_  (.CLK(clknet_leaf_231_clk_p2c),
    .RESET_B(net916),
    .D(_00140_),
    .Q_N(_06827_),
    .Q(\shift_storage.storage[1033] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1034]$_SDFFE_PN0P_  (.CLK(clknet_leaf_232_clk_p2c),
    .RESET_B(net917),
    .D(_00141_),
    .Q_N(_06826_),
    .Q(\shift_storage.storage[1034] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1035]$_SDFFE_PN0P_  (.CLK(clknet_leaf_232_clk_p2c),
    .RESET_B(net918),
    .D(_00142_),
    .Q_N(_06825_),
    .Q(\shift_storage.storage[1035] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1036]$_SDFFE_PN0P_  (.CLK(clknet_leaf_232_clk_p2c),
    .RESET_B(net919),
    .D(_00143_),
    .Q_N(_06824_),
    .Q(\shift_storage.storage[1036] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1037]$_SDFFE_PN0P_  (.CLK(clknet_leaf_231_clk_p2c),
    .RESET_B(net920),
    .D(_00144_),
    .Q_N(_06823_),
    .Q(\shift_storage.storage[1037] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1038]$_SDFFE_PN0P_  (.CLK(clknet_leaf_231_clk_p2c),
    .RESET_B(net921),
    .D(_00145_),
    .Q_N(_06822_),
    .Q(\shift_storage.storage[1038] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1039]$_SDFFE_PN0P_  (.CLK(clknet_leaf_179_clk_p2c),
    .RESET_B(net922),
    .D(_00146_),
    .Q_N(_06821_),
    .Q(\shift_storage.storage[1039] ));
 sg13g2_dfrbp_1 \shift_storage.storage[103]$_SDFFE_PN0P_  (.CLK(clknet_leaf_41_clk_p2c),
    .RESET_B(net923),
    .D(_00147_),
    .Q_N(_06820_),
    .Q(\shift_storage.storage[103] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1040]$_SDFFE_PN0P_  (.CLK(clknet_leaf_179_clk_p2c),
    .RESET_B(net924),
    .D(_00148_),
    .Q_N(_06819_),
    .Q(\shift_storage.storage[1040] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1041]$_SDFFE_PN0P_  (.CLK(clknet_leaf_193_clk_p2c),
    .RESET_B(net925),
    .D(_00149_),
    .Q_N(_06818_),
    .Q(\shift_storage.storage[1041] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1042]$_SDFFE_PN0P_  (.CLK(clknet_leaf_193_clk_p2c),
    .RESET_B(net926),
    .D(_00150_),
    .Q_N(_06817_),
    .Q(\shift_storage.storage[1042] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1043]$_SDFFE_PN0P_  (.CLK(clknet_leaf_193_clk_p2c),
    .RESET_B(net927),
    .D(_00151_),
    .Q_N(_06816_),
    .Q(\shift_storage.storage[1043] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1044]$_SDFFE_PN0P_  (.CLK(clknet_leaf_180_clk_p2c),
    .RESET_B(net928),
    .D(_00152_),
    .Q_N(_06815_),
    .Q(\shift_storage.storage[1044] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1045]$_SDFFE_PN0P_  (.CLK(clknet_leaf_180_clk_p2c),
    .RESET_B(net929),
    .D(_00153_),
    .Q_N(_06814_),
    .Q(\shift_storage.storage[1045] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1046]$_SDFFE_PN0P_  (.CLK(clknet_leaf_180_clk_p2c),
    .RESET_B(net930),
    .D(_00154_),
    .Q_N(_06813_),
    .Q(\shift_storage.storage[1046] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1047]$_SDFFE_PN0P_  (.CLK(clknet_leaf_180_clk_p2c),
    .RESET_B(net931),
    .D(_00155_),
    .Q_N(_06812_),
    .Q(\shift_storage.storage[1047] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1048]$_SDFFE_PN0P_  (.CLK(clknet_leaf_181_clk_p2c),
    .RESET_B(net932),
    .D(_00156_),
    .Q_N(_06811_),
    .Q(\shift_storage.storage[1048] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1049]$_SDFFE_PN0P_  (.CLK(clknet_leaf_181_clk_p2c),
    .RESET_B(net933),
    .D(_00157_),
    .Q_N(_06810_),
    .Q(\shift_storage.storage[1049] ));
 sg13g2_dfrbp_1 \shift_storage.storage[104]$_SDFFE_PN0P_  (.CLK(clknet_leaf_41_clk_p2c),
    .RESET_B(net934),
    .D(_00158_),
    .Q_N(_06809_),
    .Q(\shift_storage.storage[104] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1050]$_SDFFE_PN0P_  (.CLK(clknet_leaf_181_clk_p2c),
    .RESET_B(net935),
    .D(_00159_),
    .Q_N(_06808_),
    .Q(\shift_storage.storage[1050] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1051]$_SDFFE_PN0P_  (.CLK(clknet_leaf_183_clk_p2c),
    .RESET_B(net936),
    .D(_00160_),
    .Q_N(_06807_),
    .Q(\shift_storage.storage[1051] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1052]$_SDFFE_PN0P_  (.CLK(clknet_leaf_184_clk_p2c),
    .RESET_B(net937),
    .D(_00161_),
    .Q_N(_06806_),
    .Q(\shift_storage.storage[1052] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1053]$_SDFFE_PN0P_  (.CLK(clknet_leaf_183_clk_p2c),
    .RESET_B(net938),
    .D(_00162_),
    .Q_N(_06805_),
    .Q(\shift_storage.storage[1053] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1054]$_SDFFE_PN0P_  (.CLK(clknet_leaf_183_clk_p2c),
    .RESET_B(net939),
    .D(_00163_),
    .Q_N(_06804_),
    .Q(\shift_storage.storage[1054] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1055]$_SDFFE_PN0P_  (.CLK(clknet_leaf_183_clk_p2c),
    .RESET_B(net940),
    .D(_00164_),
    .Q_N(_06803_),
    .Q(\shift_storage.storage[1055] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1056]$_SDFFE_PN0P_  (.CLK(clknet_leaf_183_clk_p2c),
    .RESET_B(net941),
    .D(_00165_),
    .Q_N(_06802_),
    .Q(\shift_storage.storage[1056] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1057]$_SDFFE_PN0P_  (.CLK(clknet_leaf_186_clk_p2c),
    .RESET_B(net942),
    .D(_00166_),
    .Q_N(_06801_),
    .Q(\shift_storage.storage[1057] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1058]$_SDFFE_PN0P_  (.CLK(clknet_leaf_186_clk_p2c),
    .RESET_B(net943),
    .D(_00167_),
    .Q_N(_06800_),
    .Q(\shift_storage.storage[1058] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1059]$_SDFFE_PN0P_  (.CLK(clknet_leaf_183_clk_p2c),
    .RESET_B(net944),
    .D(_00168_),
    .Q_N(_06799_),
    .Q(\shift_storage.storage[1059] ));
 sg13g2_dfrbp_1 \shift_storage.storage[105]$_SDFFE_PN0P_  (.CLK(clknet_leaf_41_clk_p2c),
    .RESET_B(net945),
    .D(_00169_),
    .Q_N(_06798_),
    .Q(\shift_storage.storage[105] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1060]$_SDFFE_PN0P_  (.CLK(clknet_leaf_182_clk_p2c),
    .RESET_B(net946),
    .D(_00170_),
    .Q_N(_06797_),
    .Q(\shift_storage.storage[1060] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1061]$_SDFFE_PN0P_  (.CLK(clknet_leaf_191_clk_p2c),
    .RESET_B(net947),
    .D(_00171_),
    .Q_N(_06796_),
    .Q(\shift_storage.storage[1061] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1062]$_SDFFE_PN0P_  (.CLK(clknet_leaf_191_clk_p2c),
    .RESET_B(net948),
    .D(_00172_),
    .Q_N(_06795_),
    .Q(\shift_storage.storage[1062] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1063]$_SDFFE_PN0P_  (.CLK(clknet_leaf_191_clk_p2c),
    .RESET_B(net949),
    .D(_00173_),
    .Q_N(_06794_),
    .Q(\shift_storage.storage[1063] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1064]$_SDFFE_PN0P_  (.CLK(clknet_leaf_188_clk_p2c),
    .RESET_B(net950),
    .D(_00174_),
    .Q_N(_06793_),
    .Q(\shift_storage.storage[1064] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1065]$_SDFFE_PN0P_  (.CLK(clknet_leaf_187_clk_p2c),
    .RESET_B(net951),
    .D(_00175_),
    .Q_N(_06792_),
    .Q(\shift_storage.storage[1065] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1066]$_SDFFE_PN0P_  (.CLK(clknet_leaf_187_clk_p2c),
    .RESET_B(net952),
    .D(_00176_),
    .Q_N(_06791_),
    .Q(\shift_storage.storage[1066] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1067]$_SDFFE_PN0P_  (.CLK(clknet_leaf_187_clk_p2c),
    .RESET_B(net953),
    .D(_00177_),
    .Q_N(_06790_),
    .Q(\shift_storage.storage[1067] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1068]$_SDFFE_PN0P_  (.CLK(clknet_leaf_187_clk_p2c),
    .RESET_B(net954),
    .D(_00178_),
    .Q_N(_06789_),
    .Q(\shift_storage.storage[1068] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1069]$_SDFFE_PN0P_  (.CLK(clknet_leaf_187_clk_p2c),
    .RESET_B(net955),
    .D(_00179_),
    .Q_N(_06788_),
    .Q(\shift_storage.storage[1069] ));
 sg13g2_dfrbp_1 \shift_storage.storage[106]$_SDFFE_PN0P_  (.CLK(clknet_leaf_41_clk_p2c),
    .RESET_B(net956),
    .D(_00180_),
    .Q_N(_06787_),
    .Q(\shift_storage.storage[106] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1070]$_SDFFE_PN0P_  (.CLK(clknet_leaf_187_clk_p2c),
    .RESET_B(net957),
    .D(_00181_),
    .Q_N(_06786_),
    .Q(\shift_storage.storage[1070] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1071]$_SDFFE_PN0P_  (.CLK(clknet_leaf_186_clk_p2c),
    .RESET_B(net958),
    .D(_00182_),
    .Q_N(_06785_),
    .Q(\shift_storage.storage[1071] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1072]$_SDFFE_PN0P_  (.CLK(clknet_leaf_186_clk_p2c),
    .RESET_B(net959),
    .D(_00183_),
    .Q_N(_06784_),
    .Q(\shift_storage.storage[1072] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1073]$_SDFFE_PN0P_  (.CLK(clknet_leaf_186_clk_p2c),
    .RESET_B(net960),
    .D(_00184_),
    .Q_N(_06783_),
    .Q(\shift_storage.storage[1073] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1074]$_SDFFE_PN0P_  (.CLK(clknet_leaf_186_clk_p2c),
    .RESET_B(net961),
    .D(_00185_),
    .Q_N(_06782_),
    .Q(\shift_storage.storage[1074] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1075]$_SDFFE_PN0P_  (.CLK(clknet_leaf_183_clk_p2c),
    .RESET_B(net962),
    .D(_00186_),
    .Q_N(_06781_),
    .Q(\shift_storage.storage[1075] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1076]$_SDFFE_PN0P_  (.CLK(clknet_leaf_185_clk_p2c),
    .RESET_B(net963),
    .D(_00187_),
    .Q_N(_06780_),
    .Q(\shift_storage.storage[1076] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1077]$_SDFFE_PN0P_  (.CLK(clknet_leaf_185_clk_p2c),
    .RESET_B(net964),
    .D(_00188_),
    .Q_N(_06779_),
    .Q(\shift_storage.storage[1077] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1078]$_SDFFE_PN0P_  (.CLK(clknet_leaf_185_clk_p2c),
    .RESET_B(net965),
    .D(_00189_),
    .Q_N(_06778_),
    .Q(\shift_storage.storage[1078] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1079]$_SDFFE_PN0P_  (.CLK(clknet_leaf_184_clk_p2c),
    .RESET_B(net966),
    .D(_00190_),
    .Q_N(_06777_),
    .Q(\shift_storage.storage[1079] ));
 sg13g2_dfrbp_1 \shift_storage.storage[107]$_SDFFE_PN0P_  (.CLK(clknet_leaf_31_clk_p2c),
    .RESET_B(net967),
    .D(_00191_),
    .Q_N(_06776_),
    .Q(\shift_storage.storage[107] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1080]$_SDFFE_PN0P_  (.CLK(clknet_leaf_184_clk_p2c),
    .RESET_B(net968),
    .D(_00192_),
    .Q_N(_06775_),
    .Q(\shift_storage.storage[1080] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1081]$_SDFFE_PN0P_  (.CLK(clknet_leaf_184_clk_p2c),
    .RESET_B(net969),
    .D(_00193_),
    .Q_N(_06774_),
    .Q(\shift_storage.storage[1081] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1082]$_SDFFE_PN0P_  (.CLK(clknet_leaf_184_clk_p2c),
    .RESET_B(net970),
    .D(_00194_),
    .Q_N(_06773_),
    .Q(\shift_storage.storage[1082] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1083]$_SDFFE_PN0P_  (.CLK(clknet_leaf_184_clk_p2c),
    .RESET_B(net971),
    .D(_00195_),
    .Q_N(_06772_),
    .Q(\shift_storage.storage[1083] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1084]$_SDFFE_PN0P_  (.CLK(clknet_leaf_181_clk_p2c),
    .RESET_B(net972),
    .D(_00196_),
    .Q_N(_06771_),
    .Q(\shift_storage.storage[1084] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1085]$_SDFFE_PN0P_  (.CLK(clknet_leaf_181_clk_p2c),
    .RESET_B(net973),
    .D(_00197_),
    .Q_N(_06770_),
    .Q(\shift_storage.storage[1085] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1086]$_SDFFE_PN0P_  (.CLK(clknet_leaf_178_clk_p2c),
    .RESET_B(net974),
    .D(_00198_),
    .Q_N(_06769_),
    .Q(\shift_storage.storage[1086] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1087]$_SDFFE_PN0P_  (.CLK(clknet_leaf_178_clk_p2c),
    .RESET_B(net975),
    .D(_00199_),
    .Q_N(_06768_),
    .Q(\shift_storage.storage[1087] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1088]$_SDFFE_PN0P_  (.CLK(clknet_leaf_178_clk_p2c),
    .RESET_B(net976),
    .D(_00200_),
    .Q_N(_06767_),
    .Q(\shift_storage.storage[1088] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1089]$_SDFFE_PN0P_  (.CLK(clknet_leaf_179_clk_p2c),
    .RESET_B(net977),
    .D(_00201_),
    .Q_N(_06766_),
    .Q(\shift_storage.storage[1089] ));
 sg13g2_dfrbp_1 \shift_storage.storage[108]$_SDFFE_PN0P_  (.CLK(clknet_leaf_31_clk_p2c),
    .RESET_B(net978),
    .D(_00202_),
    .Q_N(_06765_),
    .Q(\shift_storage.storage[108] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1090]$_SDFFE_PN0P_  (.CLK(clknet_leaf_180_clk_p2c),
    .RESET_B(net979),
    .D(_00203_),
    .Q_N(_06764_),
    .Q(\shift_storage.storage[1090] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1091]$_SDFFE_PN0P_  (.CLK(clknet_leaf_179_clk_p2c),
    .RESET_B(net980),
    .D(_00204_),
    .Q_N(_06763_),
    .Q(\shift_storage.storage[1091] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1092]$_SDFFE_PN0P_  (.CLK(clknet_leaf_179_clk_p2c),
    .RESET_B(net981),
    .D(_00205_),
    .Q_N(_06762_),
    .Q(\shift_storage.storage[1092] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1093]$_SDFFE_PN0P_  (.CLK(clknet_leaf_232_clk_p2c),
    .RESET_B(net982),
    .D(_00206_),
    .Q_N(_06761_),
    .Q(\shift_storage.storage[1093] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1094]$_SDFFE_PN0P_  (.CLK(clknet_leaf_179_clk_p2c),
    .RESET_B(net983),
    .D(_00207_),
    .Q_N(_06760_),
    .Q(\shift_storage.storage[1094] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1095]$_SDFFE_PN0P_  (.CLK(clknet_leaf_178_clk_p2c),
    .RESET_B(net984),
    .D(_00208_),
    .Q_N(_06759_),
    .Q(\shift_storage.storage[1095] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1096]$_SDFFE_PN0P_  (.CLK(clknet_leaf_178_clk_p2c),
    .RESET_B(net985),
    .D(_00209_),
    .Q_N(_06758_),
    .Q(\shift_storage.storage[1096] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1097]$_SDFFE_PN0P_  (.CLK(clknet_leaf_177_clk_p2c),
    .RESET_B(net986),
    .D(_00210_),
    .Q_N(_06757_),
    .Q(\shift_storage.storage[1097] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1098]$_SDFFE_PN0P_  (.CLK(clknet_leaf_177_clk_p2c),
    .RESET_B(net987),
    .D(_00211_),
    .Q_N(_06756_),
    .Q(\shift_storage.storage[1098] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1099]$_SDFFE_PN0P_  (.CLK(clknet_leaf_177_clk_p2c),
    .RESET_B(net988),
    .D(_00212_),
    .Q_N(_06755_),
    .Q(\shift_storage.storage[1099] ));
 sg13g2_dfrbp_1 \shift_storage.storage[109]$_SDFFE_PN0P_  (.CLK(clknet_leaf_31_clk_p2c),
    .RESET_B(net989),
    .D(_00213_),
    .Q_N(_06754_),
    .Q(\shift_storage.storage[109] ));
 sg13g2_dfrbp_1 \shift_storage.storage[10]$_SDFFE_PN0P_  (.CLK(clknet_leaf_70_clk_p2c),
    .RESET_B(net990),
    .D(_00214_),
    .Q_N(_06753_),
    .Q(\shift_storage.storage[10] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1100]$_SDFFE_PN0P_  (.CLK(clknet_leaf_177_clk_p2c),
    .RESET_B(net991),
    .D(_00215_),
    .Q_N(_06752_),
    .Q(\shift_storage.storage[1100] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1101]$_SDFFE_PN0P_  (.CLK(clknet_leaf_233_clk_p2c),
    .RESET_B(net992),
    .D(_00216_),
    .Q_N(_06751_),
    .Q(\shift_storage.storage[1101] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1102]$_SDFFE_PN0P_  (.CLK(clknet_leaf_233_clk_p2c),
    .RESET_B(net993),
    .D(_00217_),
    .Q_N(_06750_),
    .Q(\shift_storage.storage[1102] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1103]$_SDFFE_PN0P_  (.CLK(clknet_leaf_233_clk_p2c),
    .RESET_B(net994),
    .D(_00218_),
    .Q_N(_06749_),
    .Q(\shift_storage.storage[1103] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1104]$_SDFFE_PN0P_  (.CLK(clknet_leaf_233_clk_p2c),
    .RESET_B(net995),
    .D(_00219_),
    .Q_N(_06748_),
    .Q(\shift_storage.storage[1104] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1105]$_SDFFE_PN0P_  (.CLK(clknet_leaf_235_clk_p2c),
    .RESET_B(net996),
    .D(_00220_),
    .Q_N(_06747_),
    .Q(\shift_storage.storage[1105] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1106]$_SDFFE_PN0P_  (.CLK(clknet_leaf_235_clk_p2c),
    .RESET_B(net997),
    .D(_00221_),
    .Q_N(_06746_),
    .Q(\shift_storage.storage[1106] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1107]$_SDFFE_PN0P_  (.CLK(clknet_leaf_235_clk_p2c),
    .RESET_B(net998),
    .D(_00222_),
    .Q_N(_06745_),
    .Q(\shift_storage.storage[1107] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1108]$_SDFFE_PN0P_  (.CLK(clknet_leaf_235_clk_p2c),
    .RESET_B(net999),
    .D(_00223_),
    .Q_N(_06744_),
    .Q(\shift_storage.storage[1108] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1109]$_SDFFE_PN0P_  (.CLK(clknet_leaf_235_clk_p2c),
    .RESET_B(net1000),
    .D(_00224_),
    .Q_N(_06743_),
    .Q(\shift_storage.storage[1109] ));
 sg13g2_dfrbp_1 \shift_storage.storage[110]$_SDFFE_PN0P_  (.CLK(clknet_leaf_32_clk_p2c),
    .RESET_B(net1001),
    .D(_00225_),
    .Q_N(_06742_),
    .Q(\shift_storage.storage[110] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1110]$_SDFFE_PN0P_  (.CLK(clknet_leaf_240_clk_p2c),
    .RESET_B(net1002),
    .D(_00226_),
    .Q_N(_06741_),
    .Q(\shift_storage.storage[1110] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1111]$_SDFFE_PN0P_  (.CLK(clknet_leaf_240_clk_p2c),
    .RESET_B(net1003),
    .D(_00227_),
    .Q_N(_06740_),
    .Q(\shift_storage.storage[1111] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1112]$_SDFFE_PN0P_  (.CLK(clknet_leaf_240_clk_p2c),
    .RESET_B(net1004),
    .D(_00228_),
    .Q_N(_06739_),
    .Q(\shift_storage.storage[1112] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1113]$_SDFFE_PN0P_  (.CLK(clknet_leaf_239_clk_p2c),
    .RESET_B(net1005),
    .D(_00229_),
    .Q_N(_06738_),
    .Q(\shift_storage.storage[1113] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1114]$_SDFFE_PN0P_  (.CLK(clknet_leaf_238_clk_p2c),
    .RESET_B(net1006),
    .D(_00230_),
    .Q_N(_06737_),
    .Q(\shift_storage.storage[1114] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1115]$_SDFFE_PN0P_  (.CLK(clknet_leaf_239_clk_p2c),
    .RESET_B(net1007),
    .D(_00231_),
    .Q_N(_06736_),
    .Q(\shift_storage.storage[1115] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1116]$_SDFFE_PN0P_  (.CLK(clknet_leaf_239_clk_p2c),
    .RESET_B(net1008),
    .D(_00232_),
    .Q_N(_06735_),
    .Q(\shift_storage.storage[1116] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1117]$_SDFFE_PN0P_  (.CLK(clknet_leaf_239_clk_p2c),
    .RESET_B(net1009),
    .D(_00233_),
    .Q_N(_06734_),
    .Q(\shift_storage.storage[1117] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1118]$_SDFFE_PN0P_  (.CLK(clknet_leaf_239_clk_p2c),
    .RESET_B(net1010),
    .D(_00234_),
    .Q_N(_06733_),
    .Q(\shift_storage.storage[1118] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1119]$_SDFFE_PN0P_  (.CLK(clknet_leaf_241_clk_p2c),
    .RESET_B(net1011),
    .D(_00235_),
    .Q_N(_06732_),
    .Q(\shift_storage.storage[1119] ));
 sg13g2_dfrbp_1 \shift_storage.storage[111]$_SDFFE_PN0P_  (.CLK(clknet_leaf_40_clk_p2c),
    .RESET_B(net1012),
    .D(_00236_),
    .Q_N(_06731_),
    .Q(\shift_storage.storage[111] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1120]$_SDFFE_PN0P_  (.CLK(clknet_leaf_240_clk_p2c),
    .RESET_B(net1013),
    .D(_00237_),
    .Q_N(_06730_),
    .Q(\shift_storage.storage[1120] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1121]$_SDFFE_PN0P_  (.CLK(clknet_leaf_240_clk_p2c),
    .RESET_B(net1014),
    .D(_00238_),
    .Q_N(_06729_),
    .Q(\shift_storage.storage[1121] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1122]$_SDFFE_PN0P_  (.CLK(clknet_leaf_240_clk_p2c),
    .RESET_B(net1015),
    .D(_00239_),
    .Q_N(_06728_),
    .Q(\shift_storage.storage[1122] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1123]$_SDFFE_PN0P_  (.CLK(clknet_leaf_234_clk_p2c),
    .RESET_B(net1016),
    .D(_00240_),
    .Q_N(_06727_),
    .Q(\shift_storage.storage[1123] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1124]$_SDFFE_PN0P_  (.CLK(clknet_leaf_234_clk_p2c),
    .RESET_B(net1017),
    .D(_00241_),
    .Q_N(_06726_),
    .Q(\shift_storage.storage[1124] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1125]$_SDFFE_PN0P_  (.CLK(clknet_leaf_234_clk_p2c),
    .RESET_B(net1018),
    .D(_00242_),
    .Q_N(_06725_),
    .Q(\shift_storage.storage[1125] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1126]$_SDFFE_PN0P_  (.CLK(clknet_leaf_234_clk_p2c),
    .RESET_B(net1019),
    .D(_00243_),
    .Q_N(_06724_),
    .Q(\shift_storage.storage[1126] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1127]$_SDFFE_PN0P_  (.CLK(clknet_leaf_176_clk_p2c),
    .RESET_B(net1020),
    .D(_00244_),
    .Q_N(_06723_),
    .Q(\shift_storage.storage[1127] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1128]$_SDFFE_PN0P_  (.CLK(clknet_leaf_177_clk_p2c),
    .RESET_B(net1021),
    .D(_00245_),
    .Q_N(_06722_),
    .Q(\shift_storage.storage[1128] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1129]$_SDFFE_PN0P_  (.CLK(clknet_leaf_176_clk_p2c),
    .RESET_B(net1022),
    .D(_00246_),
    .Q_N(_06721_),
    .Q(\shift_storage.storage[1129] ));
 sg13g2_dfrbp_1 \shift_storage.storage[112]$_SDFFE_PN0P_  (.CLK(clknet_leaf_32_clk_p2c),
    .RESET_B(net1023),
    .D(_00247_),
    .Q_N(_06720_),
    .Q(\shift_storage.storage[112] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1130]$_SDFFE_PN0P_  (.CLK(clknet_leaf_175_clk_p2c),
    .RESET_B(net1024),
    .D(_00248_),
    .Q_N(_06719_),
    .Q(\shift_storage.storage[1130] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1131]$_SDFFE_PN0P_  (.CLK(clknet_leaf_175_clk_p2c),
    .RESET_B(net1025),
    .D(_00249_),
    .Q_N(_06718_),
    .Q(\shift_storage.storage[1131] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1132]$_SDFFE_PN0P_  (.CLK(clknet_leaf_177_clk_p2c),
    .RESET_B(net1026),
    .D(_00250_),
    .Q_N(_06717_),
    .Q(\shift_storage.storage[1132] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1133]$_SDFFE_PN0P_  (.CLK(clknet_leaf_177_clk_p2c),
    .RESET_B(net1027),
    .D(_00251_),
    .Q_N(_06716_),
    .Q(\shift_storage.storage[1133] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1134]$_SDFFE_PN0P_  (.CLK(clknet_leaf_178_clk_p2c),
    .RESET_B(net1028),
    .D(_00252_),
    .Q_N(_06715_),
    .Q(\shift_storage.storage[1134] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1135]$_SDFFE_PN0P_  (.CLK(clknet_leaf_175_clk_p2c),
    .RESET_B(net1029),
    .D(_00253_),
    .Q_N(_06714_),
    .Q(\shift_storage.storage[1135] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1136]$_SDFFE_PN0P_  (.CLK(clknet_leaf_175_clk_p2c),
    .RESET_B(net1030),
    .D(_00254_),
    .Q_N(_06713_),
    .Q(\shift_storage.storage[1136] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1137]$_SDFFE_PN0P_  (.CLK(clknet_leaf_175_clk_p2c),
    .RESET_B(net1031),
    .D(_00255_),
    .Q_N(_06712_),
    .Q(\shift_storage.storage[1137] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1138]$_SDFFE_PN0P_  (.CLK(clknet_leaf_174_clk_p2c),
    .RESET_B(net1032),
    .D(_00256_),
    .Q_N(_06711_),
    .Q(\shift_storage.storage[1138] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1139]$_SDFFE_PN0P_  (.CLK(clknet_leaf_174_clk_p2c),
    .RESET_B(net1033),
    .D(_00257_),
    .Q_N(_06710_),
    .Q(\shift_storage.storage[1139] ));
 sg13g2_dfrbp_1 \shift_storage.storage[113]$_SDFFE_PN0P_  (.CLK(clknet_leaf_40_clk_p2c),
    .RESET_B(net1034),
    .D(_00258_),
    .Q_N(_06709_),
    .Q(\shift_storage.storage[113] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1140]$_SDFFE_PN0P_  (.CLK(clknet_leaf_174_clk_p2c),
    .RESET_B(net1035),
    .D(_00259_),
    .Q_N(_06708_),
    .Q(\shift_storage.storage[1140] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1141]$_SDFFE_PN0P_  (.CLK(clknet_leaf_174_clk_p2c),
    .RESET_B(net1036),
    .D(_00260_),
    .Q_N(_06707_),
    .Q(\shift_storage.storage[1141] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1142]$_SDFFE_PN0P_  (.CLK(clknet_leaf_174_clk_p2c),
    .RESET_B(net1037),
    .D(_00261_),
    .Q_N(_06706_),
    .Q(\shift_storage.storage[1142] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1143]$_SDFFE_PN0P_  (.CLK(clknet_leaf_185_clk_p2c),
    .RESET_B(net1038),
    .D(_00262_),
    .Q_N(_06705_),
    .Q(\shift_storage.storage[1143] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1144]$_SDFFE_PN0P_  (.CLK(clknet_leaf_185_clk_p2c),
    .RESET_B(net1039),
    .D(_00263_),
    .Q_N(_06704_),
    .Q(\shift_storage.storage[1144] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1145]$_SDFFE_PN0P_  (.CLK(clknet_leaf_173_clk_p2c),
    .RESET_B(net1040),
    .D(_00264_),
    .Q_N(_06703_),
    .Q(\shift_storage.storage[1145] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1146]$_SDFFE_PN0P_  (.CLK(clknet_leaf_173_clk_p2c),
    .RESET_B(net1041),
    .D(_00265_),
    .Q_N(_06702_),
    .Q(\shift_storage.storage[1146] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1147]$_SDFFE_PN0P_  (.CLK(clknet_leaf_151_clk_p2c),
    .RESET_B(net1042),
    .D(_00266_),
    .Q_N(_06701_),
    .Q(\shift_storage.storage[1147] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1148]$_SDFFE_PN0P_  (.CLK(clknet_leaf_151_clk_p2c),
    .RESET_B(net1043),
    .D(_00267_),
    .Q_N(_06700_),
    .Q(\shift_storage.storage[1148] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1149]$_SDFFE_PN0P_  (.CLK(clknet_leaf_151_clk_p2c),
    .RESET_B(net1044),
    .D(_00268_),
    .Q_N(_06699_),
    .Q(\shift_storage.storage[1149] ));
 sg13g2_dfrbp_1 \shift_storage.storage[114]$_SDFFE_PN0P_  (.CLK(clknet_leaf_34_clk_p2c),
    .RESET_B(net1045),
    .D(_00269_),
    .Q_N(_06698_),
    .Q(\shift_storage.storage[114] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1150]$_SDFFE_PN0P_  (.CLK(clknet_leaf_150_clk_p2c),
    .RESET_B(net1046),
    .D(_00270_),
    .Q_N(_06697_),
    .Q(\shift_storage.storage[1150] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1151]$_SDFFE_PN0P_  (.CLK(clknet_leaf_150_clk_p2c),
    .RESET_B(net1047),
    .D(_00271_),
    .Q_N(_06696_),
    .Q(\shift_storage.storage[1151] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1152]$_SDFFE_PN0P_  (.CLK(clknet_leaf_150_clk_p2c),
    .RESET_B(net1048),
    .D(_00272_),
    .Q_N(_06695_),
    .Q(\shift_storage.storage[1152] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1153]$_SDFFE_PN0P_  (.CLK(clknet_leaf_150_clk_p2c),
    .RESET_B(net1049),
    .D(_00273_),
    .Q_N(_06694_),
    .Q(\shift_storage.storage[1153] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1154]$_SDFFE_PN0P_  (.CLK(clknet_leaf_150_clk_p2c),
    .RESET_B(net1050),
    .D(_00274_),
    .Q_N(_06693_),
    .Q(\shift_storage.storage[1154] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1155]$_SDFFE_PN0P_  (.CLK(clknet_leaf_149_clk_p2c),
    .RESET_B(net1051),
    .D(_00275_),
    .Q_N(_06692_),
    .Q(\shift_storage.storage[1155] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1156]$_SDFFE_PN0P_  (.CLK(clknet_leaf_150_clk_p2c),
    .RESET_B(net1052),
    .D(_00276_),
    .Q_N(_06691_),
    .Q(\shift_storage.storage[1156] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1157]$_SDFFE_PN0P_  (.CLK(clknet_leaf_149_clk_p2c),
    .RESET_B(net1053),
    .D(_00277_),
    .Q_N(_06690_),
    .Q(\shift_storage.storage[1157] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1158]$_SDFFE_PN0P_  (.CLK(clknet_leaf_149_clk_p2c),
    .RESET_B(net1054),
    .D(_00278_),
    .Q_N(_06689_),
    .Q(\shift_storage.storage[1158] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1159]$_SDFFE_PN0P_  (.CLK(clknet_leaf_148_clk_p2c),
    .RESET_B(net1055),
    .D(_00279_),
    .Q_N(_06688_),
    .Q(\shift_storage.storage[1159] ));
 sg13g2_dfrbp_1 \shift_storage.storage[115]$_SDFFE_PN0P_  (.CLK(clknet_leaf_34_clk_p2c),
    .RESET_B(net1056),
    .D(_00280_),
    .Q_N(_06687_),
    .Q(\shift_storage.storage[115] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1160]$_SDFFE_PN0P_  (.CLK(clknet_leaf_149_clk_p2c),
    .RESET_B(net1057),
    .D(_00281_),
    .Q_N(_06686_),
    .Q(\shift_storage.storage[1160] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1161]$_SDFFE_PN0P_  (.CLK(clknet_leaf_148_clk_p2c),
    .RESET_B(net1058),
    .D(_00282_),
    .Q_N(_06685_),
    .Q(\shift_storage.storage[1161] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1162]$_SDFFE_PN0P_  (.CLK(clknet_leaf_147_clk_p2c),
    .RESET_B(net1059),
    .D(_00283_),
    .Q_N(_06684_),
    .Q(\shift_storage.storage[1162] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1163]$_SDFFE_PN0P_  (.CLK(clknet_leaf_147_clk_p2c),
    .RESET_B(net1060),
    .D(_00284_),
    .Q_N(_06683_),
    .Q(\shift_storage.storage[1163] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1164]$_SDFFE_PN0P_  (.CLK(clknet_leaf_147_clk_p2c),
    .RESET_B(net1061),
    .D(_00285_),
    .Q_N(_06682_),
    .Q(\shift_storage.storage[1164] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1165]$_SDFFE_PN0P_  (.CLK(clknet_leaf_147_clk_p2c),
    .RESET_B(net1062),
    .D(_00286_),
    .Q_N(_06681_),
    .Q(\shift_storage.storage[1165] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1166]$_SDFFE_PN0P_  (.CLK(clknet_leaf_148_clk_p2c),
    .RESET_B(net1063),
    .D(_00287_),
    .Q_N(_06680_),
    .Q(\shift_storage.storage[1166] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1167]$_SDFFE_PN0P_  (.CLK(clknet_leaf_148_clk_p2c),
    .RESET_B(net1064),
    .D(_00288_),
    .Q_N(_06679_),
    .Q(\shift_storage.storage[1167] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1168]$_SDFFE_PN0P_  (.CLK(clknet_leaf_148_clk_p2c),
    .RESET_B(net1065),
    .D(_00289_),
    .Q_N(_06678_),
    .Q(\shift_storage.storage[1168] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1169]$_SDFFE_PN0P_  (.CLK(clknet_leaf_154_clk_p2c),
    .RESET_B(net1066),
    .D(_00290_),
    .Q_N(_06677_),
    .Q(\shift_storage.storage[1169] ));
 sg13g2_dfrbp_1 \shift_storage.storage[116]$_SDFFE_PN0P_  (.CLK(clknet_leaf_35_clk_p2c),
    .RESET_B(net1067),
    .D(_00291_),
    .Q_N(_06676_),
    .Q(\shift_storage.storage[116] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1170]$_SDFFE_PN0P_  (.CLK(clknet_leaf_148_clk_p2c),
    .RESET_B(net1068),
    .D(_00292_),
    .Q_N(_06675_),
    .Q(\shift_storage.storage[1170] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1171]$_SDFFE_PN0P_  (.CLK(clknet_leaf_149_clk_p2c),
    .RESET_B(net1069),
    .D(_00293_),
    .Q_N(_06674_),
    .Q(\shift_storage.storage[1171] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1172]$_SDFFE_PN0P_  (.CLK(clknet_leaf_154_clk_p2c),
    .RESET_B(net1070),
    .D(_00294_),
    .Q_N(_06673_),
    .Q(\shift_storage.storage[1172] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1173]$_SDFFE_PN0P_  (.CLK(clknet_leaf_153_clk_p2c),
    .RESET_B(net1071),
    .D(_00295_),
    .Q_N(_06672_),
    .Q(\shift_storage.storage[1173] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1174]$_SDFFE_PN0P_  (.CLK(clknet_leaf_153_clk_p2c),
    .RESET_B(net1072),
    .D(_00296_),
    .Q_N(_06671_),
    .Q(\shift_storage.storage[1174] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1175]$_SDFFE_PN0P_  (.CLK(clknet_leaf_152_clk_p2c),
    .RESET_B(net1073),
    .D(_00297_),
    .Q_N(_06670_),
    .Q(\shift_storage.storage[1175] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1176]$_SDFFE_PN0P_  (.CLK(clknet_leaf_152_clk_p2c),
    .RESET_B(net1074),
    .D(_00298_),
    .Q_N(_06669_),
    .Q(\shift_storage.storage[1176] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1177]$_SDFFE_PN0P_  (.CLK(clknet_leaf_152_clk_p2c),
    .RESET_B(net1075),
    .D(_00299_),
    .Q_N(_06668_),
    .Q(\shift_storage.storage[1177] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1178]$_SDFFE_PN0P_  (.CLK(clknet_leaf_152_clk_p2c),
    .RESET_B(net1076),
    .D(_00300_),
    .Q_N(_06667_),
    .Q(\shift_storage.storage[1178] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1179]$_SDFFE_PN0P_  (.CLK(clknet_leaf_150_clk_p2c),
    .RESET_B(net1077),
    .D(_00301_),
    .Q_N(_06666_),
    .Q(\shift_storage.storage[1179] ));
 sg13g2_dfrbp_1 \shift_storage.storage[117]$_SDFFE_PN0P_  (.CLK(clknet_leaf_35_clk_p2c),
    .RESET_B(net1078),
    .D(_00302_),
    .Q_N(_06665_),
    .Q(\shift_storage.storage[117] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1180]$_SDFFE_PN0P_  (.CLK(clknet_leaf_151_clk_p2c),
    .RESET_B(net1079),
    .D(_00303_),
    .Q_N(_06664_),
    .Q(\shift_storage.storage[1180] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1181]$_SDFFE_PN0P_  (.CLK(clknet_leaf_151_clk_p2c),
    .RESET_B(net1080),
    .D(_00304_),
    .Q_N(_06663_),
    .Q(\shift_storage.storage[1181] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1182]$_SDFFE_PN0P_  (.CLK(clknet_leaf_152_clk_p2c),
    .RESET_B(net1081),
    .D(_00305_),
    .Q_N(_06662_),
    .Q(\shift_storage.storage[1182] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1183]$_SDFFE_PN0P_  (.CLK(clknet_leaf_162_clk_p2c),
    .RESET_B(net1082),
    .D(_00306_),
    .Q_N(_06661_),
    .Q(\shift_storage.storage[1183] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1184]$_SDFFE_PN0P_  (.CLK(clknet_leaf_162_clk_p2c),
    .RESET_B(net1083),
    .D(_00307_),
    .Q_N(_06660_),
    .Q(\shift_storage.storage[1184] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1185]$_SDFFE_PN0P_  (.CLK(clknet_leaf_151_clk_p2c),
    .RESET_B(net1084),
    .D(_00308_),
    .Q_N(_06659_),
    .Q(\shift_storage.storage[1185] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1186]$_SDFFE_PN0P_  (.CLK(clknet_leaf_162_clk_p2c),
    .RESET_B(net1085),
    .D(_00309_),
    .Q_N(_06658_),
    .Q(\shift_storage.storage[1186] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1187]$_SDFFE_PN0P_  (.CLK(clknet_leaf_162_clk_p2c),
    .RESET_B(net1086),
    .D(_00310_),
    .Q_N(_06657_),
    .Q(\shift_storage.storage[1187] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1188]$_SDFFE_PN0P_  (.CLK(clknet_leaf_163_clk_p2c),
    .RESET_B(net1087),
    .D(_00311_),
    .Q_N(_06656_),
    .Q(\shift_storage.storage[1188] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1189]$_SDFFE_PN0P_  (.CLK(clknet_leaf_163_clk_p2c),
    .RESET_B(net1088),
    .D(_00312_),
    .Q_N(_06655_),
    .Q(\shift_storage.storage[1189] ));
 sg13g2_dfrbp_1 \shift_storage.storage[118]$_SDFFE_PN0P_  (.CLK(clknet_leaf_35_clk_p2c),
    .RESET_B(net1089),
    .D(_00313_),
    .Q_N(_06654_),
    .Q(\shift_storage.storage[118] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1190]$_SDFFE_PN0P_  (.CLK(clknet_leaf_173_clk_p2c),
    .RESET_B(net1090),
    .D(_00314_),
    .Q_N(_06653_),
    .Q(\shift_storage.storage[1190] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1191]$_SDFFE_PN0P_  (.CLK(clknet_leaf_173_clk_p2c),
    .RESET_B(net1091),
    .D(_00315_),
    .Q_N(_06652_),
    .Q(\shift_storage.storage[1191] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1192]$_SDFFE_PN0P_  (.CLK(clknet_leaf_173_clk_p2c),
    .RESET_B(net1092),
    .D(_00316_),
    .Q_N(_06651_),
    .Q(\shift_storage.storage[1192] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1193]$_SDFFE_PN0P_  (.CLK(clknet_leaf_173_clk_p2c),
    .RESET_B(net1093),
    .D(_00317_),
    .Q_N(_06650_),
    .Q(\shift_storage.storage[1193] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1194]$_SDFFE_PN0P_  (.CLK(clknet_leaf_174_clk_p2c),
    .RESET_B(net1094),
    .D(_00318_),
    .Q_N(_06649_),
    .Q(\shift_storage.storage[1194] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1195]$_SDFFE_PN0P_  (.CLK(clknet_leaf_174_clk_p2c),
    .RESET_B(net1095),
    .D(_00319_),
    .Q_N(_06648_),
    .Q(\shift_storage.storage[1195] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1196]$_SDFFE_PN0P_  (.CLK(clknet_leaf_176_clk_p2c),
    .RESET_B(net1096),
    .D(_00320_),
    .Q_N(_06647_),
    .Q(\shift_storage.storage[1196] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1197]$_SDFFE_PN0P_  (.CLK(clknet_leaf_176_clk_p2c),
    .RESET_B(net1097),
    .D(_00321_),
    .Q_N(_06646_),
    .Q(\shift_storage.storage[1197] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1198]$_SDFFE_PN0P_  (.CLK(clknet_leaf_176_clk_p2c),
    .RESET_B(net1098),
    .D(_00322_),
    .Q_N(_06645_),
    .Q(\shift_storage.storage[1198] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1199]$_SDFFE_PN0P_  (.CLK(clknet_leaf_171_clk_p2c),
    .RESET_B(net1099),
    .D(_00323_),
    .Q_N(_06644_),
    .Q(\shift_storage.storage[1199] ));
 sg13g2_dfrbp_1 \shift_storage.storage[119]$_SDFFE_PN0P_  (.CLK(clknet_leaf_35_clk_p2c),
    .RESET_B(net1100),
    .D(_00324_),
    .Q_N(_06643_),
    .Q(\shift_storage.storage[119] ));
 sg13g2_dfrbp_1 \shift_storage.storage[11]$_SDFFE_PN0P_  (.CLK(clknet_leaf_70_clk_p2c),
    .RESET_B(net1101),
    .D(_00325_),
    .Q_N(_06642_),
    .Q(\shift_storage.storage[11] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1200]$_SDFFE_PN0P_  (.CLK(clknet_leaf_176_clk_p2c),
    .RESET_B(net1102),
    .D(_00326_),
    .Q_N(_06641_),
    .Q(\shift_storage.storage[1200] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1201]$_SDFFE_PN0P_  (.CLK(clknet_leaf_176_clk_p2c),
    .RESET_B(net1103),
    .D(_00327_),
    .Q_N(_06640_),
    .Q(\shift_storage.storage[1201] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1202]$_SDFFE_PN0P_  (.CLK(clknet_leaf_241_clk_p2c),
    .RESET_B(net1104),
    .D(_00328_),
    .Q_N(_06639_),
    .Q(\shift_storage.storage[1202] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1203]$_SDFFE_PN0P_  (.CLK(clknet_leaf_241_clk_p2c),
    .RESET_B(net1105),
    .D(_00329_),
    .Q_N(_06638_),
    .Q(\shift_storage.storage[1203] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1204]$_SDFFE_PN0P_  (.CLK(clknet_leaf_241_clk_p2c),
    .RESET_B(net1106),
    .D(_00330_),
    .Q_N(_06637_),
    .Q(\shift_storage.storage[1204] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1205]$_SDFFE_PN0P_  (.CLK(clknet_leaf_171_clk_p2c),
    .RESET_B(net1107),
    .D(_00331_),
    .Q_N(_06636_),
    .Q(\shift_storage.storage[1205] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1206]$_SDFFE_PN0P_  (.CLK(clknet_leaf_171_clk_p2c),
    .RESET_B(net1108),
    .D(_00332_),
    .Q_N(_06635_),
    .Q(\shift_storage.storage[1206] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1207]$_SDFFE_PN0P_  (.CLK(clknet_leaf_170_clk_p2c),
    .RESET_B(net1109),
    .D(_00333_),
    .Q_N(_06634_),
    .Q(\shift_storage.storage[1207] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1208]$_SDFFE_PN0P_  (.CLK(clknet_leaf_170_clk_p2c),
    .RESET_B(net1110),
    .D(_00334_),
    .Q_N(_06633_),
    .Q(\shift_storage.storage[1208] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1209]$_SDFFE_PN0P_  (.CLK(clknet_leaf_169_clk_p2c),
    .RESET_B(net1111),
    .D(_00335_),
    .Q_N(_06632_),
    .Q(\shift_storage.storage[1209] ));
 sg13g2_dfrbp_1 \shift_storage.storage[120]$_SDFFE_PN0P_  (.CLK(clknet_leaf_36_clk_p2c),
    .RESET_B(net1112),
    .D(_00336_),
    .Q_N(_06631_),
    .Q(\shift_storage.storage[120] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1210]$_SDFFE_PN0P_  (.CLK(clknet_leaf_169_clk_p2c),
    .RESET_B(net1113),
    .D(_00337_),
    .Q_N(_06630_),
    .Q(\shift_storage.storage[1210] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1211]$_SDFFE_PN0P_  (.CLK(clknet_leaf_169_clk_p2c),
    .RESET_B(net1114),
    .D(_00338_),
    .Q_N(_06629_),
    .Q(\shift_storage.storage[1211] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1212]$_SDFFE_PN0P_  (.CLK(clknet_leaf_167_clk_p2c),
    .RESET_B(net1115),
    .D(_00339_),
    .Q_N(_06628_),
    .Q(\shift_storage.storage[1212] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1213]$_SDFFE_PN0P_  (.CLK(clknet_leaf_167_clk_p2c),
    .RESET_B(net1116),
    .D(_00340_),
    .Q_N(_06627_),
    .Q(\shift_storage.storage[1213] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1214]$_SDFFE_PN0P_  (.CLK(clknet_leaf_170_clk_p2c),
    .RESET_B(net1117),
    .D(_00341_),
    .Q_N(_06626_),
    .Q(\shift_storage.storage[1214] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1215]$_SDFFE_PN0P_  (.CLK(clknet_leaf_170_clk_p2c),
    .RESET_B(net1118),
    .D(_00342_),
    .Q_N(_06625_),
    .Q(\shift_storage.storage[1215] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1216]$_SDFFE_PN0P_  (.CLK(clknet_leaf_172_clk_p2c),
    .RESET_B(net1119),
    .D(_00343_),
    .Q_N(_06624_),
    .Q(\shift_storage.storage[1216] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1217]$_SDFFE_PN0P_  (.CLK(clknet_leaf_164_clk_p2c),
    .RESET_B(net1120),
    .D(_00344_),
    .Q_N(_06623_),
    .Q(\shift_storage.storage[1217] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1218]$_SDFFE_PN0P_  (.CLK(clknet_leaf_164_clk_p2c),
    .RESET_B(net1121),
    .D(_00345_),
    .Q_N(_06622_),
    .Q(\shift_storage.storage[1218] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1219]$_SDFFE_PN0P_  (.CLK(clknet_leaf_164_clk_p2c),
    .RESET_B(net1122),
    .D(_00346_),
    .Q_N(_06621_),
    .Q(\shift_storage.storage[1219] ));
 sg13g2_dfrbp_1 \shift_storage.storage[121]$_SDFFE_PN0P_  (.CLK(clknet_leaf_36_clk_p2c),
    .RESET_B(net1123),
    .D(_00347_),
    .Q_N(_06620_),
    .Q(\shift_storage.storage[121] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1220]$_SDFFE_PN0P_  (.CLK(clknet_leaf_164_clk_p2c),
    .RESET_B(net1124),
    .D(_00348_),
    .Q_N(_06619_),
    .Q(\shift_storage.storage[1220] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1221]$_SDFFE_PN0P_  (.CLK(clknet_leaf_164_clk_p2c),
    .RESET_B(net1125),
    .D(_00349_),
    .Q_N(_06618_),
    .Q(\shift_storage.storage[1221] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1222]$_SDFFE_PN0P_  (.CLK(clknet_leaf_165_clk_p2c),
    .RESET_B(net1126),
    .D(_00350_),
    .Q_N(_06617_),
    .Q(\shift_storage.storage[1222] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1223]$_SDFFE_PN0P_  (.CLK(clknet_leaf_160_clk_p2c),
    .RESET_B(net1127),
    .D(_00351_),
    .Q_N(_06616_),
    .Q(\shift_storage.storage[1223] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1224]$_SDFFE_PN0P_  (.CLK(clknet_leaf_160_clk_p2c),
    .RESET_B(net1128),
    .D(_00352_),
    .Q_N(_06615_),
    .Q(\shift_storage.storage[1224] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1225]$_SDFFE_PN0P_  (.CLK(clknet_leaf_165_clk_p2c),
    .RESET_B(net1129),
    .D(_00353_),
    .Q_N(_06614_),
    .Q(\shift_storage.storage[1225] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1226]$_SDFFE_PN0P_  (.CLK(clknet_leaf_165_clk_p2c),
    .RESET_B(net1130),
    .D(_00354_),
    .Q_N(_06613_),
    .Q(\shift_storage.storage[1226] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1227]$_SDFFE_PN0P_  (.CLK(clknet_leaf_165_clk_p2c),
    .RESET_B(net1131),
    .D(_00355_),
    .Q_N(_06612_),
    .Q(\shift_storage.storage[1227] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1228]$_SDFFE_PN0P_  (.CLK(clknet_leaf_166_clk_p2c),
    .RESET_B(net1132),
    .D(_00356_),
    .Q_N(_06611_),
    .Q(\shift_storage.storage[1228] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1229]$_SDFFE_PN0P_  (.CLK(clknet_leaf_166_clk_p2c),
    .RESET_B(net1133),
    .D(_00357_),
    .Q_N(_06610_),
    .Q(\shift_storage.storage[1229] ));
 sg13g2_dfrbp_1 \shift_storage.storage[122]$_SDFFE_PN0P_  (.CLK(clknet_leaf_244_clk_p2c),
    .RESET_B(net1134),
    .D(_00358_),
    .Q_N(_06609_),
    .Q(\shift_storage.storage[122] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1230]$_SDFFE_PN0P_  (.CLK(clknet_leaf_164_clk_p2c),
    .RESET_B(net1135),
    .D(_00359_),
    .Q_N(_06608_),
    .Q(\shift_storage.storage[1230] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1231]$_SDFFE_PN0P_  (.CLK(clknet_leaf_167_clk_p2c),
    .RESET_B(net1136),
    .D(_00360_),
    .Q_N(_06607_),
    .Q(\shift_storage.storage[1231] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1232]$_SDFFE_PN0P_  (.CLK(clknet_leaf_167_clk_p2c),
    .RESET_B(net1137),
    .D(_00361_),
    .Q_N(_06606_),
    .Q(\shift_storage.storage[1232] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1233]$_SDFFE_PN0P_  (.CLK(clknet_leaf_167_clk_p2c),
    .RESET_B(net1138),
    .D(_00362_),
    .Q_N(_06605_),
    .Q(\shift_storage.storage[1233] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1234]$_SDFFE_PN0P_  (.CLK(clknet_leaf_167_clk_p2c),
    .RESET_B(net1139),
    .D(_00363_),
    .Q_N(_06604_),
    .Q(\shift_storage.storage[1234] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1235]$_SDFFE_PN0P_  (.CLK(clknet_leaf_167_clk_p2c),
    .RESET_B(net1140),
    .D(_00364_),
    .Q_N(_06603_),
    .Q(\shift_storage.storage[1235] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1236]$_SDFFE_PN0P_  (.CLK(clknet_leaf_168_clk_p2c),
    .RESET_B(net1141),
    .D(_00365_),
    .Q_N(_06602_),
    .Q(\shift_storage.storage[1236] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1237]$_SDFFE_PN0P_  (.CLK(clknet_leaf_168_clk_p2c),
    .RESET_B(net1142),
    .D(_00366_),
    .Q_N(_06601_),
    .Q(\shift_storage.storage[1237] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1238]$_SDFFE_PN0P_  (.CLK(clknet_leaf_168_clk_p2c),
    .RESET_B(net1143),
    .D(_00367_),
    .Q_N(_06600_),
    .Q(\shift_storage.storage[1238] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1239]$_SDFFE_PN0P_  (.CLK(clknet_leaf_108_clk_p2c),
    .RESET_B(net1144),
    .D(_00368_),
    .Q_N(_06599_),
    .Q(\shift_storage.storage[1239] ));
 sg13g2_dfrbp_1 \shift_storage.storage[123]$_SDFFE_PN0P_  (.CLK(clknet_leaf_244_clk_p2c),
    .RESET_B(net1145),
    .D(_00369_),
    .Q_N(_06598_),
    .Q(\shift_storage.storage[123] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1240]$_SDFFE_PN0P_  (.CLK(clknet_leaf_108_clk_p2c),
    .RESET_B(net1146),
    .D(_00370_),
    .Q_N(_06597_),
    .Q(\shift_storage.storage[1240] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1241]$_SDFFE_PN0P_  (.CLK(clknet_leaf_109_clk_p2c),
    .RESET_B(net1147),
    .D(_00371_),
    .Q_N(_06596_),
    .Q(\shift_storage.storage[1241] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1242]$_SDFFE_PN0P_  (.CLK(clknet_leaf_109_clk_p2c),
    .RESET_B(net1148),
    .D(_00372_),
    .Q_N(_06595_),
    .Q(\shift_storage.storage[1242] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1243]$_SDFFE_PN0P_  (.CLK(clknet_leaf_109_clk_p2c),
    .RESET_B(net1149),
    .D(_00373_),
    .Q_N(_06594_),
    .Q(\shift_storage.storage[1243] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1244]$_SDFFE_PN0P_  (.CLK(clknet_leaf_111_clk_p2c),
    .RESET_B(net1150),
    .D(_00374_),
    .Q_N(_06593_),
    .Q(\shift_storage.storage[1244] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1245]$_SDFFE_PN0P_  (.CLK(clknet_leaf_112_clk_p2c),
    .RESET_B(net1151),
    .D(_00375_),
    .Q_N(_06592_),
    .Q(\shift_storage.storage[1245] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1246]$_SDFFE_PN0P_  (.CLK(clknet_leaf_112_clk_p2c),
    .RESET_B(net1152),
    .D(_00376_),
    .Q_N(_06591_),
    .Q(\shift_storage.storage[1246] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1247]$_SDFFE_PN0P_  (.CLK(clknet_leaf_103_clk_p2c),
    .RESET_B(net1153),
    .D(_00377_),
    .Q_N(_06590_),
    .Q(\shift_storage.storage[1247] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1248]$_SDFFE_PN0P_  (.CLK(clknet_leaf_103_clk_p2c),
    .RESET_B(net1154),
    .D(_00378_),
    .Q_N(_06589_),
    .Q(\shift_storage.storage[1248] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1249]$_SDFFE_PN0P_  (.CLK(clknet_leaf_103_clk_p2c),
    .RESET_B(net1155),
    .D(_00379_),
    .Q_N(_06588_),
    .Q(\shift_storage.storage[1249] ));
 sg13g2_dfrbp_1 \shift_storage.storage[124]$_SDFFE_PN0P_  (.CLK(clknet_leaf_35_clk_p2c),
    .RESET_B(net1156),
    .D(_00380_),
    .Q_N(_06587_),
    .Q(\shift_storage.storage[124] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1250]$_SDFFE_PN0P_  (.CLK(clknet_leaf_103_clk_p2c),
    .RESET_B(net1157),
    .D(_00381_),
    .Q_N(_06586_),
    .Q(\shift_storage.storage[1250] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1251]$_SDFFE_PN0P_  (.CLK(clknet_leaf_103_clk_p2c),
    .RESET_B(net1158),
    .D(_00382_),
    .Q_N(_06585_),
    .Q(\shift_storage.storage[1251] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1252]$_SDFFE_PN0P_  (.CLK(clknet_leaf_102_clk_p2c),
    .RESET_B(net1159),
    .D(_00383_),
    .Q_N(_06584_),
    .Q(\shift_storage.storage[1252] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1253]$_SDFFE_PN0P_  (.CLK(clknet_leaf_113_clk_p2c),
    .RESET_B(net1160),
    .D(_00384_),
    .Q_N(_06583_),
    .Q(\shift_storage.storage[1253] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1254]$_SDFFE_PN0P_  (.CLK(clknet_leaf_113_clk_p2c),
    .RESET_B(net1161),
    .D(_00385_),
    .Q_N(_06582_),
    .Q(\shift_storage.storage[1254] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1255]$_SDFFE_PN0P_  (.CLK(clknet_leaf_113_clk_p2c),
    .RESET_B(net1162),
    .D(_00386_),
    .Q_N(_06581_),
    .Q(\shift_storage.storage[1255] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1256]$_SDFFE_PN0P_  (.CLK(clknet_leaf_101_clk_p2c),
    .RESET_B(net1163),
    .D(_00387_),
    .Q_N(_06580_),
    .Q(\shift_storage.storage[1256] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1257]$_SDFFE_PN0P_  (.CLK(clknet_leaf_101_clk_p2c),
    .RESET_B(net1164),
    .D(_00388_),
    .Q_N(_06579_),
    .Q(\shift_storage.storage[1257] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1258]$_SDFFE_PN0P_  (.CLK(clknet_leaf_90_clk_p2c),
    .RESET_B(net1165),
    .D(_00389_),
    .Q_N(_06578_),
    .Q(\shift_storage.storage[1258] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1259]$_SDFFE_PN0P_  (.CLK(clknet_leaf_90_clk_p2c),
    .RESET_B(net1166),
    .D(_00390_),
    .Q_N(_06577_),
    .Q(\shift_storage.storage[1259] ));
 sg13g2_dfrbp_1 \shift_storage.storage[125]$_SDFFE_PN0P_  (.CLK(clknet_leaf_34_clk_p2c),
    .RESET_B(net1167),
    .D(_00391_),
    .Q_N(_06576_),
    .Q(\shift_storage.storage[125] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1260]$_SDFFE_PN0P_  (.CLK(clknet_leaf_90_clk_p2c),
    .RESET_B(net1168),
    .D(_00392_),
    .Q_N(_06575_),
    .Q(\shift_storage.storage[1260] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1261]$_SDFFE_PN0P_  (.CLK(clknet_leaf_90_clk_p2c),
    .RESET_B(net1169),
    .D(_00393_),
    .Q_N(_06574_),
    .Q(\shift_storage.storage[1261] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1262]$_SDFFE_PN0P_  (.CLK(clknet_leaf_89_clk_p2c),
    .RESET_B(net1170),
    .D(_00394_),
    .Q_N(_06573_),
    .Q(\shift_storage.storage[1262] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1263]$_SDFFE_PN0P_  (.CLK(clknet_leaf_88_clk_p2c),
    .RESET_B(net1171),
    .D(_00395_),
    .Q_N(_06572_),
    .Q(\shift_storage.storage[1263] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1264]$_SDFFE_PN0P_  (.CLK(clknet_leaf_88_clk_p2c),
    .RESET_B(net1172),
    .D(_00396_),
    .Q_N(_06571_),
    .Q(\shift_storage.storage[1264] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1265]$_SDFFE_PN0P_  (.CLK(clknet_leaf_88_clk_p2c),
    .RESET_B(net1173),
    .D(_00397_),
    .Q_N(_06570_),
    .Q(\shift_storage.storage[1265] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1266]$_SDFFE_PN0P_  (.CLK(clknet_leaf_88_clk_p2c),
    .RESET_B(net1174),
    .D(_00398_),
    .Q_N(_06569_),
    .Q(\shift_storage.storage[1266] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1267]$_SDFFE_PN0P_  (.CLK(clknet_leaf_88_clk_p2c),
    .RESET_B(net1175),
    .D(_00399_),
    .Q_N(_06568_),
    .Q(\shift_storage.storage[1267] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1268]$_SDFFE_PN0P_  (.CLK(clknet_leaf_88_clk_p2c),
    .RESET_B(net1176),
    .D(_00400_),
    .Q_N(_06567_),
    .Q(\shift_storage.storage[1268] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1269]$_SDFFE_PN0P_  (.CLK(clknet_leaf_89_clk_p2c),
    .RESET_B(net1177),
    .D(_00401_),
    .Q_N(_06566_),
    .Q(\shift_storage.storage[1269] ));
 sg13g2_dfrbp_1 \shift_storage.storage[126]$_SDFFE_PN0P_  (.CLK(clknet_leaf_35_clk_p2c),
    .RESET_B(net1178),
    .D(_00402_),
    .Q_N(_06565_),
    .Q(\shift_storage.storage[126] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1270]$_SDFFE_PN0P_  (.CLK(clknet_leaf_89_clk_p2c),
    .RESET_B(net1179),
    .D(_00403_),
    .Q_N(_06564_),
    .Q(\shift_storage.storage[1270] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1271]$_SDFFE_PN0P_  (.CLK(clknet_leaf_89_clk_p2c),
    .RESET_B(net1180),
    .D(_00404_),
    .Q_N(_06563_),
    .Q(\shift_storage.storage[1271] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1272]$_SDFFE_PN0P_  (.CLK(clknet_leaf_89_clk_p2c),
    .RESET_B(net1181),
    .D(_00405_),
    .Q_N(_06562_),
    .Q(\shift_storage.storage[1272] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1273]$_SDFFE_PN0P_  (.CLK(clknet_leaf_89_clk_p2c),
    .RESET_B(net1182),
    .D(_00406_),
    .Q_N(_06561_),
    .Q(\shift_storage.storage[1273] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1274]$_SDFFE_PN0P_  (.CLK(clknet_leaf_122_clk_p2c),
    .RESET_B(net1183),
    .D(_00407_),
    .Q_N(_06560_),
    .Q(\shift_storage.storage[1274] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1275]$_SDFFE_PN0P_  (.CLK(clknet_leaf_121_clk_p2c),
    .RESET_B(net1184),
    .D(_00408_),
    .Q_N(_06559_),
    .Q(\shift_storage.storage[1275] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1276]$_SDFFE_PN0P_  (.CLK(clknet_leaf_122_clk_p2c),
    .RESET_B(net1185),
    .D(_00409_),
    .Q_N(_06558_),
    .Q(\shift_storage.storage[1276] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1277]$_SDFFE_PN0P_  (.CLK(clknet_leaf_121_clk_p2c),
    .RESET_B(net1186),
    .D(_00410_),
    .Q_N(_06557_),
    .Q(\shift_storage.storage[1277] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1278]$_SDFFE_PN0P_  (.CLK(clknet_leaf_113_clk_p2c),
    .RESET_B(net1187),
    .D(_00411_),
    .Q_N(_06556_),
    .Q(\shift_storage.storage[1278] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1279]$_SDFFE_PN0P_  (.CLK(clknet_leaf_113_clk_p2c),
    .RESET_B(net1188),
    .D(_00412_),
    .Q_N(_06555_),
    .Q(\shift_storage.storage[1279] ));
 sg13g2_dfrbp_1 \shift_storage.storage[127]$_SDFFE_PN0P_  (.CLK(clknet_leaf_34_clk_p2c),
    .RESET_B(net1189),
    .D(_00413_),
    .Q_N(_06554_),
    .Q(\shift_storage.storage[127] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1280]$_SDFFE_PN0P_  (.CLK(clknet_leaf_114_clk_p2c),
    .RESET_B(net1190),
    .D(_00414_),
    .Q_N(_06553_),
    .Q(\shift_storage.storage[1280] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1281]$_SDFFE_PN0P_  (.CLK(clknet_leaf_113_clk_p2c),
    .RESET_B(net1191),
    .D(_00415_),
    .Q_N(_06552_),
    .Q(\shift_storage.storage[1281] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1282]$_SDFFE_PN0P_  (.CLK(clknet_leaf_121_clk_p2c),
    .RESET_B(net1192),
    .D(_00416_),
    .Q_N(_06551_),
    .Q(\shift_storage.storage[1282] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1283]$_SDFFE_PN0P_  (.CLK(clknet_leaf_121_clk_p2c),
    .RESET_B(net1193),
    .D(_00417_),
    .Q_N(_06550_),
    .Q(\shift_storage.storage[1283] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1284]$_SDFFE_PN0P_  (.CLK(clknet_leaf_121_clk_p2c),
    .RESET_B(net1194),
    .D(_00418_),
    .Q_N(_06549_),
    .Q(\shift_storage.storage[1284] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1285]$_SDFFE_PN0P_  (.CLK(clknet_leaf_121_clk_p2c),
    .RESET_B(net1195),
    .D(_00419_),
    .Q_N(_06548_),
    .Q(\shift_storage.storage[1285] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1286]$_SDFFE_PN0P_  (.CLK(clknet_leaf_120_clk_p2c),
    .RESET_B(net1196),
    .D(_00420_),
    .Q_N(_06547_),
    .Q(\shift_storage.storage[1286] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1287]$_SDFFE_PN0P_  (.CLK(clknet_leaf_122_clk_p2c),
    .RESET_B(net1197),
    .D(_00421_),
    .Q_N(_06546_),
    .Q(\shift_storage.storage[1287] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1288]$_SDFFE_PN0P_  (.CLK(clknet_leaf_122_clk_p2c),
    .RESET_B(net1198),
    .D(_00422_),
    .Q_N(_06545_),
    .Q(\shift_storage.storage[1288] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1289]$_SDFFE_PN0P_  (.CLK(clknet_leaf_123_clk_p2c),
    .RESET_B(net1199),
    .D(_00423_),
    .Q_N(_06544_),
    .Q(\shift_storage.storage[1289] ));
 sg13g2_dfrbp_1 \shift_storage.storage[128]$_SDFFE_PN0P_  (.CLK(clknet_leaf_34_clk_p2c),
    .RESET_B(net1200),
    .D(_00424_),
    .Q_N(_06543_),
    .Q(\shift_storage.storage[128] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1290]$_SDFFE_PN0P_  (.CLK(clknet_leaf_123_clk_p2c),
    .RESET_B(net1201),
    .D(_00425_),
    .Q_N(_06542_),
    .Q(\shift_storage.storage[1290] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1291]$_SDFFE_PN0P_  (.CLK(clknet_leaf_123_clk_p2c),
    .RESET_B(net1202),
    .D(_00426_),
    .Q_N(_06541_),
    .Q(\shift_storage.storage[1291] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1292]$_SDFFE_PN0P_  (.CLK(clknet_leaf_123_clk_p2c),
    .RESET_B(net1203),
    .D(_00427_),
    .Q_N(_06540_),
    .Q(\shift_storage.storage[1292] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1293]$_SDFFE_PN0P_  (.CLK(clknet_leaf_124_clk_p2c),
    .RESET_B(net1204),
    .D(_00428_),
    .Q_N(_06539_),
    .Q(\shift_storage.storage[1293] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1294]$_SDFFE_PN0P_  (.CLK(clknet_leaf_124_clk_p2c),
    .RESET_B(net1205),
    .D(_00429_),
    .Q_N(_06538_),
    .Q(\shift_storage.storage[1294] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1295]$_SDFFE_PN0P_  (.CLK(clknet_leaf_124_clk_p2c),
    .RESET_B(net1206),
    .D(_00430_),
    .Q_N(_06537_),
    .Q(\shift_storage.storage[1295] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1296]$_SDFFE_PN0P_  (.CLK(clknet_leaf_124_clk_p2c),
    .RESET_B(net1207),
    .D(_00431_),
    .Q_N(_06536_),
    .Q(\shift_storage.storage[1296] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1297]$_SDFFE_PN0P_  (.CLK(clknet_leaf_125_clk_p2c),
    .RESET_B(net1208),
    .D(_00432_),
    .Q_N(_06535_),
    .Q(\shift_storage.storage[1297] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1298]$_SDFFE_PN0P_  (.CLK(clknet_leaf_125_clk_p2c),
    .RESET_B(net1209),
    .D(_00433_),
    .Q_N(_06534_),
    .Q(\shift_storage.storage[1298] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1299]$_SDFFE_PN0P_  (.CLK(clknet_leaf_123_clk_p2c),
    .RESET_B(net1210),
    .D(_00434_),
    .Q_N(_06533_),
    .Q(\shift_storage.storage[1299] ));
 sg13g2_dfrbp_1 \shift_storage.storage[129]$_SDFFE_PN0P_  (.CLK(clknet_leaf_33_clk_p2c),
    .RESET_B(net1211),
    .D(_00435_),
    .Q_N(_06532_),
    .Q(\shift_storage.storage[129] ));
 sg13g2_dfrbp_1 \shift_storage.storage[12]$_SDFFE_PN0P_  (.CLK(clknet_leaf_70_clk_p2c),
    .RESET_B(net1212),
    .D(_00436_),
    .Q_N(_06531_),
    .Q(\shift_storage.storage[12] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1300]$_SDFFE_PN0P_  (.CLK(clknet_leaf_125_clk_p2c),
    .RESET_B(net1213),
    .D(_00437_),
    .Q_N(_06530_),
    .Q(\shift_storage.storage[1300] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1301]$_SDFFE_PN0P_  (.CLK(clknet_leaf_125_clk_p2c),
    .RESET_B(net1214),
    .D(_00438_),
    .Q_N(_06529_),
    .Q(\shift_storage.storage[1301] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1302]$_SDFFE_PN0P_  (.CLK(clknet_leaf_125_clk_p2c),
    .RESET_B(net1215),
    .D(_00439_),
    .Q_N(_06528_),
    .Q(\shift_storage.storage[1302] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1303]$_SDFFE_PN0P_  (.CLK(clknet_leaf_87_clk_p2c),
    .RESET_B(net1216),
    .D(_00440_),
    .Q_N(_06527_),
    .Q(\shift_storage.storage[1303] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1304]$_SDFFE_PN0P_  (.CLK(clknet_leaf_125_clk_p2c),
    .RESET_B(net1217),
    .D(_00441_),
    .Q_N(_06526_),
    .Q(\shift_storage.storage[1304] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1305]$_SDFFE_PN0P_  (.CLK(clknet_leaf_126_clk_p2c),
    .RESET_B(net1218),
    .D(_00442_),
    .Q_N(_06525_),
    .Q(\shift_storage.storage[1305] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1306]$_SDFFE_PN0P_  (.CLK(clknet_leaf_126_clk_p2c),
    .RESET_B(net1219),
    .D(_00443_),
    .Q_N(_06524_),
    .Q(\shift_storage.storage[1306] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1307]$_SDFFE_PN0P_  (.CLK(clknet_leaf_126_clk_p2c),
    .RESET_B(net1220),
    .D(_00444_),
    .Q_N(_06523_),
    .Q(\shift_storage.storage[1307] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1308]$_SDFFE_PN0P_  (.CLK(clknet_leaf_126_clk_p2c),
    .RESET_B(net1221),
    .D(_00445_),
    .Q_N(_06522_),
    .Q(\shift_storage.storage[1308] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1309]$_SDFFE_PN0P_  (.CLK(clknet_leaf_126_clk_p2c),
    .RESET_B(net1222),
    .D(_00446_),
    .Q_N(_06521_),
    .Q(\shift_storage.storage[1309] ));
 sg13g2_dfrbp_1 \shift_storage.storage[130]$_SDFFE_PN0P_  (.CLK(clknet_leaf_33_clk_p2c),
    .RESET_B(net1223),
    .D(_00447_),
    .Q_N(_06520_),
    .Q(\shift_storage.storage[130] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1310]$_SDFFE_PN0P_  (.CLK(clknet_leaf_127_clk_p2c),
    .RESET_B(net1224),
    .D(_00448_),
    .Q_N(_06519_),
    .Q(\shift_storage.storage[1310] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1311]$_SDFFE_PN0P_  (.CLK(clknet_leaf_127_clk_p2c),
    .RESET_B(net1225),
    .D(_00449_),
    .Q_N(_06518_),
    .Q(\shift_storage.storage[1311] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1312]$_SDFFE_PN0P_  (.CLK(clknet_leaf_127_clk_p2c),
    .RESET_B(net1226),
    .D(_00450_),
    .Q_N(_06517_),
    .Q(\shift_storage.storage[1312] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1313]$_SDFFE_PN0P_  (.CLK(clknet_leaf_127_clk_p2c),
    .RESET_B(net1227),
    .D(_00451_),
    .Q_N(_06516_),
    .Q(\shift_storage.storage[1313] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1314]$_SDFFE_PN0P_  (.CLK(clknet_leaf_127_clk_p2c),
    .RESET_B(net1228),
    .D(_00452_),
    .Q_N(_06515_),
    .Q(\shift_storage.storage[1314] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1315]$_SDFFE_PN0P_  (.CLK(clknet_leaf_130_clk_p2c),
    .RESET_B(net1229),
    .D(_00453_),
    .Q_N(_06514_),
    .Q(\shift_storage.storage[1315] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1316]$_SDFFE_PN0P_  (.CLK(clknet_leaf_130_clk_p2c),
    .RESET_B(net1230),
    .D(_00454_),
    .Q_N(_06513_),
    .Q(\shift_storage.storage[1316] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1317]$_SDFFE_PN0P_  (.CLK(clknet_leaf_131_clk_p2c),
    .RESET_B(net1231),
    .D(_00455_),
    .Q_N(_06512_),
    .Q(\shift_storage.storage[1317] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1318]$_SDFFE_PN0P_  (.CLK(clknet_leaf_131_clk_p2c),
    .RESET_B(net1232),
    .D(_00456_),
    .Q_N(_06511_),
    .Q(\shift_storage.storage[1318] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1319]$_SDFFE_PN0P_  (.CLK(clknet_leaf_131_clk_p2c),
    .RESET_B(net1233),
    .D(_00457_),
    .Q_N(_06510_),
    .Q(\shift_storage.storage[1319] ));
 sg13g2_dfrbp_1 \shift_storage.storage[131]$_SDFFE_PN0P_  (.CLK(clknet_leaf_32_clk_p2c),
    .RESET_B(net1234),
    .D(_00458_),
    .Q_N(_06509_),
    .Q(\shift_storage.storage[131] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1320]$_SDFFE_PN0P_  (.CLK(clknet_leaf_132_clk_p2c),
    .RESET_B(net1235),
    .D(_00459_),
    .Q_N(_06508_),
    .Q(\shift_storage.storage[1320] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1321]$_SDFFE_PN0P_  (.CLK(clknet_leaf_135_clk_p2c),
    .RESET_B(net1236),
    .D(_00460_),
    .Q_N(_06507_),
    .Q(\shift_storage.storage[1321] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1322]$_SDFFE_PN0P_  (.CLK(clknet_leaf_135_clk_p2c),
    .RESET_B(net1237),
    .D(_00461_),
    .Q_N(_06506_),
    .Q(\shift_storage.storage[1322] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1323]$_SDFFE_PN0P_  (.CLK(clknet_leaf_135_clk_p2c),
    .RESET_B(net1238),
    .D(_00462_),
    .Q_N(_06505_),
    .Q(\shift_storage.storage[1323] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1324]$_SDFFE_PN0P_  (.CLK(clknet_leaf_136_clk_p2c),
    .RESET_B(net1239),
    .D(_00463_),
    .Q_N(_06504_),
    .Q(\shift_storage.storage[1324] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1325]$_SDFFE_PN0P_  (.CLK(clknet_leaf_136_clk_p2c),
    .RESET_B(net1240),
    .D(_00464_),
    .Q_N(_06503_),
    .Q(\shift_storage.storage[1325] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1326]$_SDFFE_PN0P_  (.CLK(clknet_leaf_136_clk_p2c),
    .RESET_B(net1241),
    .D(_00465_),
    .Q_N(_06502_),
    .Q(\shift_storage.storage[1326] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1327]$_SDFFE_PN0P_  (.CLK(clknet_leaf_138_clk_p2c),
    .RESET_B(net1242),
    .D(_00466_),
    .Q_N(_06501_),
    .Q(\shift_storage.storage[1327] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1328]$_SDFFE_PN0P_  (.CLK(clknet_leaf_137_clk_p2c),
    .RESET_B(net1243),
    .D(_00467_),
    .Q_N(_06500_),
    .Q(\shift_storage.storage[1328] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1329]$_SDFFE_PN0P_  (.CLK(clknet_leaf_138_clk_p2c),
    .RESET_B(net1244),
    .D(_00468_),
    .Q_N(_06499_),
    .Q(\shift_storage.storage[1329] ));
 sg13g2_dfrbp_1 \shift_storage.storage[132]$_SDFFE_PN0P_  (.CLK(clknet_leaf_32_clk_p2c),
    .RESET_B(net1245),
    .D(_00469_),
    .Q_N(_06498_),
    .Q(\shift_storage.storage[132] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1330]$_SDFFE_PN0P_  (.CLK(clknet_leaf_138_clk_p2c),
    .RESET_B(net1246),
    .D(_00470_),
    .Q_N(_06497_),
    .Q(\shift_storage.storage[1330] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1331]$_SDFFE_PN0P_  (.CLK(clknet_leaf_138_clk_p2c),
    .RESET_B(net1247),
    .D(_00471_),
    .Q_N(_06496_),
    .Q(\shift_storage.storage[1331] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1332]$_SDFFE_PN0P_  (.CLK(clknet_leaf_139_clk_p2c),
    .RESET_B(net1248),
    .D(_00472_),
    .Q_N(_06495_),
    .Q(\shift_storage.storage[1332] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1333]$_SDFFE_PN0P_  (.CLK(clknet_leaf_138_clk_p2c),
    .RESET_B(net1249),
    .D(_00473_),
    .Q_N(_06494_),
    .Q(\shift_storage.storage[1333] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1334]$_SDFFE_PN0P_  (.CLK(clknet_leaf_139_clk_p2c),
    .RESET_B(net1250),
    .D(_00474_),
    .Q_N(_06493_),
    .Q(\shift_storage.storage[1334] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1335]$_SDFFE_PN0P_  (.CLK(clknet_leaf_139_clk_p2c),
    .RESET_B(net1251),
    .D(_00475_),
    .Q_N(_06492_),
    .Q(\shift_storage.storage[1335] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1336]$_SDFFE_PN0P_  (.CLK(clknet_leaf_139_clk_p2c),
    .RESET_B(net1252),
    .D(_00476_),
    .Q_N(_06491_),
    .Q(\shift_storage.storage[1336] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1337]$_SDFFE_PN0P_  (.CLK(clknet_leaf_139_clk_p2c),
    .RESET_B(net1253),
    .D(_00477_),
    .Q_N(_06490_),
    .Q(\shift_storage.storage[1337] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1338]$_SDFFE_PN0P_  (.CLK(clknet_leaf_140_clk_p2c),
    .RESET_B(net1254),
    .D(_00478_),
    .Q_N(_06489_),
    .Q(\shift_storage.storage[1338] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1339]$_SDFFE_PN0P_  (.CLK(clknet_leaf_137_clk_p2c),
    .RESET_B(net1255),
    .D(_00479_),
    .Q_N(_06488_),
    .Q(\shift_storage.storage[1339] ));
 sg13g2_dfrbp_1 \shift_storage.storage[133]$_SDFFE_PN0P_  (.CLK(clknet_leaf_34_clk_p2c),
    .RESET_B(net1256),
    .D(_00480_),
    .Q_N(_06487_),
    .Q(\shift_storage.storage[133] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1340]$_SDFFE_PN0P_  (.CLK(clknet_leaf_138_clk_p2c),
    .RESET_B(net1257),
    .D(_00481_),
    .Q_N(_06486_),
    .Q(\shift_storage.storage[1340] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1341]$_SDFFE_PN0P_  (.CLK(clknet_leaf_137_clk_p2c),
    .RESET_B(net1258),
    .D(_00482_),
    .Q_N(_06485_),
    .Q(\shift_storage.storage[1341] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1342]$_SDFFE_PN0P_  (.CLK(clknet_leaf_137_clk_p2c),
    .RESET_B(net1259),
    .D(_00483_),
    .Q_N(_06484_),
    .Q(\shift_storage.storage[1342] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1343]$_SDFFE_PN0P_  (.CLK(clknet_leaf_137_clk_p2c),
    .RESET_B(net1260),
    .D(_00484_),
    .Q_N(_06483_),
    .Q(\shift_storage.storage[1343] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1344]$_SDFFE_PN0P_  (.CLK(clknet_leaf_136_clk_p2c),
    .RESET_B(net1261),
    .D(_00485_),
    .Q_N(_06482_),
    .Q(\shift_storage.storage[1344] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1345]$_SDFFE_PN0P_  (.CLK(clknet_leaf_136_clk_p2c),
    .RESET_B(net1262),
    .D(_00486_),
    .Q_N(_06481_),
    .Q(\shift_storage.storage[1345] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1346]$_SDFFE_PN0P_  (.CLK(clknet_leaf_135_clk_p2c),
    .RESET_B(net1263),
    .D(_00487_),
    .Q_N(_06480_),
    .Q(\shift_storage.storage[1346] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1347]$_SDFFE_PN0P_  (.CLK(clknet_leaf_131_clk_p2c),
    .RESET_B(net1264),
    .D(_00488_),
    .Q_N(_06479_),
    .Q(\shift_storage.storage[1347] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1348]$_SDFFE_PN0P_  (.CLK(clknet_leaf_130_clk_p2c),
    .RESET_B(net1265),
    .D(_00489_),
    .Q_N(_06478_),
    .Q(\shift_storage.storage[1348] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1349]$_SDFFE_PN0P_  (.CLK(clknet_leaf_129_clk_p2c),
    .RESET_B(net1266),
    .D(_00490_),
    .Q_N(_06477_),
    .Q(\shift_storage.storage[1349] ));
 sg13g2_dfrbp_1 \shift_storage.storage[134]$_SDFFE_PN0P_  (.CLK(clknet_leaf_32_clk_p2c),
    .RESET_B(net1267),
    .D(_00491_),
    .Q_N(_06476_),
    .Q(\shift_storage.storage[134] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1350]$_SDFFE_PN0P_  (.CLK(clknet_leaf_130_clk_p2c),
    .RESET_B(net1268),
    .D(_00492_),
    .Q_N(_06475_),
    .Q(\shift_storage.storage[1350] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1351]$_SDFFE_PN0P_  (.CLK(clknet_leaf_129_clk_p2c),
    .RESET_B(net1269),
    .D(_00493_),
    .Q_N(_06474_),
    .Q(\shift_storage.storage[1351] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1352]$_SDFFE_PN0P_  (.CLK(clknet_leaf_127_clk_p2c),
    .RESET_B(net1270),
    .D(_00494_),
    .Q_N(_06473_),
    .Q(\shift_storage.storage[1352] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1353]$_SDFFE_PN0P_  (.CLK(clknet_leaf_126_clk_p2c),
    .RESET_B(net1271),
    .D(_00495_),
    .Q_N(_06472_),
    .Q(\shift_storage.storage[1353] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1354]$_SDFFE_PN0P_  (.CLK(clknet_leaf_128_clk_p2c),
    .RESET_B(net1272),
    .D(_00496_),
    .Q_N(_06471_),
    .Q(\shift_storage.storage[1354] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1355]$_SDFFE_PN0P_  (.CLK(clknet_leaf_128_clk_p2c),
    .RESET_B(net1273),
    .D(_00497_),
    .Q_N(_06470_),
    .Q(\shift_storage.storage[1355] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1356]$_SDFFE_PN0P_  (.CLK(clknet_leaf_128_clk_p2c),
    .RESET_B(net1274),
    .D(_00498_),
    .Q_N(_06469_),
    .Q(\shift_storage.storage[1356] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1357]$_SDFFE_PN0P_  (.CLK(clknet_leaf_128_clk_p2c),
    .RESET_B(net1275),
    .D(_00499_),
    .Q_N(_06468_),
    .Q(\shift_storage.storage[1357] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1358]$_SDFFE_PN0P_  (.CLK(clknet_leaf_124_clk_p2c),
    .RESET_B(net1276),
    .D(_00500_),
    .Q_N(_06467_),
    .Q(\shift_storage.storage[1358] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1359]$_SDFFE_PN0P_  (.CLK(clknet_leaf_124_clk_p2c),
    .RESET_B(net1277),
    .D(_00501_),
    .Q_N(_06466_),
    .Q(\shift_storage.storage[1359] ));
 sg13g2_dfrbp_1 \shift_storage.storage[135]$_SDFFE_PN0P_  (.CLK(clknet_leaf_31_clk_p2c),
    .RESET_B(net1278),
    .D(_00502_),
    .Q_N(_06465_),
    .Q(\shift_storage.storage[135] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1360]$_SDFFE_PN0P_  (.CLK(clknet_leaf_123_clk_p2c),
    .RESET_B(net1279),
    .D(_00503_),
    .Q_N(_06464_),
    .Q(\shift_storage.storage[1360] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1361]$_SDFFE_PN0P_  (.CLK(clknet_leaf_119_clk_p2c),
    .RESET_B(net1280),
    .D(_00504_),
    .Q_N(_06463_),
    .Q(\shift_storage.storage[1361] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1362]$_SDFFE_PN0P_  (.CLK(clknet_leaf_119_clk_p2c),
    .RESET_B(net1281),
    .D(_00505_),
    .Q_N(_06462_),
    .Q(\shift_storage.storage[1362] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1363]$_SDFFE_PN0P_  (.CLK(clknet_leaf_119_clk_p2c),
    .RESET_B(net1282),
    .D(_00506_),
    .Q_N(_06461_),
    .Q(\shift_storage.storage[1363] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1364]$_SDFFE_PN0P_  (.CLK(clknet_leaf_120_clk_p2c),
    .RESET_B(net1283),
    .D(_00507_),
    .Q_N(_06460_),
    .Q(\shift_storage.storage[1364] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1365]$_SDFFE_PN0P_  (.CLK(clknet_leaf_120_clk_p2c),
    .RESET_B(net1284),
    .D(_00508_),
    .Q_N(_06459_),
    .Q(\shift_storage.storage[1365] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1366]$_SDFFE_PN0P_  (.CLK(clknet_leaf_120_clk_p2c),
    .RESET_B(net1285),
    .D(_00509_),
    .Q_N(_06458_),
    .Q(\shift_storage.storage[1366] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1367]$_SDFFE_PN0P_  (.CLK(clknet_leaf_120_clk_p2c),
    .RESET_B(net1286),
    .D(_00510_),
    .Q_N(_06457_),
    .Q(\shift_storage.storage[1367] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1368]$_SDFFE_PN0P_  (.CLK(clknet_leaf_120_clk_p2c),
    .RESET_B(net1287),
    .D(_00511_),
    .Q_N(_06456_),
    .Q(\shift_storage.storage[1368] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1369]$_SDFFE_PN0P_  (.CLK(clknet_leaf_114_clk_p2c),
    .RESET_B(net1288),
    .D(_00512_),
    .Q_N(_06455_),
    .Q(\shift_storage.storage[1369] ));
 sg13g2_dfrbp_1 \shift_storage.storage[136]$_SDFFE_PN0P_  (.CLK(clknet_leaf_31_clk_p2c),
    .RESET_B(net1289),
    .D(_00513_),
    .Q_N(_06454_),
    .Q(\shift_storage.storage[136] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1370]$_SDFFE_PN0P_  (.CLK(clknet_leaf_114_clk_p2c),
    .RESET_B(net1290),
    .D(_00514_),
    .Q_N(_06453_),
    .Q(\shift_storage.storage[1370] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1371]$_SDFFE_PN0P_  (.CLK(clknet_leaf_114_clk_p2c),
    .RESET_B(net1291),
    .D(_00515_),
    .Q_N(_06452_),
    .Q(\shift_storage.storage[1371] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1372]$_SDFFE_PN0P_  (.CLK(clknet_leaf_114_clk_p2c),
    .RESET_B(net1292),
    .D(_00516_),
    .Q_N(_06451_),
    .Q(\shift_storage.storage[1372] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1373]$_SDFFE_PN0P_  (.CLK(clknet_leaf_114_clk_p2c),
    .RESET_B(net1293),
    .D(_00517_),
    .Q_N(_06450_),
    .Q(\shift_storage.storage[1373] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1374]$_SDFFE_PN0P_  (.CLK(clknet_leaf_115_clk_p2c),
    .RESET_B(net1294),
    .D(_00518_),
    .Q_N(_06449_),
    .Q(\shift_storage.storage[1374] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1375]$_SDFFE_PN0P_  (.CLK(clknet_leaf_115_clk_p2c),
    .RESET_B(net1295),
    .D(_00519_),
    .Q_N(_06448_),
    .Q(\shift_storage.storage[1375] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1376]$_SDFFE_PN0P_  (.CLK(clknet_leaf_115_clk_p2c),
    .RESET_B(net1296),
    .D(_00520_),
    .Q_N(_06447_),
    .Q(\shift_storage.storage[1376] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1377]$_SDFFE_PN0P_  (.CLK(clknet_leaf_116_clk_p2c),
    .RESET_B(net1297),
    .D(_00521_),
    .Q_N(_06446_),
    .Q(\shift_storage.storage[1377] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1378]$_SDFFE_PN0P_  (.CLK(clknet_leaf_116_clk_p2c),
    .RESET_B(net1298),
    .D(_00522_),
    .Q_N(_06445_),
    .Q(\shift_storage.storage[1378] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1379]$_SDFFE_PN0P_  (.CLK(clknet_leaf_159_clk_p2c),
    .RESET_B(net1299),
    .D(_00523_),
    .Q_N(_06444_),
    .Q(\shift_storage.storage[1379] ));
 sg13g2_dfrbp_1 \shift_storage.storage[137]$_SDFFE_PN0P_  (.CLK(clknet_leaf_32_clk_p2c),
    .RESET_B(net1300),
    .D(_00524_),
    .Q_N(_06443_),
    .Q(\shift_storage.storage[137] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1380]$_SDFFE_PN0P_  (.CLK(clknet_leaf_159_clk_p2c),
    .RESET_B(net1301),
    .D(_00525_),
    .Q_N(_06442_),
    .Q(\shift_storage.storage[1380] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1381]$_SDFFE_PN0P_  (.CLK(clknet_leaf_158_clk_p2c),
    .RESET_B(net1302),
    .D(_00526_),
    .Q_N(_06441_),
    .Q(\shift_storage.storage[1381] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1382]$_SDFFE_PN0P_  (.CLK(clknet_leaf_158_clk_p2c),
    .RESET_B(net1303),
    .D(_00527_),
    .Q_N(_06440_),
    .Q(\shift_storage.storage[1382] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1383]$_SDFFE_PN0P_  (.CLK(clknet_leaf_161_clk_p2c),
    .RESET_B(net1304),
    .D(_00528_),
    .Q_N(_06439_),
    .Q(\shift_storage.storage[1383] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1384]$_SDFFE_PN0P_  (.CLK(clknet_leaf_161_clk_p2c),
    .RESET_B(net1305),
    .D(_00529_),
    .Q_N(_06438_),
    .Q(\shift_storage.storage[1384] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1385]$_SDFFE_PN0P_  (.CLK(clknet_leaf_160_clk_p2c),
    .RESET_B(net1306),
    .D(_00530_),
    .Q_N(_06437_),
    .Q(\shift_storage.storage[1385] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1386]$_SDFFE_PN0P_  (.CLK(clknet_leaf_160_clk_p2c),
    .RESET_B(net1307),
    .D(_00531_),
    .Q_N(_06436_),
    .Q(\shift_storage.storage[1386] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1387]$_SDFFE_PN0P_  (.CLK(clknet_leaf_160_clk_p2c),
    .RESET_B(net1308),
    .D(_00532_),
    .Q_N(_06435_),
    .Q(\shift_storage.storage[1387] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1388]$_SDFFE_PN0P_  (.CLK(clknet_leaf_165_clk_p2c),
    .RESET_B(net1309),
    .D(_00533_),
    .Q_N(_06434_),
    .Q(\shift_storage.storage[1388] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1389]$_SDFFE_PN0P_  (.CLK(clknet_leaf_166_clk_p2c),
    .RESET_B(net1310),
    .D(_00534_),
    .Q_N(_06433_),
    .Q(\shift_storage.storage[1389] ));
 sg13g2_dfrbp_1 \shift_storage.storage[138]$_SDFFE_PN0P_  (.CLK(clknet_leaf_29_clk_p2c),
    .RESET_B(net1311),
    .D(_00535_),
    .Q_N(_06432_),
    .Q(\shift_storage.storage[138] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1390]$_SDFFE_PN0P_  (.CLK(clknet_leaf_110_clk_p2c),
    .RESET_B(net1312),
    .D(_00536_),
    .Q_N(_06431_),
    .Q(\shift_storage.storage[1390] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1391]$_SDFFE_PN0P_  (.CLK(clknet_leaf_110_clk_p2c),
    .RESET_B(net1313),
    .D(_00537_),
    .Q_N(_06430_),
    .Q(\shift_storage.storage[1391] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1392]$_SDFFE_PN0P_  (.CLK(clknet_leaf_116_clk_p2c),
    .RESET_B(net1314),
    .D(_00538_),
    .Q_N(_06429_),
    .Q(\shift_storage.storage[1392] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1393]$_SDFFE_PN0P_  (.CLK(clknet_leaf_111_clk_p2c),
    .RESET_B(net1315),
    .D(_00539_),
    .Q_N(_06428_),
    .Q(\shift_storage.storage[1393] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1394]$_SDFFE_PN0P_  (.CLK(clknet_leaf_115_clk_p2c),
    .RESET_B(net1316),
    .D(_00540_),
    .Q_N(_06427_),
    .Q(\shift_storage.storage[1394] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1395]$_SDFFE_PN0P_  (.CLK(clknet_leaf_111_clk_p2c),
    .RESET_B(net1317),
    .D(_00541_),
    .Q_N(_06426_),
    .Q(\shift_storage.storage[1395] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1396]$_SDFFE_PN0P_  (.CLK(clknet_leaf_115_clk_p2c),
    .RESET_B(net1318),
    .D(_00542_),
    .Q_N(_06425_),
    .Q(\shift_storage.storage[1396] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1397]$_SDFFE_PN0P_  (.CLK(clknet_leaf_115_clk_p2c),
    .RESET_B(net1319),
    .D(_00543_),
    .Q_N(_06424_),
    .Q(\shift_storage.storage[1397] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1398]$_SDFFE_PN0P_  (.CLK(clknet_leaf_114_clk_p2c),
    .RESET_B(net1320),
    .D(_00544_),
    .Q_N(_06423_),
    .Q(\shift_storage.storage[1398] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1399]$_SDFFE_PN0P_  (.CLK(clknet_leaf_112_clk_p2c),
    .RESET_B(net1321),
    .D(_00545_),
    .Q_N(_06422_),
    .Q(\shift_storage.storage[1399] ));
 sg13g2_dfrbp_1 \shift_storage.storage[139]$_SDFFE_PN0P_  (.CLK(clknet_leaf_28_clk_p2c),
    .RESET_B(net1322),
    .D(_00546_),
    .Q_N(_06421_),
    .Q(\shift_storage.storage[139] ));
 sg13g2_dfrbp_1 \shift_storage.storage[13]$_SDFFE_PN0P_  (.CLK(clknet_leaf_70_clk_p2c),
    .RESET_B(net1323),
    .D(_00547_),
    .Q_N(_06420_),
    .Q(\shift_storage.storage[13] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1400]$_SDFFE_PN0P_  (.CLK(clknet_leaf_112_clk_p2c),
    .RESET_B(net1324),
    .D(_00548_),
    .Q_N(_06419_),
    .Q(\shift_storage.storage[1400] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1401]$_SDFFE_PN0P_  (.CLK(clknet_leaf_112_clk_p2c),
    .RESET_B(net1325),
    .D(_00549_),
    .Q_N(_06418_),
    .Q(\shift_storage.storage[1401] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1402]$_SDFFE_PN0P_  (.CLK(clknet_leaf_112_clk_p2c),
    .RESET_B(net1326),
    .D(_00550_),
    .Q_N(_06417_),
    .Q(\shift_storage.storage[1402] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1403]$_SDFFE_PN0P_  (.CLK(clknet_leaf_111_clk_p2c),
    .RESET_B(net1327),
    .D(_00551_),
    .Q_N(_06416_),
    .Q(\shift_storage.storage[1403] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1404]$_SDFFE_PN0P_  (.CLK(clknet_leaf_111_clk_p2c),
    .RESET_B(net1328),
    .D(_00552_),
    .Q_N(_06415_),
    .Q(\shift_storage.storage[1404] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1405]$_SDFFE_PN0P_  (.CLK(clknet_leaf_111_clk_p2c),
    .RESET_B(net1329),
    .D(_00553_),
    .Q_N(_06414_),
    .Q(\shift_storage.storage[1405] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1406]$_SDFFE_PN0P_  (.CLK(clknet_leaf_110_clk_p2c),
    .RESET_B(net1330),
    .D(_00554_),
    .Q_N(_06413_),
    .Q(\shift_storage.storage[1406] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1407]$_SDFFE_PN0P_  (.CLK(clknet_leaf_110_clk_p2c),
    .RESET_B(net1331),
    .D(_00555_),
    .Q_N(_06412_),
    .Q(\shift_storage.storage[1407] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1408]$_SDFFE_PN0P_  (.CLK(clknet_leaf_110_clk_p2c),
    .RESET_B(net1332),
    .D(_00556_),
    .Q_N(_06411_),
    .Q(\shift_storage.storage[1408] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1409]$_SDFFE_PN0P_  (.CLK(clknet_leaf_110_clk_p2c),
    .RESET_B(net1333),
    .D(_00557_),
    .Q_N(_06410_),
    .Q(\shift_storage.storage[1409] ));
 sg13g2_dfrbp_1 \shift_storage.storage[140]$_SDFFE_PN0P_  (.CLK(clknet_leaf_29_clk_p2c),
    .RESET_B(net1334),
    .D(_00558_),
    .Q_N(_06409_),
    .Q(\shift_storage.storage[140] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1410]$_SDFFE_PN0P_  (.CLK(clknet_leaf_166_clk_p2c),
    .RESET_B(net1335),
    .D(_00559_),
    .Q_N(_06408_),
    .Q(\shift_storage.storage[1410] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1411]$_SDFFE_PN0P_  (.CLK(clknet_leaf_166_clk_p2c),
    .RESET_B(net1336),
    .D(_00560_),
    .Q_N(_06407_),
    .Q(\shift_storage.storage[1411] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1412]$_SDFFE_PN0P_  (.CLK(clknet_leaf_166_clk_p2c),
    .RESET_B(net1337),
    .D(_00561_),
    .Q_N(_06406_),
    .Q(\shift_storage.storage[1412] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1413]$_SDFFE_PN0P_  (.CLK(clknet_leaf_168_clk_p2c),
    .RESET_B(net1338),
    .D(_00562_),
    .Q_N(_06405_),
    .Q(\shift_storage.storage[1413] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1414]$_SDFFE_PN0P_  (.CLK(clknet_leaf_108_clk_p2c),
    .RESET_B(net1339),
    .D(_00563_),
    .Q_N(_06404_),
    .Q(\shift_storage.storage[1414] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1415]$_SDFFE_PN0P_  (.CLK(clknet_leaf_108_clk_p2c),
    .RESET_B(net1340),
    .D(_00564_),
    .Q_N(_06403_),
    .Q(\shift_storage.storage[1415] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1416]$_SDFFE_PN0P_  (.CLK(clknet_leaf_108_clk_p2c),
    .RESET_B(net1341),
    .D(_00565_),
    .Q_N(_06402_),
    .Q(\shift_storage.storage[1416] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1417]$_SDFFE_PN0P_  (.CLK(clknet_leaf_108_clk_p2c),
    .RESET_B(net1342),
    .D(_00566_),
    .Q_N(_06401_),
    .Q(\shift_storage.storage[1417] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1418]$_SDFFE_PN0P_  (.CLK(clknet_leaf_107_clk_p2c),
    .RESET_B(net1343),
    .D(_00567_),
    .Q_N(_06400_),
    .Q(\shift_storage.storage[1418] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1419]$_SDFFE_PN0P_  (.CLK(clknet_leaf_107_clk_p2c),
    .RESET_B(net1344),
    .D(_00568_),
    .Q_N(_06399_),
    .Q(\shift_storage.storage[1419] ));
 sg13g2_dfrbp_1 \shift_storage.storage[141]$_SDFFE_PN0P_  (.CLK(clknet_leaf_30_clk_p2c),
    .RESET_B(net1345),
    .D(_00569_),
    .Q_N(_06398_),
    .Q(\shift_storage.storage[141] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1420]$_SDFFE_PN0P_  (.CLK(clknet_leaf_107_clk_p2c),
    .RESET_B(net1346),
    .D(_00570_),
    .Q_N(_06397_),
    .Q(\shift_storage.storage[1420] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1421]$_SDFFE_PN0P_  (.CLK(clknet_leaf_107_clk_p2c),
    .RESET_B(net1347),
    .D(_00571_),
    .Q_N(_06396_),
    .Q(\shift_storage.storage[1421] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1422]$_SDFFE_PN0P_  (.CLK(clknet_leaf_109_clk_p2c),
    .RESET_B(net1348),
    .D(_00572_),
    .Q_N(_06395_),
    .Q(\shift_storage.storage[1422] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1423]$_SDFFE_PN0P_  (.CLK(clknet_leaf_109_clk_p2c),
    .RESET_B(net1349),
    .D(_00573_),
    .Q_N(_06394_),
    .Q(\shift_storage.storage[1423] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1424]$_SDFFE_PN0P_  (.CLK(clknet_leaf_109_clk_p2c),
    .RESET_B(net1350),
    .D(_00574_),
    .Q_N(_06393_),
    .Q(\shift_storage.storage[1424] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1425]$_SDFFE_PN0P_  (.CLK(clknet_leaf_109_clk_p2c),
    .RESET_B(net1351),
    .D(_00575_),
    .Q_N(_06392_),
    .Q(\shift_storage.storage[1425] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1426]$_SDFFE_PN0P_  (.CLK(clknet_leaf_106_clk_p2c),
    .RESET_B(net1352),
    .D(_00576_),
    .Q_N(_06391_),
    .Q(\shift_storage.storage[1426] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1427]$_SDFFE_PN0P_  (.CLK(clknet_leaf_106_clk_p2c),
    .RESET_B(net1353),
    .D(_00577_),
    .Q_N(_06390_),
    .Q(\shift_storage.storage[1427] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1428]$_SDFFE_PN0P_  (.CLK(clknet_leaf_103_clk_p2c),
    .RESET_B(net1354),
    .D(_00578_),
    .Q_N(_06389_),
    .Q(\shift_storage.storage[1428] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1429]$_SDFFE_PN0P_  (.CLK(clknet_leaf_104_clk_p2c),
    .RESET_B(net1355),
    .D(_00579_),
    .Q_N(_06388_),
    .Q(\shift_storage.storage[1429] ));
 sg13g2_dfrbp_1 \shift_storage.storage[142]$_SDFFE_PN0P_  (.CLK(clknet_leaf_30_clk_p2c),
    .RESET_B(net1356),
    .D(_00580_),
    .Q_N(_06387_),
    .Q(\shift_storage.storage[142] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1430]$_SDFFE_PN0P_  (.CLK(clknet_leaf_104_clk_p2c),
    .RESET_B(net1357),
    .D(_00581_),
    .Q_N(_06386_),
    .Q(\shift_storage.storage[1430] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1431]$_SDFFE_PN0P_  (.CLK(clknet_leaf_104_clk_p2c),
    .RESET_B(net1358),
    .D(_00582_),
    .Q_N(_06385_),
    .Q(\shift_storage.storage[1431] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1432]$_SDFFE_PN0P_  (.CLK(clknet_leaf_104_clk_p2c),
    .RESET_B(net1359),
    .D(_00583_),
    .Q_N(_06384_),
    .Q(\shift_storage.storage[1432] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1433]$_SDFFE_PN0P_  (.CLK(clknet_leaf_104_clk_p2c),
    .RESET_B(net1360),
    .D(_00584_),
    .Q_N(_06383_),
    .Q(\shift_storage.storage[1433] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1434]$_SDFFE_PN0P_  (.CLK(clknet_leaf_102_clk_p2c),
    .RESET_B(net1361),
    .D(_00585_),
    .Q_N(_06382_),
    .Q(\shift_storage.storage[1434] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1435]$_SDFFE_PN0P_  (.CLK(clknet_leaf_102_clk_p2c),
    .RESET_B(net1362),
    .D(_00586_),
    .Q_N(_06381_),
    .Q(\shift_storage.storage[1435] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1436]$_SDFFE_PN0P_  (.CLK(clknet_leaf_102_clk_p2c),
    .RESET_B(net1363),
    .D(_00587_),
    .Q_N(_06380_),
    .Q(\shift_storage.storage[1436] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1437]$_SDFFE_PN0P_  (.CLK(clknet_leaf_102_clk_p2c),
    .RESET_B(net1364),
    .D(_00588_),
    .Q_N(_06379_),
    .Q(\shift_storage.storage[1437] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1438]$_SDFFE_PN0P_  (.CLK(clknet_leaf_102_clk_p2c),
    .RESET_B(net1365),
    .D(_00589_),
    .Q_N(_06378_),
    .Q(\shift_storage.storage[1438] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1439]$_SDFFE_PN0P_  (.CLK(clknet_leaf_100_clk_p2c),
    .RESET_B(net1366),
    .D(_00590_),
    .Q_N(_06377_),
    .Q(\shift_storage.storage[1439] ));
 sg13g2_dfrbp_1 \shift_storage.storage[143]$_SDFFE_PN0P_  (.CLK(clknet_leaf_30_clk_p2c),
    .RESET_B(net1367),
    .D(_00591_),
    .Q_N(_06376_),
    .Q(\shift_storage.storage[143] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1440]$_SDFFE_PN0P_  (.CLK(clknet_leaf_101_clk_p2c),
    .RESET_B(net1368),
    .D(_00592_),
    .Q_N(_06375_),
    .Q(\shift_storage.storage[1440] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1441]$_SDFFE_PN0P_  (.CLK(clknet_leaf_101_clk_p2c),
    .RESET_B(net1369),
    .D(_00593_),
    .Q_N(_06374_),
    .Q(\shift_storage.storage[1441] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1442]$_SDFFE_PN0P_  (.CLK(clknet_leaf_101_clk_p2c),
    .RESET_B(net1370),
    .D(_00594_),
    .Q_N(_06373_),
    .Q(\shift_storage.storage[1442] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1443]$_SDFFE_PN0P_  (.CLK(clknet_leaf_90_clk_p2c),
    .RESET_B(net1371),
    .D(_00595_),
    .Q_N(_06372_),
    .Q(\shift_storage.storage[1443] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1444]$_SDFFE_PN0P_  (.CLK(clknet_leaf_91_clk_p2c),
    .RESET_B(net1372),
    .D(_00596_),
    .Q_N(_06371_),
    .Q(\shift_storage.storage[1444] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1445]$_SDFFE_PN0P_  (.CLK(clknet_leaf_90_clk_p2c),
    .RESET_B(net1373),
    .D(_00597_),
    .Q_N(_06370_),
    .Q(\shift_storage.storage[1445] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1446]$_SDFFE_PN0P_  (.CLK(clknet_leaf_91_clk_p2c),
    .RESET_B(net1374),
    .D(_00598_),
    .Q_N(_06369_),
    .Q(\shift_storage.storage[1446] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1447]$_SDFFE_PN0P_  (.CLK(clknet_leaf_92_clk_p2c),
    .RESET_B(net1375),
    .D(_00599_),
    .Q_N(_06368_),
    .Q(\shift_storage.storage[1447] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1448]$_SDFFE_PN0P_  (.CLK(clknet_leaf_92_clk_p2c),
    .RESET_B(net1376),
    .D(_00600_),
    .Q_N(_06367_),
    .Q(\shift_storage.storage[1448] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1449]$_SDFFE_PN0P_  (.CLK(clknet_leaf_92_clk_p2c),
    .RESET_B(net1377),
    .D(_00601_),
    .Q_N(_06366_),
    .Q(\shift_storage.storage[1449] ));
 sg13g2_dfrbp_1 \shift_storage.storage[144]$_SDFFE_PN0P_  (.CLK(clknet_leaf_30_clk_p2c),
    .RESET_B(net1378),
    .D(_00602_),
    .Q_N(_06365_),
    .Q(\shift_storage.storage[144] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1450]$_SDFFE_PN0P_  (.CLK(clknet_leaf_92_clk_p2c),
    .RESET_B(net1379),
    .D(_00603_),
    .Q_N(_06364_),
    .Q(\shift_storage.storage[1450] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1451]$_SDFFE_PN0P_  (.CLK(clknet_leaf_87_clk_p2c),
    .RESET_B(net1380),
    .D(_00604_),
    .Q_N(_06363_),
    .Q(\shift_storage.storage[1451] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1452]$_SDFFE_PN0P_  (.CLK(clknet_leaf_87_clk_p2c),
    .RESET_B(net1381),
    .D(_00605_),
    .Q_N(_06362_),
    .Q(\shift_storage.storage[1452] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1453]$_SDFFE_PN0P_  (.CLK(clknet_leaf_87_clk_p2c),
    .RESET_B(net1382),
    .D(_00606_),
    .Q_N(_06361_),
    .Q(\shift_storage.storage[1453] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1454]$_SDFFE_PN0P_  (.CLK(clknet_leaf_87_clk_p2c),
    .RESET_B(net1383),
    .D(_00607_),
    .Q_N(_06360_),
    .Q(\shift_storage.storage[1454] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1455]$_SDFFE_PN0P_  (.CLK(clknet_leaf_87_clk_p2c),
    .RESET_B(net1384),
    .D(_00608_),
    .Q_N(_06359_),
    .Q(\shift_storage.storage[1455] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1456]$_SDFFE_PN0P_  (.CLK(clknet_leaf_86_clk_p2c),
    .RESET_B(net1385),
    .D(_00609_),
    .Q_N(_06358_),
    .Q(\shift_storage.storage[1456] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1457]$_SDFFE_PN0P_  (.CLK(clknet_leaf_86_clk_p2c),
    .RESET_B(net1386),
    .D(_00610_),
    .Q_N(_06357_),
    .Q(\shift_storage.storage[1457] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1458]$_SDFFE_PN0P_  (.CLK(clknet_leaf_93_clk_p2c),
    .RESET_B(net1387),
    .D(_00611_),
    .Q_N(_06356_),
    .Q(\shift_storage.storage[1458] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1459]$_SDFFE_PN0P_  (.CLK(clknet_leaf_92_clk_p2c),
    .RESET_B(net1388),
    .D(_00612_),
    .Q_N(_06355_),
    .Q(\shift_storage.storage[1459] ));
 sg13g2_dfrbp_1 \shift_storage.storage[145]$_SDFFE_PN0P_  (.CLK(clknet_leaf_31_clk_p2c),
    .RESET_B(net1389),
    .D(_00613_),
    .Q_N(_06354_),
    .Q(\shift_storage.storage[145] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1460]$_SDFFE_PN0P_  (.CLK(clknet_leaf_84_clk_p2c),
    .RESET_B(net1390),
    .D(_00614_),
    .Q_N(_06353_),
    .Q(\shift_storage.storage[1460] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1461]$_SDFFE_PN0P_  (.CLK(clknet_leaf_93_clk_p2c),
    .RESET_B(net1391),
    .D(_00615_),
    .Q_N(_06352_),
    .Q(\shift_storage.storage[1461] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1462]$_SDFFE_PN0P_  (.CLK(clknet_leaf_93_clk_p2c),
    .RESET_B(net1392),
    .D(_00616_),
    .Q_N(_06351_),
    .Q(\shift_storage.storage[1462] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1463]$_SDFFE_PN0P_  (.CLK(clknet_leaf_93_clk_p2c),
    .RESET_B(net1393),
    .D(_00617_),
    .Q_N(_06350_),
    .Q(\shift_storage.storage[1463] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1464]$_SDFFE_PN0P_  (.CLK(clknet_leaf_84_clk_p2c),
    .RESET_B(net1394),
    .D(_00618_),
    .Q_N(_06349_),
    .Q(\shift_storage.storage[1464] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1465]$_SDFFE_PN0P_  (.CLK(clknet_leaf_84_clk_p2c),
    .RESET_B(net1395),
    .D(_00619_),
    .Q_N(_06348_),
    .Q(\shift_storage.storage[1465] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1466]$_SDFFE_PN0P_  (.CLK(clknet_leaf_84_clk_p2c),
    .RESET_B(net1396),
    .D(_00620_),
    .Q_N(_06347_),
    .Q(\shift_storage.storage[1466] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1467]$_SDFFE_PN0P_  (.CLK(clknet_leaf_84_clk_p2c),
    .RESET_B(net1397),
    .D(_00621_),
    .Q_N(_06346_),
    .Q(\shift_storage.storage[1467] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1468]$_SDFFE_PN0P_  (.CLK(clknet_leaf_85_clk_p2c),
    .RESET_B(net1398),
    .D(_00622_),
    .Q_N(_06345_),
    .Q(\shift_storage.storage[1468] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1469]$_SDFFE_PN0P_  (.CLK(clknet_leaf_85_clk_p2c),
    .RESET_B(net1399),
    .D(_00623_),
    .Q_N(_06344_),
    .Q(\shift_storage.storage[1469] ));
 sg13g2_dfrbp_1 \shift_storage.storage[146]$_SDFFE_PN0P_  (.CLK(clknet_leaf_30_clk_p2c),
    .RESET_B(net1400),
    .D(_00624_),
    .Q_N(_06343_),
    .Q(\shift_storage.storage[146] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1470]$_SDFFE_PN0P_  (.CLK(clknet_leaf_85_clk_p2c),
    .RESET_B(net1401),
    .D(_00625_),
    .Q_N(_06342_),
    .Q(\shift_storage.storage[1470] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1471]$_SDFFE_PN0P_  (.CLK(clknet_leaf_85_clk_p2c),
    .RESET_B(net1402),
    .D(_00626_),
    .Q_N(_06341_),
    .Q(\shift_storage.storage[1471] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1472]$_SDFFE_PN0P_  (.CLK(clknet_leaf_86_clk_p2c),
    .RESET_B(net1403),
    .D(_00627_),
    .Q_N(_06340_),
    .Q(\shift_storage.storage[1472] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1473]$_SDFFE_PN0P_  (.CLK(clknet_leaf_86_clk_p2c),
    .RESET_B(net1404),
    .D(_00628_),
    .Q_N(_06339_),
    .Q(\shift_storage.storage[1473] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1474]$_SDFFE_PN0P_  (.CLK(clknet_leaf_85_clk_p2c),
    .RESET_B(net1405),
    .D(_00629_),
    .Q_N(_06338_),
    .Q(\shift_storage.storage[1474] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1475]$_SDFFE_PN0P_  (.CLK(clknet_leaf_85_clk_p2c),
    .RESET_B(net1406),
    .D(_00630_),
    .Q_N(_06337_),
    .Q(\shift_storage.storage[1475] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1476]$_SDFFE_PN0P_  (.CLK(clknet_leaf_83_clk_p2c),
    .RESET_B(net1407),
    .D(_00631_),
    .Q_N(_06336_),
    .Q(\shift_storage.storage[1476] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1477]$_SDFFE_PN0P_  (.CLK(clknet_leaf_83_clk_p2c),
    .RESET_B(net1408),
    .D(_00632_),
    .Q_N(_06335_),
    .Q(\shift_storage.storage[1477] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1478]$_SDFFE_PN0P_  (.CLK(clknet_leaf_83_clk_p2c),
    .RESET_B(net1409),
    .D(_00633_),
    .Q_N(_06334_),
    .Q(\shift_storage.storage[1478] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1479]$_SDFFE_PN0P_  (.CLK(clknet_leaf_83_clk_p2c),
    .RESET_B(net1410),
    .D(_00634_),
    .Q_N(_06333_),
    .Q(\shift_storage.storage[1479] ));
 sg13g2_dfrbp_1 \shift_storage.storage[147]$_SDFFE_PN0P_  (.CLK(clknet_leaf_31_clk_p2c),
    .RESET_B(net1411),
    .D(_00635_),
    .Q_N(_06332_),
    .Q(\shift_storage.storage[147] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1480]$_SDFFE_PN0P_  (.CLK(clknet_leaf_83_clk_p2c),
    .RESET_B(net1412),
    .D(_00636_),
    .Q_N(_06331_),
    .Q(\shift_storage.storage[1480] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1481]$_SDFFE_PN0P_  (.CLK(clknet_leaf_83_clk_p2c),
    .RESET_B(net1413),
    .D(_00637_),
    .Q_N(_06330_),
    .Q(\shift_storage.storage[1481] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1482]$_SDFFE_PN0P_  (.CLK(clknet_leaf_95_clk_p2c),
    .RESET_B(net1414),
    .D(_00638_),
    .Q_N(_06329_),
    .Q(\shift_storage.storage[1482] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1483]$_SDFFE_PN0P_  (.CLK(clknet_leaf_95_clk_p2c),
    .RESET_B(net1415),
    .D(_00639_),
    .Q_N(_06328_),
    .Q(\shift_storage.storage[1483] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1484]$_SDFFE_PN0P_  (.CLK(clknet_leaf_94_clk_p2c),
    .RESET_B(net1416),
    .D(_00640_),
    .Q_N(_06327_),
    .Q(\shift_storage.storage[1484] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1485]$_SDFFE_PN0P_  (.CLK(clknet_leaf_94_clk_p2c),
    .RESET_B(net1417),
    .D(_00641_),
    .Q_N(_06326_),
    .Q(\shift_storage.storage[1485] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1486]$_SDFFE_PN0P_  (.CLK(clknet_leaf_93_clk_p2c),
    .RESET_B(net1418),
    .D(_00642_),
    .Q_N(_06325_),
    .Q(\shift_storage.storage[1486] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1487]$_SDFFE_PN0P_  (.CLK(clknet_leaf_94_clk_p2c),
    .RESET_B(net1419),
    .D(_00643_),
    .Q_N(_06324_),
    .Q(\shift_storage.storage[1487] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1488]$_SDFFE_PN0P_  (.CLK(clknet_leaf_93_clk_p2c),
    .RESET_B(net1420),
    .D(_00644_),
    .Q_N(_06323_),
    .Q(\shift_storage.storage[1488] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1489]$_SDFFE_PN0P_  (.CLK(clknet_leaf_92_clk_p2c),
    .RESET_B(net1421),
    .D(_00645_),
    .Q_N(_06322_),
    .Q(\shift_storage.storage[1489] ));
 sg13g2_dfrbp_1 \shift_storage.storage[148]$_SDFFE_PN0P_  (.CLK(clknet_leaf_42_clk_p2c),
    .RESET_B(net1422),
    .D(_00646_),
    .Q_N(_06321_),
    .Q(\shift_storage.storage[148] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1490]$_SDFFE_PN0P_  (.CLK(clknet_leaf_91_clk_p2c),
    .RESET_B(net1423),
    .D(_00647_),
    .Q_N(_06320_),
    .Q(\shift_storage.storage[1490] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1491]$_SDFFE_PN0P_  (.CLK(clknet_leaf_91_clk_p2c),
    .RESET_B(net1424),
    .D(_00648_),
    .Q_N(_06319_),
    .Q(\shift_storage.storage[1491] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1492]$_SDFFE_PN0P_  (.CLK(clknet_leaf_91_clk_p2c),
    .RESET_B(net1425),
    .D(_00649_),
    .Q_N(_06318_),
    .Q(\shift_storage.storage[1492] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1493]$_SDFFE_PN0P_  (.CLK(clknet_leaf_91_clk_p2c),
    .RESET_B(net1426),
    .D(_00650_),
    .Q_N(_06317_),
    .Q(\shift_storage.storage[1493] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1494]$_SDFFE_PN0P_  (.CLK(clknet_leaf_100_clk_p2c),
    .RESET_B(net1427),
    .D(_00651_),
    .Q_N(_06316_),
    .Q(\shift_storage.storage[1494] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1495]$_SDFFE_PN0P_  (.CLK(clknet_leaf_100_clk_p2c),
    .RESET_B(net1428),
    .D(_00652_),
    .Q_N(_06315_),
    .Q(\shift_storage.storage[1495] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1496]$_SDFFE_PN0P_  (.CLK(clknet_leaf_100_clk_p2c),
    .RESET_B(net1429),
    .D(_00653_),
    .Q_N(_06314_),
    .Q(\shift_storage.storage[1496] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1497]$_SDFFE_PN0P_  (.CLK(clknet_leaf_99_clk_p2c),
    .RESET_B(net1430),
    .D(_00654_),
    .Q_N(_06313_),
    .Q(\shift_storage.storage[1497] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1498]$_SDFFE_PN0P_  (.CLK(clknet_leaf_99_clk_p2c),
    .RESET_B(net1431),
    .D(_00655_),
    .Q_N(_06312_),
    .Q(\shift_storage.storage[1498] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1499]$_SDFFE_PN0P_  (.CLK(clknet_leaf_99_clk_p2c),
    .RESET_B(net1432),
    .D(_00656_),
    .Q_N(_06311_),
    .Q(\shift_storage.storage[1499] ));
 sg13g2_dfrbp_1 \shift_storage.storage[149]$_SDFFE_PN0P_  (.CLK(clknet_leaf_42_clk_p2c),
    .RESET_B(net1433),
    .D(_00657_),
    .Q_N(_06310_),
    .Q(\shift_storage.storage[149] ));
 sg13g2_dfrbp_1 \shift_storage.storage[14]$_SDFFE_PN0P_  (.CLK(clknet_leaf_70_clk_p2c),
    .RESET_B(net1434),
    .D(_00658_),
    .Q_N(_06309_),
    .Q(\shift_storage.storage[14] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1500]$_SDFFE_PN0P_  (.CLK(clknet_leaf_99_clk_p2c),
    .RESET_B(net1435),
    .D(_00659_),
    .Q_N(_06308_),
    .Q(\shift_storage.storage[1500] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1501]$_SDFFE_PN0P_  (.CLK(clknet_leaf_98_clk_p2c),
    .RESET_B(net1436),
    .D(_00660_),
    .Q_N(_06307_),
    .Q(\shift_storage.storage[1501] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1502]$_SDFFE_PN0P_  (.CLK(clknet_leaf_105_clk_p2c),
    .RESET_B(net1437),
    .D(_00661_),
    .Q_N(_06306_),
    .Q(\shift_storage.storage[1502] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1503]$_SDFFE_PN0P_  (.CLK(clknet_leaf_105_clk_p2c),
    .RESET_B(net1438),
    .D(_00662_),
    .Q_N(_06305_),
    .Q(\shift_storage.storage[1503] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1504]$_SDFFE_PN0P_  (.CLK(clknet_leaf_105_clk_p2c),
    .RESET_B(net1439),
    .D(_00663_),
    .Q_N(_06304_),
    .Q(\shift_storage.storage[1504] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1505]$_SDFFE_PN0P_  (.CLK(clknet_leaf_104_clk_p2c),
    .RESET_B(net1440),
    .D(_00664_),
    .Q_N(_06303_),
    .Q(\shift_storage.storage[1505] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1506]$_SDFFE_PN0P_  (.CLK(clknet_leaf_105_clk_p2c),
    .RESET_B(net1441),
    .D(_00665_),
    .Q_N(_06302_),
    .Q(\shift_storage.storage[1506] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1507]$_SDFFE_PN0P_  (.CLK(clknet_leaf_106_clk_p2c),
    .RESET_B(net1442),
    .D(_00666_),
    .Q_N(_06301_),
    .Q(\shift_storage.storage[1507] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1508]$_SDFFE_PN0P_  (.CLK(clknet_leaf_106_clk_p2c),
    .RESET_B(net1443),
    .D(_00667_),
    .Q_N(_06300_),
    .Q(\shift_storage.storage[1508] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1509]$_SDFFE_PN0P_  (.CLK(clknet_leaf_106_clk_p2c),
    .RESET_B(net1444),
    .D(_00668_),
    .Q_N(_06299_),
    .Q(\shift_storage.storage[1509] ));
 sg13g2_dfrbp_1 \shift_storage.storage[150]$_SDFFE_PN0P_  (.CLK(clknet_leaf_42_clk_p2c),
    .RESET_B(net1445),
    .D(_00669_),
    .Q_N(_06298_),
    .Q(\shift_storage.storage[150] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1510]$_SDFFE_PN0P_  (.CLK(clknet_leaf_107_clk_p2c),
    .RESET_B(net1446),
    .D(_00670_),
    .Q_N(_06297_),
    .Q(\shift_storage.storage[1510] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1511]$_SDFFE_PN0P_  (.CLK(clknet_leaf_107_clk_p2c),
    .RESET_B(net1447),
    .D(_00671_),
    .Q_N(_06296_),
    .Q(\shift_storage.storage[1511] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1512]$_SDFFE_PN0P_  (.CLK(clknet_leaf_107_clk_p2c),
    .RESET_B(net1448),
    .D(_00672_),
    .Q_N(_06295_),
    .Q(\shift_storage.storage[1512] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1513]$_SDFFE_PN0P_  (.CLK(clknet_leaf_38_clk_p2c),
    .RESET_B(net1449),
    .D(_00673_),
    .Q_N(_06294_),
    .Q(\shift_storage.storage[1513] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1514]$_SDFFE_PN0P_  (.CLK(clknet_leaf_37_clk_p2c),
    .RESET_B(net1450),
    .D(_00674_),
    .Q_N(_06293_),
    .Q(\shift_storage.storage[1514] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1515]$_SDFFE_PN0P_  (.CLK(clknet_leaf_37_clk_p2c),
    .RESET_B(net1451),
    .D(_00675_),
    .Q_N(_06292_),
    .Q(\shift_storage.storage[1515] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1516]$_SDFFE_PN0P_  (.CLK(clknet_leaf_37_clk_p2c),
    .RESET_B(net1452),
    .D(_00676_),
    .Q_N(_06291_),
    .Q(\shift_storage.storage[1516] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1517]$_SDFFE_PN0P_  (.CLK(clknet_leaf_37_clk_p2c),
    .RESET_B(net1453),
    .D(_00677_),
    .Q_N(_06290_),
    .Q(\shift_storage.storage[1517] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1518]$_SDFFE_PN0P_  (.CLK(clknet_leaf_36_clk_p2c),
    .RESET_B(net1454),
    .D(_00678_),
    .Q_N(_06289_),
    .Q(\shift_storage.storage[1518] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1519]$_SDFFE_PN0P_  (.CLK(clknet_leaf_36_clk_p2c),
    .RESET_B(net1455),
    .D(_00679_),
    .Q_N(_06288_),
    .Q(\shift_storage.storage[1519] ));
 sg13g2_dfrbp_1 \shift_storage.storage[151]$_SDFFE_PN0P_  (.CLK(clknet_leaf_41_clk_p2c),
    .RESET_B(net1456),
    .D(_00680_),
    .Q_N(_06287_),
    .Q(\shift_storage.storage[151] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1520]$_SDFFE_PN0P_  (.CLK(clknet_leaf_36_clk_p2c),
    .RESET_B(net1457),
    .D(_00681_),
    .Q_N(_06286_),
    .Q(\shift_storage.storage[1520] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1521]$_SDFFE_PN0P_  (.CLK(clknet_leaf_36_clk_p2c),
    .RESET_B(net1458),
    .D(_00682_),
    .Q_N(_06285_),
    .Q(\shift_storage.storage[1521] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1522]$_SDFFE_PN0P_  (.CLK(clknet_leaf_243_clk_p2c),
    .RESET_B(net1459),
    .D(_00683_),
    .Q_N(_06284_),
    .Q(\shift_storage.storage[1522] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1523]$_SDFFE_PN0P_  (.CLK(clknet_leaf_243_clk_p2c),
    .RESET_B(net1460),
    .D(_00684_),
    .Q_N(_06283_),
    .Q(\shift_storage.storage[1523] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1524]$_SDFFE_PN0P_  (.CLK(clknet_leaf_168_clk_p2c),
    .RESET_B(net1461),
    .D(_00685_),
    .Q_N(_06282_),
    .Q(\shift_storage.storage[1524] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1525]$_SDFFE_PN0P_  (.CLK(clknet_leaf_168_clk_p2c),
    .RESET_B(net1462),
    .D(_00686_),
    .Q_N(_06281_),
    .Q(\shift_storage.storage[1525] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1526]$_SDFFE_PN0P_  (.CLK(clknet_leaf_169_clk_p2c),
    .RESET_B(net1463),
    .D(_00687_),
    .Q_N(_06280_),
    .Q(\shift_storage.storage[1526] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1527]$_SDFFE_PN0P_  (.CLK(clknet_leaf_169_clk_p2c),
    .RESET_B(net1464),
    .D(_00688_),
    .Q_N(_06279_),
    .Q(\shift_storage.storage[1527] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1528]$_SDFFE_PN0P_  (.CLK(clknet_leaf_169_clk_p2c),
    .RESET_B(net1465),
    .D(_00689_),
    .Q_N(_06278_),
    .Q(\shift_storage.storage[1528] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1529]$_SDFFE_PN0P_  (.CLK(clknet_leaf_242_clk_p2c),
    .RESET_B(net1466),
    .D(_00690_),
    .Q_N(_06277_),
    .Q(\shift_storage.storage[1529] ));
 sg13g2_dfrbp_1 \shift_storage.storage[152]$_SDFFE_PN0P_  (.CLK(clknet_leaf_42_clk_p2c),
    .RESET_B(net1467),
    .D(_00691_),
    .Q_N(_06276_),
    .Q(\shift_storage.storage[152] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1530]$_SDFFE_PN0P_  (.CLK(clknet_leaf_243_clk_p2c),
    .RESET_B(net1468),
    .D(_00692_),
    .Q_N(_06275_),
    .Q(\shift_storage.storage[1530] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1531]$_SDFFE_PN0P_  (.CLK(clknet_leaf_243_clk_p2c),
    .RESET_B(net1469),
    .D(_00693_),
    .Q_N(_06274_),
    .Q(\shift_storage.storage[1531] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1532]$_SDFFE_PN0P_  (.CLK(clknet_leaf_243_clk_p2c),
    .RESET_B(net1470),
    .D(_00694_),
    .Q_N(_06273_),
    .Q(\shift_storage.storage[1532] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1533]$_SDFFE_PN0P_  (.CLK(clknet_leaf_243_clk_p2c),
    .RESET_B(net1471),
    .D(_00695_),
    .Q_N(_06272_),
    .Q(\shift_storage.storage[1533] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1534]$_SDFFE_PN0P_  (.CLK(clknet_leaf_244_clk_p2c),
    .RESET_B(net1472),
    .D(_00696_),
    .Q_N(_06271_),
    .Q(\shift_storage.storage[1534] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1535]$_SDFFE_PN0P_  (.CLK(clknet_leaf_244_clk_p2c),
    .RESET_B(net1473),
    .D(_00697_),
    .Q_N(_06270_),
    .Q(\shift_storage.storage[1535] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1536]$_SDFFE_PN0P_  (.CLK(clknet_leaf_244_clk_p2c),
    .RESET_B(net1474),
    .D(_00698_),
    .Q_N(_06269_),
    .Q(\shift_storage.storage[1536] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1537]$_SDFFE_PN0P_  (.CLK(clknet_leaf_248_clk_p2c),
    .RESET_B(net1475),
    .D(_00699_),
    .Q_N(_06268_),
    .Q(\shift_storage.storage[1537] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1538]$_SDFFE_PN0P_  (.CLK(clknet_leaf_245_clk_p2c),
    .RESET_B(net1476),
    .D(_00700_),
    .Q_N(_06267_),
    .Q(\shift_storage.storage[1538] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1539]$_SDFFE_PN0P_  (.CLK(clknet_leaf_242_clk_p2c),
    .RESET_B(net1477),
    .D(_00701_),
    .Q_N(_06266_),
    .Q(\shift_storage.storage[1539] ));
 sg13g2_dfrbp_1 \shift_storage.storage[153]$_SDFFE_PN0P_  (.CLK(clknet_leaf_42_clk_p2c),
    .RESET_B(net1478),
    .D(_00702_),
    .Q_N(_06265_),
    .Q(\shift_storage.storage[153] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1540]$_SDFFE_PN0P_  (.CLK(clknet_leaf_242_clk_p2c),
    .RESET_B(net1479),
    .D(_00703_),
    .Q_N(_06264_),
    .Q(\shift_storage.storage[1540] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1541]$_SDFFE_PN0P_  (.CLK(clknet_leaf_242_clk_p2c),
    .RESET_B(net1480),
    .D(_00704_),
    .Q_N(_06263_),
    .Q(\shift_storage.storage[1541] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1542]$_SDFFE_PN0P_  (.CLK(clknet_leaf_242_clk_p2c),
    .RESET_B(net1481),
    .D(_00705_),
    .Q_N(_06262_),
    .Q(\shift_storage.storage[1542] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1543]$_SDFFE_PN0P_  (.CLK(clknet_leaf_242_clk_p2c),
    .RESET_B(net1482),
    .D(_00706_),
    .Q_N(_06261_),
    .Q(\shift_storage.storage[1543] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1544]$_SDFFE_PN0P_  (.CLK(clknet_leaf_241_clk_p2c),
    .RESET_B(net1483),
    .D(_00707_),
    .Q_N(_06260_),
    .Q(\shift_storage.storage[1544] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1545]$_SDFFE_PN0P_  (.CLK(clknet_leaf_170_clk_p2c),
    .RESET_B(net1484),
    .D(_00708_),
    .Q_N(_06259_),
    .Q(\shift_storage.storage[1545] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1546]$_SDFFE_PN0P_  (.CLK(clknet_leaf_241_clk_p2c),
    .RESET_B(net1485),
    .D(_00709_),
    .Q_N(_06258_),
    .Q(\shift_storage.storage[1546] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1547]$_SDFFE_PN0P_  (.CLK(clknet_leaf_170_clk_p2c),
    .RESET_B(net1486),
    .D(_00710_),
    .Q_N(_06257_),
    .Q(\shift_storage.storage[1547] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1548]$_SDFFE_PN0P_  (.CLK(clknet_leaf_171_clk_p2c),
    .RESET_B(net1487),
    .D(_00711_),
    .Q_N(_06256_),
    .Q(\shift_storage.storage[1548] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1549]$_SDFFE_PN0P_  (.CLK(clknet_leaf_171_clk_p2c),
    .RESET_B(net1488),
    .D(_00712_),
    .Q_N(_06255_),
    .Q(\shift_storage.storage[1549] ));
 sg13g2_dfrbp_1 \shift_storage.storage[154]$_SDFFE_PN0P_  (.CLK(clknet_leaf_43_clk_p2c),
    .RESET_B(net1489),
    .D(_00713_),
    .Q_N(_06254_),
    .Q(\shift_storage.storage[154] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1550]$_SDFFE_PN0P_  (.CLK(clknet_leaf_172_clk_p2c),
    .RESET_B(net1490),
    .D(_00714_),
    .Q_N(_06253_),
    .Q(\shift_storage.storage[1550] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1551]$_SDFFE_PN0P_  (.CLK(clknet_leaf_171_clk_p2c),
    .RESET_B(net1491),
    .D(_00715_),
    .Q_N(_06252_),
    .Q(\shift_storage.storage[1551] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1552]$_SDFFE_PN0P_  (.CLK(clknet_leaf_172_clk_p2c),
    .RESET_B(net1492),
    .D(_00716_),
    .Q_N(_06251_),
    .Q(\shift_storage.storage[1552] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1553]$_SDFFE_PN0P_  (.CLK(clknet_leaf_172_clk_p2c),
    .RESET_B(net1493),
    .D(_00717_),
    .Q_N(_06250_),
    .Q(\shift_storage.storage[1553] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1554]$_SDFFE_PN0P_  (.CLK(clknet_leaf_172_clk_p2c),
    .RESET_B(net1494),
    .D(_00718_),
    .Q_N(_06249_),
    .Q(\shift_storage.storage[1554] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1555]$_SDFFE_PN0P_  (.CLK(clknet_leaf_172_clk_p2c),
    .RESET_B(net1495),
    .D(_00719_),
    .Q_N(_06248_),
    .Q(\shift_storage.storage[1555] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1556]$_SDFFE_PN0P_  (.CLK(clknet_leaf_163_clk_p2c),
    .RESET_B(net1496),
    .D(_00720_),
    .Q_N(_06247_),
    .Q(\shift_storage.storage[1556] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1557]$_SDFFE_PN0P_  (.CLK(clknet_leaf_163_clk_p2c),
    .RESET_B(net1497),
    .D(_00721_),
    .Q_N(_06246_),
    .Q(\shift_storage.storage[1557] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1558]$_SDFFE_PN0P_  (.CLK(clknet_leaf_163_clk_p2c),
    .RESET_B(net1498),
    .D(_00722_),
    .Q_N(_06245_),
    .Q(\shift_storage.storage[1558] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1559]$_SDFFE_PN0P_  (.CLK(clknet_leaf_163_clk_p2c),
    .RESET_B(net1499),
    .D(_00723_),
    .Q_N(_06244_),
    .Q(\shift_storage.storage[1559] ));
 sg13g2_dfrbp_1 \shift_storage.storage[155]$_SDFFE_PN0P_  (.CLK(clknet_leaf_52_clk_p2c),
    .RESET_B(net1500),
    .D(_00724_),
    .Q_N(_06243_),
    .Q(\shift_storage.storage[155] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1560]$_SDFFE_PN0P_  (.CLK(clknet_leaf_162_clk_p2c),
    .RESET_B(net1501),
    .D(_00725_),
    .Q_N(_06242_),
    .Q(\shift_storage.storage[1560] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1561]$_SDFFE_PN0P_  (.CLK(clknet_leaf_162_clk_p2c),
    .RESET_B(net1502),
    .D(_00726_),
    .Q_N(_06241_),
    .Q(\shift_storage.storage[1561] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1562]$_SDFFE_PN0P_  (.CLK(clknet_leaf_161_clk_p2c),
    .RESET_B(net1503),
    .D(_00727_),
    .Q_N(_06240_),
    .Q(\shift_storage.storage[1562] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1563]$_SDFFE_PN0P_  (.CLK(clknet_leaf_161_clk_p2c),
    .RESET_B(net1504),
    .D(_00728_),
    .Q_N(_06239_),
    .Q(\shift_storage.storage[1563] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1564]$_SDFFE_PN0P_  (.CLK(clknet_leaf_161_clk_p2c),
    .RESET_B(net1505),
    .D(_00729_),
    .Q_N(_06238_),
    .Q(\shift_storage.storage[1564] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1565]$_SDFFE_PN0P_  (.CLK(clknet_leaf_161_clk_p2c),
    .RESET_B(net1506),
    .D(_00730_),
    .Q_N(_06237_),
    .Q(\shift_storage.storage[1565] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1566]$_SDFFE_PN0P_  (.CLK(clknet_leaf_153_clk_p2c),
    .RESET_B(net1507),
    .D(_00731_),
    .Q_N(_06236_),
    .Q(\shift_storage.storage[1566] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1567]$_SDFFE_PN0P_  (.CLK(clknet_leaf_158_clk_p2c),
    .RESET_B(net1508),
    .D(_00732_),
    .Q_N(_06235_),
    .Q(\shift_storage.storage[1567] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1568]$_SDFFE_PN0P_  (.CLK(clknet_leaf_158_clk_p2c),
    .RESET_B(net1509),
    .D(_00733_),
    .Q_N(_06234_),
    .Q(\shift_storage.storage[1568] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1569]$_SDFFE_PN0P_  (.CLK(clknet_leaf_153_clk_p2c),
    .RESET_B(net1510),
    .D(_00734_),
    .Q_N(_06233_),
    .Q(\shift_storage.storage[1569] ));
 sg13g2_dfrbp_1 \shift_storage.storage[156]$_SDFFE_PN0P_  (.CLK(clknet_leaf_52_clk_p2c),
    .RESET_B(net1511),
    .D(_00735_),
    .Q_N(_06232_),
    .Q(\shift_storage.storage[156] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1570]$_SDFFE_PN0P_  (.CLK(clknet_leaf_156_clk_p2c),
    .RESET_B(net1512),
    .D(_00736_),
    .Q_N(_06231_),
    .Q(\shift_storage.storage[1570] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1571]$_SDFFE_PN0P_  (.CLK(clknet_leaf_153_clk_p2c),
    .RESET_B(net1513),
    .D(_00737_),
    .Q_N(_06230_),
    .Q(\shift_storage.storage[1571] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1572]$_SDFFE_PN0P_  (.CLK(clknet_leaf_153_clk_p2c),
    .RESET_B(net1514),
    .D(_00738_),
    .Q_N(_06229_),
    .Q(\shift_storage.storage[1572] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1573]$_SDFFE_PN0P_  (.CLK(clknet_leaf_155_clk_p2c),
    .RESET_B(net1515),
    .D(_00739_),
    .Q_N(_06228_),
    .Q(\shift_storage.storage[1573] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1574]$_SDFFE_PN0P_  (.CLK(clknet_leaf_154_clk_p2c),
    .RESET_B(net1516),
    .D(_00740_),
    .Q_N(_06227_),
    .Q(\shift_storage.storage[1574] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1575]$_SDFFE_PN0P_  (.CLK(clknet_leaf_154_clk_p2c),
    .RESET_B(net1517),
    .D(_00741_),
    .Q_N(_06226_),
    .Q(\shift_storage.storage[1575] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1576]$_SDFFE_PN0P_  (.CLK(clknet_leaf_154_clk_p2c),
    .RESET_B(net1518),
    .D(_00742_),
    .Q_N(_06225_),
    .Q(\shift_storage.storage[1576] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1577]$_SDFFE_PN0P_  (.CLK(clknet_leaf_154_clk_p2c),
    .RESET_B(net1519),
    .D(_00743_),
    .Q_N(_06224_),
    .Q(\shift_storage.storage[1577] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1578]$_SDFFE_PN0P_  (.CLK(clknet_leaf_147_clk_p2c),
    .RESET_B(net1520),
    .D(_00744_),
    .Q_N(_06223_),
    .Q(\shift_storage.storage[1578] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1579]$_SDFFE_PN0P_  (.CLK(clknet_leaf_147_clk_p2c),
    .RESET_B(net1521),
    .D(_00745_),
    .Q_N(_06222_),
    .Q(\shift_storage.storage[1579] ));
 sg13g2_dfrbp_1 \shift_storage.storage[157]$_SDFFE_PN0P_  (.CLK(clknet_leaf_44_clk_p2c),
    .RESET_B(net1522),
    .D(_00746_),
    .Q_N(_06221_),
    .Q(\shift_storage.storage[157] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1580]$_SDFFE_PN0P_  (.CLK(clknet_leaf_146_clk_p2c),
    .RESET_B(net1523),
    .D(_00747_),
    .Q_N(_06220_),
    .Q(\shift_storage.storage[1580] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1581]$_SDFFE_PN0P_  (.CLK(clknet_leaf_145_clk_p2c),
    .RESET_B(net1524),
    .D(_00748_),
    .Q_N(_06219_),
    .Q(\shift_storage.storage[1581] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1582]$_SDFFE_PN0P_  (.CLK(clknet_leaf_145_clk_p2c),
    .RESET_B(net1525),
    .D(_00749_),
    .Q_N(_06218_),
    .Q(\shift_storage.storage[1582] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1583]$_SDFFE_PN0P_  (.CLK(clknet_leaf_145_clk_p2c),
    .RESET_B(net1526),
    .D(_00750_),
    .Q_N(_06217_),
    .Q(\shift_storage.storage[1583] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1584]$_SDFFE_PN0P_  (.CLK(clknet_leaf_146_clk_p2c),
    .RESET_B(net1527),
    .D(_00751_),
    .Q_N(_06216_),
    .Q(\shift_storage.storage[1584] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1585]$_SDFFE_PN0P_  (.CLK(clknet_leaf_146_clk_p2c),
    .RESET_B(net1528),
    .D(_00752_),
    .Q_N(_06215_),
    .Q(\shift_storage.storage[1585] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1586]$_SDFFE_PN0P_  (.CLK(clknet_leaf_146_clk_p2c),
    .RESET_B(net1529),
    .D(_00753_),
    .Q_N(_06214_),
    .Q(\shift_storage.storage[1586] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1587]$_SDFFE_PN0P_  (.CLK(clknet_leaf_142_clk_p2c),
    .RESET_B(net1530),
    .D(_00754_),
    .Q_N(_06213_),
    .Q(\shift_storage.storage[1587] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1588]$_SDFFE_PN0P_  (.CLK(clknet_leaf_142_clk_p2c),
    .RESET_B(net1531),
    .D(_00755_),
    .Q_N(_06212_),
    .Q(\shift_storage.storage[1588] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1589]$_SDFFE_PN0P_  (.CLK(clknet_leaf_142_clk_p2c),
    .RESET_B(net1532),
    .D(_00756_),
    .Q_N(_06211_),
    .Q(\shift_storage.storage[1589] ));
 sg13g2_dfrbp_1 \shift_storage.storage[158]$_SDFFE_PN0P_  (.CLK(clknet_leaf_47_clk_p2c),
    .RESET_B(net1533),
    .D(_00757_),
    .Q_N(_06210_),
    .Q(\shift_storage.storage[158] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1590]$_SDFFE_PN0P_  (.CLK(clknet_leaf_141_clk_p2c),
    .RESET_B(net1534),
    .D(_00758_),
    .Q_N(_06209_),
    .Q(\shift_storage.storage[1590] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1591]$_SDFFE_PN0P_  (.CLK(clknet_leaf_141_clk_p2c),
    .RESET_B(net1535),
    .D(_00759_),
    .Q_N(_06208_),
    .Q(\shift_storage.storage[1591] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1592]$_SDFFE_PN0P_  (.CLK(clknet_leaf_141_clk_p2c),
    .RESET_B(net1536),
    .D(_00760_),
    .Q_N(_06207_),
    .Q(\shift_storage.storage[1592] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1593]$_SDFFE_PN0P_  (.CLK(clknet_leaf_141_clk_p2c),
    .RESET_B(net1537),
    .D(_00761_),
    .Q_N(_06206_),
    .Q(\shift_storage.storage[1593] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1594]$_SDFFE_PN0P_  (.CLK(clknet_leaf_141_clk_p2c),
    .RESET_B(net1538),
    .D(_00762_),
    .Q_N(_06205_),
    .Q(\shift_storage.storage[1594] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1595]$_SDFFE_PN0P_  (.CLK(clknet_leaf_140_clk_p2c),
    .RESET_B(net1539),
    .D(_00763_),
    .Q_N(_06204_),
    .Q(\shift_storage.storage[1595] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1596]$_SDFFE_PN0P_  (.CLK(clknet_leaf_140_clk_p2c),
    .RESET_B(net1540),
    .D(_00764_),
    .Q_N(_06203_),
    .Q(\shift_storage.storage[1596] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1597]$_SDFFE_PN0P_  (.CLK(clknet_leaf_140_clk_p2c),
    .RESET_B(net1541),
    .D(_00765_),
    .Q_N(_06202_),
    .Q(\shift_storage.storage[1597] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1598]$_SDFFE_PN0P_  (.CLK(clknet_leaf_140_clk_p2c),
    .RESET_B(net1542),
    .D(_00766_),
    .Q_N(_06201_),
    .Q(\shift_storage.storage[1598] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1599]$_SDFFE_PN0P_  (.CLK(clknet_leaf_139_clk_p2c),
    .RESET_B(net1543),
    .D(_00767_),
    .Q_N(_06200_),
    .Q(\shift_storage.shreg_out ));
 sg13g2_dfrbp_1 \shift_storage.storage[159]$_SDFFE_PN0P_  (.CLK(clknet_leaf_49_clk_p2c),
    .RESET_B(net1544),
    .D(_00768_),
    .Q_N(_06199_),
    .Q(\shift_storage.storage[159] ));
 sg13g2_dfrbp_1 \shift_storage.storage[15]$_SDFFE_PN0P_  (.CLK(clknet_leaf_69_clk_p2c),
    .RESET_B(net1545),
    .D(_00769_),
    .Q_N(_06198_),
    .Q(\shift_storage.storage[15] ));
 sg13g2_dfrbp_1 \shift_storage.storage[160]$_SDFFE_PN0P_  (.CLK(clknet_leaf_46_clk_p2c),
    .RESET_B(net1546),
    .D(_00770_),
    .Q_N(_06197_),
    .Q(\shift_storage.storage[160] ));
 sg13g2_dfrbp_1 \shift_storage.storage[161]$_SDFFE_PN0P_  (.CLK(clknet_leaf_49_clk_p2c),
    .RESET_B(net1547),
    .D(_00771_),
    .Q_N(_06196_),
    .Q(\shift_storage.storage[161] ));
 sg13g2_dfrbp_1 \shift_storage.storage[162]$_SDFFE_PN0P_  (.CLK(clknet_leaf_49_clk_p2c),
    .RESET_B(net1548),
    .D(_00772_),
    .Q_N(_06195_),
    .Q(\shift_storage.storage[162] ));
 sg13g2_dfrbp_1 \shift_storage.storage[163]$_SDFFE_PN0P_  (.CLK(clknet_leaf_52_clk_p2c),
    .RESET_B(net1549),
    .D(_00773_),
    .Q_N(_06194_),
    .Q(\shift_storage.storage[163] ));
 sg13g2_dfrbp_1 \shift_storage.storage[164]$_SDFFE_PN0P_  (.CLK(clknet_leaf_52_clk_p2c),
    .RESET_B(net1550),
    .D(_00774_),
    .Q_N(_06193_),
    .Q(\shift_storage.storage[164] ));
 sg13g2_dfrbp_1 \shift_storage.storage[165]$_SDFFE_PN0P_  (.CLK(clknet_leaf_52_clk_p2c),
    .RESET_B(net1551),
    .D(_00775_),
    .Q_N(_06192_),
    .Q(\shift_storage.storage[165] ));
 sg13g2_dfrbp_1 \shift_storage.storage[166]$_SDFFE_PN0P_  (.CLK(clknet_leaf_51_clk_p2c),
    .RESET_B(net1552),
    .D(_00776_),
    .Q_N(_06191_),
    .Q(\shift_storage.storage[166] ));
 sg13g2_dfrbp_1 \shift_storage.storage[167]$_SDFFE_PN0P_  (.CLK(clknet_leaf_51_clk_p2c),
    .RESET_B(net1553),
    .D(_00777_),
    .Q_N(_06190_),
    .Q(\shift_storage.storage[167] ));
 sg13g2_dfrbp_1 \shift_storage.storage[168]$_SDFFE_PN0P_  (.CLK(clknet_leaf_51_clk_p2c),
    .RESET_B(net1554),
    .D(_00778_),
    .Q_N(_06189_),
    .Q(\shift_storage.storage[168] ));
 sg13g2_dfrbp_1 \shift_storage.storage[169]$_SDFFE_PN0P_  (.CLK(clknet_leaf_51_clk_p2c),
    .RESET_B(net1555),
    .D(_00779_),
    .Q_N(_06188_),
    .Q(\shift_storage.storage[169] ));
 sg13g2_dfrbp_1 \shift_storage.storage[16]$_SDFFE_PN0P_  (.CLK(clknet_leaf_68_clk_p2c),
    .RESET_B(net1556),
    .D(_00780_),
    .Q_N(_06187_),
    .Q(\shift_storage.storage[16] ));
 sg13g2_dfrbp_1 \shift_storage.storage[170]$_SDFFE_PN0P_  (.CLK(clknet_leaf_52_clk_p2c),
    .RESET_B(net1557),
    .D(_00781_),
    .Q_N(_06186_),
    .Q(\shift_storage.storage[170] ));
 sg13g2_dfrbp_1 \shift_storage.storage[171]$_SDFFE_PN0P_  (.CLK(clknet_leaf_52_clk_p2c),
    .RESET_B(net1558),
    .D(_00782_),
    .Q_N(_06185_),
    .Q(\shift_storage.storage[171] ));
 sg13g2_dfrbp_1 \shift_storage.storage[172]$_SDFFE_PN0P_  (.CLK(clknet_leaf_53_clk_p2c),
    .RESET_B(net1559),
    .D(_00783_),
    .Q_N(_06184_),
    .Q(\shift_storage.storage[172] ));
 sg13g2_dfrbp_1 \shift_storage.storage[173]$_SDFFE_PN0P_  (.CLK(clknet_leaf_53_clk_p2c),
    .RESET_B(net1560),
    .D(_00784_),
    .Q_N(_06183_),
    .Q(\shift_storage.storage[173] ));
 sg13g2_dfrbp_1 \shift_storage.storage[174]$_SDFFE_PN0P_  (.CLK(clknet_leaf_53_clk_p2c),
    .RESET_B(net1561),
    .D(_00785_),
    .Q_N(_06182_),
    .Q(\shift_storage.storage[174] ));
 sg13g2_dfrbp_1 \shift_storage.storage[175]$_SDFFE_PN0P_  (.CLK(clknet_leaf_53_clk_p2c),
    .RESET_B(net1562),
    .D(_00786_),
    .Q_N(_06181_),
    .Q(\shift_storage.storage[175] ));
 sg13g2_dfrbp_1 \shift_storage.storage[176]$_SDFFE_PN0P_  (.CLK(clknet_leaf_53_clk_p2c),
    .RESET_B(net1563),
    .D(_00787_),
    .Q_N(_06180_),
    .Q(\shift_storage.storage[176] ));
 sg13g2_dfrbp_1 \shift_storage.storage[177]$_SDFFE_PN0P_  (.CLK(clknet_leaf_42_clk_p2c),
    .RESET_B(net1564),
    .D(_00788_),
    .Q_N(_06179_),
    .Q(\shift_storage.storage[177] ));
 sg13g2_dfrbp_1 \shift_storage.storage[178]$_SDFFE_PN0P_  (.CLK(clknet_leaf_53_clk_p2c),
    .RESET_B(net1565),
    .D(_00789_),
    .Q_N(_06178_),
    .Q(\shift_storage.storage[178] ));
 sg13g2_dfrbp_1 \shift_storage.storage[179]$_SDFFE_PN0P_  (.CLK(clknet_leaf_20_clk_p2c),
    .RESET_B(net1566),
    .D(_00790_),
    .Q_N(_06177_),
    .Q(\shift_storage.storage[179] ));
 sg13g2_dfrbp_1 \shift_storage.storage[17]$_SDFFE_PN0P_  (.CLK(clknet_leaf_68_clk_p2c),
    .RESET_B(net1567),
    .D(_00791_),
    .Q_N(_06176_),
    .Q(\shift_storage.storage[17] ));
 sg13g2_dfrbp_1 \shift_storage.storage[180]$_SDFFE_PN0P_  (.CLK(clknet_leaf_20_clk_p2c),
    .RESET_B(net1568),
    .D(_00792_),
    .Q_N(_06175_),
    .Q(\shift_storage.storage[180] ));
 sg13g2_dfrbp_1 \shift_storage.storage[181]$_SDFFE_PN0P_  (.CLK(clknet_leaf_20_clk_p2c),
    .RESET_B(net1569),
    .D(_00793_),
    .Q_N(_06174_),
    .Q(\shift_storage.storage[181] ));
 sg13g2_dfrbp_1 \shift_storage.storage[182]$_SDFFE_PN0P_  (.CLK(clknet_leaf_20_clk_p2c),
    .RESET_B(net1570),
    .D(_00794_),
    .Q_N(_06173_),
    .Q(\shift_storage.storage[182] ));
 sg13g2_dfrbp_1 \shift_storage.storage[183]$_SDFFE_PN0P_  (.CLK(clknet_leaf_19_clk_p2c),
    .RESET_B(net1571),
    .D(_00795_),
    .Q_N(_06172_),
    .Q(\shift_storage.storage[183] ));
 sg13g2_dfrbp_1 \shift_storage.storage[184]$_SDFFE_PN0P_  (.CLK(clknet_leaf_20_clk_p2c),
    .RESET_B(net1572),
    .D(_00796_),
    .Q_N(_06171_),
    .Q(\shift_storage.storage[184] ));
 sg13g2_dfrbp_1 \shift_storage.storage[185]$_SDFFE_PN0P_  (.CLK(clknet_leaf_19_clk_p2c),
    .RESET_B(net1573),
    .D(_00797_),
    .Q_N(_06170_),
    .Q(\shift_storage.storage[185] ));
 sg13g2_dfrbp_1 \shift_storage.storage[186]$_SDFFE_PN0P_  (.CLK(clknet_leaf_19_clk_p2c),
    .RESET_B(net1574),
    .D(_00798_),
    .Q_N(_06169_),
    .Q(\shift_storage.storage[186] ));
 sg13g2_dfrbp_1 \shift_storage.storage[187]$_SDFFE_PN0P_  (.CLK(clknet_leaf_19_clk_p2c),
    .RESET_B(net1575),
    .D(_00799_),
    .Q_N(_06168_),
    .Q(\shift_storage.storage[187] ));
 sg13g2_dfrbp_1 \shift_storage.storage[188]$_SDFFE_PN0P_  (.CLK(clknet_leaf_19_clk_p2c),
    .RESET_B(net1576),
    .D(_00800_),
    .Q_N(_06167_),
    .Q(\shift_storage.storage[188] ));
 sg13g2_dfrbp_1 \shift_storage.storage[189]$_SDFFE_PN0P_  (.CLK(clknet_leaf_19_clk_p2c),
    .RESET_B(net1577),
    .D(_00801_),
    .Q_N(_06166_),
    .Q(\shift_storage.storage[189] ));
 sg13g2_dfrbp_1 \shift_storage.storage[18]$_SDFFE_PN0P_  (.CLK(clknet_leaf_68_clk_p2c),
    .RESET_B(net1578),
    .D(_00802_),
    .Q_N(_06165_),
    .Q(\shift_storage.storage[18] ));
 sg13g2_dfrbp_1 \shift_storage.storage[190]$_SDFFE_PN0P_  (.CLK(clknet_leaf_54_clk_p2c),
    .RESET_B(net1579),
    .D(_00803_),
    .Q_N(_06164_),
    .Q(\shift_storage.storage[190] ));
 sg13g2_dfrbp_1 \shift_storage.storage[191]$_SDFFE_PN0P_  (.CLK(clknet_leaf_54_clk_p2c),
    .RESET_B(net1580),
    .D(_00804_),
    .Q_N(_06163_),
    .Q(\shift_storage.storage[191] ));
 sg13g2_dfrbp_1 \shift_storage.storage[192]$_SDFFE_PN0P_  (.CLK(clknet_leaf_54_clk_p2c),
    .RESET_B(net1581),
    .D(_00805_),
    .Q_N(_06162_),
    .Q(\shift_storage.storage[192] ));
 sg13g2_dfrbp_1 \shift_storage.storage[193]$_SDFFE_PN0P_  (.CLK(clknet_leaf_53_clk_p2c),
    .RESET_B(net1582),
    .D(_00806_),
    .Q_N(_06161_),
    .Q(\shift_storage.storage[193] ));
 sg13g2_dfrbp_1 \shift_storage.storage[194]$_SDFFE_PN0P_  (.CLK(clknet_leaf_54_clk_p2c),
    .RESET_B(net1583),
    .D(_00807_),
    .Q_N(_06160_),
    .Q(\shift_storage.storage[194] ));
 sg13g2_dfrbp_1 \shift_storage.storage[195]$_SDFFE_PN0P_  (.CLK(clknet_leaf_54_clk_p2c),
    .RESET_B(net1584),
    .D(_00808_),
    .Q_N(_06159_),
    .Q(\shift_storage.storage[195] ));
 sg13g2_dfrbp_1 \shift_storage.storage[196]$_SDFFE_PN0P_  (.CLK(clknet_leaf_55_clk_p2c),
    .RESET_B(net1585),
    .D(_00809_),
    .Q_N(_06158_),
    .Q(\shift_storage.storage[196] ));
 sg13g2_dfrbp_1 \shift_storage.storage[197]$_SDFFE_PN0P_  (.CLK(clknet_leaf_55_clk_p2c),
    .RESET_B(net1586),
    .D(_00810_),
    .Q_N(_06157_),
    .Q(\shift_storage.storage[197] ));
 sg13g2_dfrbp_1 \shift_storage.storage[198]$_SDFFE_PN0P_  (.CLK(clknet_leaf_55_clk_p2c),
    .RESET_B(net1587),
    .D(_00811_),
    .Q_N(_06156_),
    .Q(\shift_storage.storage[198] ));
 sg13g2_dfrbp_1 \shift_storage.storage[199]$_SDFFE_PN0P_  (.CLK(clknet_leaf_51_clk_p2c),
    .RESET_B(net1588),
    .D(_00812_),
    .Q_N(_06155_),
    .Q(\shift_storage.storage[199] ));
 sg13g2_dfrbp_1 \shift_storage.storage[19]$_SDFFE_PN0P_  (.CLK(clknet_leaf_68_clk_p2c),
    .RESET_B(net1589),
    .D(_00813_),
    .Q_N(_06154_),
    .Q(\shift_storage.storage[19] ));
 sg13g2_dfrbp_1 \shift_storage.storage[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_76_clk_p2c),
    .RESET_B(net1590),
    .D(_00814_),
    .Q_N(_06153_),
    .Q(\shift_storage.storage[1] ));
 sg13g2_dfrbp_1 \shift_storage.storage[200]$_SDFFE_PN0P_  (.CLK(clknet_leaf_51_clk_p2c),
    .RESET_B(net1591),
    .D(_00815_),
    .Q_N(_06152_),
    .Q(\shift_storage.storage[200] ));
 sg13g2_dfrbp_1 \shift_storage.storage[201]$_SDFFE_PN0P_  (.CLK(clknet_leaf_50_clk_p2c),
    .RESET_B(net1592),
    .D(_00816_),
    .Q_N(_06151_),
    .Q(\shift_storage.storage[201] ));
 sg13g2_dfrbp_1 \shift_storage.storage[202]$_SDFFE_PN0P_  (.CLK(clknet_leaf_50_clk_p2c),
    .RESET_B(net1593),
    .D(_00817_),
    .Q_N(_06150_),
    .Q(\shift_storage.storage[202] ));
 sg13g2_dfrbp_1 \shift_storage.storage[203]$_SDFFE_PN0P_  (.CLK(clknet_leaf_50_clk_p2c),
    .RESET_B(net1594),
    .D(_00818_),
    .Q_N(_06149_),
    .Q(\shift_storage.storage[203] ));
 sg13g2_dfrbp_1 \shift_storage.storage[204]$_SDFFE_PN0P_  (.CLK(clknet_leaf_50_clk_p2c),
    .RESET_B(net1595),
    .D(_00819_),
    .Q_N(_06148_),
    .Q(\shift_storage.storage[204] ));
 sg13g2_dfrbp_1 \shift_storage.storage[205]$_SDFFE_PN0P_  (.CLK(clknet_leaf_66_clk_p2c),
    .RESET_B(net1596),
    .D(_00820_),
    .Q_N(_06147_),
    .Q(\shift_storage.storage[205] ));
 sg13g2_dfrbp_1 \shift_storage.storage[206]$_SDFFE_PN0P_  (.CLK(clknet_leaf_65_clk_p2c),
    .RESET_B(net1597),
    .D(_00821_),
    .Q_N(_06146_),
    .Q(\shift_storage.storage[206] ));
 sg13g2_dfrbp_1 \shift_storage.storage[207]$_SDFFE_PN0P_  (.CLK(clknet_leaf_65_clk_p2c),
    .RESET_B(net1598),
    .D(_00822_),
    .Q_N(_06145_),
    .Q(\shift_storage.storage[207] ));
 sg13g2_dfrbp_1 \shift_storage.storage[208]$_SDFFE_PN0P_  (.CLK(clknet_leaf_65_clk_p2c),
    .RESET_B(net1599),
    .D(_00823_),
    .Q_N(_06144_),
    .Q(\shift_storage.storage[208] ));
 sg13g2_dfrbp_1 \shift_storage.storage[209]$_SDFFE_PN0P_  (.CLK(clknet_leaf_62_clk_p2c),
    .RESET_B(net1600),
    .D(_00824_),
    .Q_N(_06143_),
    .Q(\shift_storage.storage[209] ));
 sg13g2_dfrbp_1 \shift_storage.storage[20]$_SDFFE_PN0P_  (.CLK(clknet_leaf_68_clk_p2c),
    .RESET_B(net1601),
    .D(_00825_),
    .Q_N(_06142_),
    .Q(\shift_storage.storage[20] ));
 sg13g2_dfrbp_1 \shift_storage.storage[210]$_SDFFE_PN0P_  (.CLK(clknet_leaf_62_clk_p2c),
    .RESET_B(net1602),
    .D(_00826_),
    .Q_N(_06141_),
    .Q(\shift_storage.storage[210] ));
 sg13g2_dfrbp_1 \shift_storage.storage[211]$_SDFFE_PN0P_  (.CLK(clknet_leaf_62_clk_p2c),
    .RESET_B(net1603),
    .D(_00827_),
    .Q_N(_06140_),
    .Q(\shift_storage.storage[211] ));
 sg13g2_dfrbp_1 \shift_storage.storage[212]$_SDFFE_PN0P_  (.CLK(clknet_leaf_61_clk_p2c),
    .RESET_B(net1604),
    .D(_00828_),
    .Q_N(_06139_),
    .Q(\shift_storage.storage[212] ));
 sg13g2_dfrbp_1 \shift_storage.storage[213]$_SDFFE_PN0P_  (.CLK(clknet_leaf_61_clk_p2c),
    .RESET_B(net1605),
    .D(_00829_),
    .Q_N(_06138_),
    .Q(\shift_storage.storage[213] ));
 sg13g2_dfrbp_1 \shift_storage.storage[214]$_SDFFE_PN0P_  (.CLK(clknet_leaf_61_clk_p2c),
    .RESET_B(net1606),
    .D(_00830_),
    .Q_N(_06137_),
    .Q(\shift_storage.storage[214] ));
 sg13g2_dfrbp_1 \shift_storage.storage[215]$_SDFFE_PN0P_  (.CLK(clknet_leaf_61_clk_p2c),
    .RESET_B(net1607),
    .D(_00831_),
    .Q_N(_06136_),
    .Q(\shift_storage.storage[215] ));
 sg13g2_dfrbp_1 \shift_storage.storage[216]$_SDFFE_PN0P_  (.CLK(clknet_leaf_56_clk_p2c),
    .RESET_B(net1608),
    .D(_00832_),
    .Q_N(_06135_),
    .Q(\shift_storage.storage[216] ));
 sg13g2_dfrbp_1 \shift_storage.storage[217]$_SDFFE_PN0P_  (.CLK(clknet_leaf_56_clk_p2c),
    .RESET_B(net1609),
    .D(_00833_),
    .Q_N(_06134_),
    .Q(\shift_storage.storage[217] ));
 sg13g2_dfrbp_1 \shift_storage.storage[218]$_SDFFE_PN0P_  (.CLK(clknet_leaf_57_clk_p2c),
    .RESET_B(net1610),
    .D(_00834_),
    .Q_N(_06133_),
    .Q(\shift_storage.storage[218] ));
 sg13g2_dfrbp_1 \shift_storage.storage[219]$_SDFFE_PN0P_  (.CLK(clknet_leaf_57_clk_p2c),
    .RESET_B(net1611),
    .D(_00835_),
    .Q_N(_06132_),
    .Q(\shift_storage.storage[219] ));
 sg13g2_dfrbp_1 \shift_storage.storage[21]$_SDFFE_PN0P_  (.CLK(clknet_leaf_67_clk_p2c),
    .RESET_B(net1612),
    .D(_00836_),
    .Q_N(_06131_),
    .Q(\shift_storage.storage[21] ));
 sg13g2_dfrbp_1 \shift_storage.storage[220]$_SDFFE_PN0P_  (.CLK(clknet_leaf_58_clk_p2c),
    .RESET_B(net1613),
    .D(_00837_),
    .Q_N(_06130_),
    .Q(\shift_storage.storage[220] ));
 sg13g2_dfrbp_1 \shift_storage.storage[221]$_SDFFE_PN0P_  (.CLK(clknet_leaf_58_clk_p2c),
    .RESET_B(net1614),
    .D(_00838_),
    .Q_N(_06129_),
    .Q(\shift_storage.storage[221] ));
 sg13g2_dfrbp_1 \shift_storage.storage[222]$_SDFFE_PN0P_  (.CLK(clknet_leaf_58_clk_p2c),
    .RESET_B(net1615),
    .D(_00839_),
    .Q_N(_06128_),
    .Q(\shift_storage.storage[222] ));
 sg13g2_dfrbp_1 \shift_storage.storage[223]$_SDFFE_PN0P_  (.CLK(clknet_leaf_58_clk_p2c),
    .RESET_B(net1616),
    .D(_00840_),
    .Q_N(_06127_),
    .Q(\shift_storage.storage[223] ));
 sg13g2_dfrbp_1 \shift_storage.storage[224]$_SDFFE_PN0P_  (.CLK(clknet_leaf_58_clk_p2c),
    .RESET_B(net1617),
    .D(_00841_),
    .Q_N(_06126_),
    .Q(\shift_storage.storage[224] ));
 sg13g2_dfrbp_1 \shift_storage.storage[225]$_SDFFE_PN0P_  (.CLK(clknet_leaf_15_clk_p2c),
    .RESET_B(net1618),
    .D(_00842_),
    .Q_N(_06125_),
    .Q(\shift_storage.storage[225] ));
 sg13g2_dfrbp_1 \shift_storage.storage[226]$_SDFFE_PN0P_  (.CLK(clknet_leaf_15_clk_p2c),
    .RESET_B(net1619),
    .D(_00843_),
    .Q_N(_06124_),
    .Q(\shift_storage.storage[226] ));
 sg13g2_dfrbp_1 \shift_storage.storage[227]$_SDFFE_PN0P_  (.CLK(clknet_leaf_15_clk_p2c),
    .RESET_B(net1620),
    .D(_00844_),
    .Q_N(_06123_),
    .Q(\shift_storage.storage[227] ));
 sg13g2_dfrbp_1 \shift_storage.storage[228]$_SDFFE_PN0P_  (.CLK(clknet_leaf_16_clk_p2c),
    .RESET_B(net1621),
    .D(_00845_),
    .Q_N(_06122_),
    .Q(\shift_storage.storage[228] ));
 sg13g2_dfrbp_1 \shift_storage.storage[229]$_SDFFE_PN0P_  (.CLK(clknet_leaf_16_clk_p2c),
    .RESET_B(net1622),
    .D(_00846_),
    .Q_N(_06121_),
    .Q(\shift_storage.storage[229] ));
 sg13g2_dfrbp_1 \shift_storage.storage[22]$_SDFFE_PN0P_  (.CLK(clknet_leaf_67_clk_p2c),
    .RESET_B(net1623),
    .D(_00847_),
    .Q_N(_06120_),
    .Q(\shift_storage.storage[22] ));
 sg13g2_dfrbp_1 \shift_storage.storage[230]$_SDFFE_PN0P_  (.CLK(clknet_leaf_17_clk_p2c),
    .RESET_B(net1624),
    .D(_00848_),
    .Q_N(_06119_),
    .Q(\shift_storage.storage[230] ));
 sg13g2_dfrbp_1 \shift_storage.storage[231]$_SDFFE_PN0P_  (.CLK(clknet_leaf_15_clk_p2c),
    .RESET_B(net1625),
    .D(_00849_),
    .Q_N(_06118_),
    .Q(\shift_storage.storage[231] ));
 sg13g2_dfrbp_1 \shift_storage.storage[232]$_SDFFE_PN0P_  (.CLK(clknet_leaf_13_clk_p2c),
    .RESET_B(net1626),
    .D(_00850_),
    .Q_N(_06117_),
    .Q(\shift_storage.storage[232] ));
 sg13g2_dfrbp_1 \shift_storage.storage[233]$_SDFFE_PN0P_  (.CLK(clknet_leaf_13_clk_p2c),
    .RESET_B(net1627),
    .D(_00851_),
    .Q_N(_06116_),
    .Q(\shift_storage.storage[233] ));
 sg13g2_dfrbp_1 \shift_storage.storage[234]$_SDFFE_PN0P_  (.CLK(clknet_leaf_14_clk_p2c),
    .RESET_B(net1628),
    .D(_00852_),
    .Q_N(_06115_),
    .Q(\shift_storage.storage[234] ));
 sg13g2_dfrbp_1 \shift_storage.storage[235]$_SDFFE_PN0P_  (.CLK(clknet_leaf_13_clk_p2c),
    .RESET_B(net1629),
    .D(_00853_),
    .Q_N(_06114_),
    .Q(\shift_storage.storage[235] ));
 sg13g2_dfrbp_1 \shift_storage.storage[236]$_SDFFE_PN0P_  (.CLK(clknet_leaf_14_clk_p2c),
    .RESET_B(net1630),
    .D(_00854_),
    .Q_N(_06113_),
    .Q(\shift_storage.storage[236] ));
 sg13g2_dfrbp_1 \shift_storage.storage[237]$_SDFFE_PN0P_  (.CLK(clknet_leaf_14_clk_p2c),
    .RESET_B(net1631),
    .D(_00855_),
    .Q_N(_06112_),
    .Q(\shift_storage.storage[237] ));
 sg13g2_dfrbp_1 \shift_storage.storage[238]$_SDFFE_PN0P_  (.CLK(clknet_leaf_14_clk_p2c),
    .RESET_B(net1632),
    .D(_00856_),
    .Q_N(_06111_),
    .Q(\shift_storage.storage[238] ));
 sg13g2_dfrbp_1 \shift_storage.storage[239]$_SDFFE_PN0P_  (.CLK(clknet_leaf_14_clk_p2c),
    .RESET_B(net1633),
    .D(_00857_),
    .Q_N(_06110_),
    .Q(\shift_storage.storage[239] ));
 sg13g2_dfrbp_1 \shift_storage.storage[23]$_SDFFE_PN0P_  (.CLK(clknet_leaf_67_clk_p2c),
    .RESET_B(net1634),
    .D(_00858_),
    .Q_N(_06109_),
    .Q(\shift_storage.storage[23] ));
 sg13g2_dfrbp_1 \shift_storage.storage[240]$_SDFFE_PN0P_  (.CLK(clknet_leaf_14_clk_p2c),
    .RESET_B(net1635),
    .D(_00859_),
    .Q_N(_06108_),
    .Q(\shift_storage.storage[240] ));
 sg13g2_dfrbp_1 \shift_storage.storage[241]$_SDFFE_PN0P_  (.CLK(clknet_leaf_59_clk_p2c),
    .RESET_B(net1636),
    .D(_00860_),
    .Q_N(_06107_),
    .Q(\shift_storage.storage[241] ));
 sg13g2_dfrbp_1 \shift_storage.storage[242]$_SDFFE_PN0P_  (.CLK(clknet_leaf_59_clk_p2c),
    .RESET_B(net1637),
    .D(_00861_),
    .Q_N(_06106_),
    .Q(\shift_storage.storage[242] ));
 sg13g2_dfrbp_1 \shift_storage.storage[243]$_SDFFE_PN0P_  (.CLK(clknet_leaf_15_clk_p2c),
    .RESET_B(net1638),
    .D(_00862_),
    .Q_N(_06105_),
    .Q(\shift_storage.storage[243] ));
 sg13g2_dfrbp_1 \shift_storage.storage[244]$_SDFFE_PN0P_  (.CLK(clknet_leaf_58_clk_p2c),
    .RESET_B(net1639),
    .D(_00863_),
    .Q_N(_06104_),
    .Q(\shift_storage.storage[244] ));
 sg13g2_dfrbp_1 \shift_storage.storage[245]$_SDFFE_PN0P_  (.CLK(clknet_leaf_59_clk_p2c),
    .RESET_B(net1640),
    .D(_00864_),
    .Q_N(_06103_),
    .Q(\shift_storage.storage[245] ));
 sg13g2_dfrbp_1 \shift_storage.storage[246]$_SDFFE_PN0P_  (.CLK(clknet_leaf_59_clk_p2c),
    .RESET_B(net1641),
    .D(_00865_),
    .Q_N(_06102_),
    .Q(\shift_storage.storage[246] ));
 sg13g2_dfrbp_1 \shift_storage.storage[247]$_SDFFE_PN0P_  (.CLK(clknet_leaf_59_clk_p2c),
    .RESET_B(net1642),
    .D(_00866_),
    .Q_N(_06101_),
    .Q(\shift_storage.storage[247] ));
 sg13g2_dfrbp_1 \shift_storage.storage[248]$_SDFFE_PN0P_  (.CLK(clknet_leaf_60_clk_p2c),
    .RESET_B(net1643),
    .D(_00867_),
    .Q_N(_06100_),
    .Q(\shift_storage.storage[248] ));
 sg13g2_dfrbp_1 \shift_storage.storage[249]$_SDFFE_PN0P_  (.CLK(clknet_leaf_60_clk_p2c),
    .RESET_B(net1644),
    .D(_00868_),
    .Q_N(_06099_),
    .Q(\shift_storage.storage[249] ));
 sg13g2_dfrbp_1 \shift_storage.storage[24]$_SDFFE_PN0P_  (.CLK(clknet_leaf_67_clk_p2c),
    .RESET_B(net1645),
    .D(_00869_),
    .Q_N(_06098_),
    .Q(\shift_storage.storage[24] ));
 sg13g2_dfrbp_1 \shift_storage.storage[250]$_SDFFE_PN0P_  (.CLK(clknet_leaf_60_clk_p2c),
    .RESET_B(net1646),
    .D(_00870_),
    .Q_N(_06097_),
    .Q(\shift_storage.storage[250] ));
 sg13g2_dfrbp_1 \shift_storage.storage[251]$_SDFFE_PN0P_  (.CLK(clknet_leaf_60_clk_p2c),
    .RESET_B(net1647),
    .D(_00871_),
    .Q_N(_06096_),
    .Q(\shift_storage.storage[251] ));
 sg13g2_dfrbp_1 \shift_storage.storage[252]$_SDFFE_PN0P_  (.CLK(clknet_leaf_61_clk_p2c),
    .RESET_B(net1648),
    .D(_00872_),
    .Q_N(_06095_),
    .Q(\shift_storage.storage[252] ));
 sg13g2_dfrbp_1 \shift_storage.storage[253]$_SDFFE_PN0P_  (.CLK(clknet_leaf_60_clk_p2c),
    .RESET_B(net1649),
    .D(_00873_),
    .Q_N(_06094_),
    .Q(\shift_storage.storage[253] ));
 sg13g2_dfrbp_1 \shift_storage.storage[254]$_SDFFE_PN0P_  (.CLK(clknet_leaf_60_clk_p2c),
    .RESET_B(net1650),
    .D(_00874_),
    .Q_N(_06093_),
    .Q(\shift_storage.storage[254] ));
 sg13g2_dfrbp_1 \shift_storage.storage[255]$_SDFFE_PN0P_  (.CLK(clknet_leaf_61_clk_p2c),
    .RESET_B(net1651),
    .D(_00875_),
    .Q_N(_06092_),
    .Q(\shift_storage.storage[255] ));
 sg13g2_dfrbp_1 \shift_storage.storage[256]$_SDFFE_PN0P_  (.CLK(clknet_leaf_62_clk_p2c),
    .RESET_B(net1652),
    .D(_00876_),
    .Q_N(_06091_),
    .Q(\shift_storage.storage[256] ));
 sg13g2_dfrbp_1 \shift_storage.storage[257]$_SDFFE_PN0P_  (.CLK(clknet_leaf_63_clk_p2c),
    .RESET_B(net1653),
    .D(_00877_),
    .Q_N(_06090_),
    .Q(\shift_storage.storage[257] ));
 sg13g2_dfrbp_1 \shift_storage.storage[258]$_SDFFE_PN0P_  (.CLK(clknet_leaf_62_clk_p2c),
    .RESET_B(net1654),
    .D(_00878_),
    .Q_N(_06089_),
    .Q(\shift_storage.storage[258] ));
 sg13g2_dfrbp_1 \shift_storage.storage[259]$_SDFFE_PN0P_  (.CLK(clknet_leaf_62_clk_p2c),
    .RESET_B(net1655),
    .D(_00879_),
    .Q_N(_06088_),
    .Q(\shift_storage.storage[259] ));
 sg13g2_dfrbp_1 \shift_storage.storage[25]$_SDFFE_PN0P_  (.CLK(clknet_leaf_67_clk_p2c),
    .RESET_B(net1656),
    .D(_00880_),
    .Q_N(_06087_),
    .Q(\shift_storage.storage[25] ));
 sg13g2_dfrbp_1 \shift_storage.storage[260]$_SDFFE_PN0P_  (.CLK(clknet_leaf_63_clk_p2c),
    .RESET_B(net1657),
    .D(_00881_),
    .Q_N(_06086_),
    .Q(\shift_storage.storage[260] ));
 sg13g2_dfrbp_1 \shift_storage.storage[261]$_SDFFE_PN0P_  (.CLK(clknet_leaf_63_clk_p2c),
    .RESET_B(net1658),
    .D(_00882_),
    .Q_N(_06085_),
    .Q(\shift_storage.storage[261] ));
 sg13g2_dfrbp_1 \shift_storage.storage[262]$_SDFFE_PN0P_  (.CLK(clknet_leaf_64_clk_p2c),
    .RESET_B(net1659),
    .D(_00883_),
    .Q_N(_06084_),
    .Q(\shift_storage.storage[262] ));
 sg13g2_dfrbp_1 \shift_storage.storage[263]$_SDFFE_PN0P_  (.CLK(clknet_leaf_63_clk_p2c),
    .RESET_B(net1660),
    .D(_00884_),
    .Q_N(_06083_),
    .Q(\shift_storage.storage[263] ));
 sg13g2_dfrbp_1 \shift_storage.storage[264]$_SDFFE_PN0P_  (.CLK(clknet_leaf_64_clk_p2c),
    .RESET_B(net1661),
    .D(_00885_),
    .Q_N(_06082_),
    .Q(\shift_storage.storage[264] ));
 sg13g2_dfrbp_1 \shift_storage.storage[265]$_SDFFE_PN0P_  (.CLK(clknet_leaf_63_clk_p2c),
    .RESET_B(net1662),
    .D(_00886_),
    .Q_N(_06081_),
    .Q(\shift_storage.storage[265] ));
 sg13g2_dfrbp_1 \shift_storage.storage[266]$_SDFFE_PN0P_  (.CLK(clknet_leaf_64_clk_p2c),
    .RESET_B(net1663),
    .D(_00887_),
    .Q_N(_06080_),
    .Q(\shift_storage.storage[266] ));
 sg13g2_dfrbp_1 \shift_storage.storage[267]$_SDFFE_PN0P_  (.CLK(clknet_leaf_64_clk_p2c),
    .RESET_B(net1664),
    .D(_00888_),
    .Q_N(_06079_),
    .Q(\shift_storage.storage[267] ));
 sg13g2_dfrbp_1 \shift_storage.storage[268]$_SDFFE_PN0P_  (.CLK(clknet_leaf_64_clk_p2c),
    .RESET_B(net1665),
    .D(_00889_),
    .Q_N(_06078_),
    .Q(\shift_storage.storage[268] ));
 sg13g2_dfrbp_1 \shift_storage.storage[269]$_SDFFE_PN0P_  (.CLK(clknet_leaf_71_clk_p2c),
    .RESET_B(net1666),
    .D(_00890_),
    .Q_N(_06077_),
    .Q(\shift_storage.storage[269] ));
 sg13g2_dfrbp_1 \shift_storage.storage[26]$_SDFFE_PN0P_  (.CLK(clknet_leaf_49_clk_p2c),
    .RESET_B(net1667),
    .D(_00891_),
    .Q_N(_06076_),
    .Q(\shift_storage.storage[26] ));
 sg13g2_dfrbp_1 \shift_storage.storage[270]$_SDFFE_PN0P_  (.CLK(clknet_leaf_71_clk_p2c),
    .RESET_B(net1668),
    .D(_00892_),
    .Q_N(_06075_),
    .Q(\shift_storage.storage[270] ));
 sg13g2_dfrbp_1 \shift_storage.storage[271]$_SDFFE_PN0P_  (.CLK(clknet_leaf_71_clk_p2c),
    .RESET_B(net1669),
    .D(_00893_),
    .Q_N(_06074_),
    .Q(\shift_storage.storage[271] ));
 sg13g2_dfrbp_1 \shift_storage.storage[272]$_SDFFE_PN0P_  (.CLK(clknet_leaf_72_clk_p2c),
    .RESET_B(net1670),
    .D(_00894_),
    .Q_N(_06073_),
    .Q(\shift_storage.storage[272] ));
 sg13g2_dfrbp_1 \shift_storage.storage[273]$_SDFFE_PN0P_  (.CLK(clknet_leaf_72_clk_p2c),
    .RESET_B(net1671),
    .D(_00895_),
    .Q_N(_06072_),
    .Q(\shift_storage.storage[273] ));
 sg13g2_dfrbp_1 \shift_storage.storage[274]$_SDFFE_PN0P_  (.CLK(clknet_leaf_72_clk_p2c),
    .RESET_B(net1672),
    .D(_00896_),
    .Q_N(_06071_),
    .Q(\shift_storage.storage[274] ));
 sg13g2_dfrbp_1 \shift_storage.storage[275]$_SDFFE_PN0P_  (.CLK(clknet_leaf_72_clk_p2c),
    .RESET_B(net1673),
    .D(_00897_),
    .Q_N(_06070_),
    .Q(\shift_storage.storage[275] ));
 sg13g2_dfrbp_1 \shift_storage.storage[276]$_SDFFE_PN0P_  (.CLK(clknet_leaf_73_clk_p2c),
    .RESET_B(net1674),
    .D(_00898_),
    .Q_N(_06069_),
    .Q(\shift_storage.storage[276] ));
 sg13g2_dfrbp_1 \shift_storage.storage[277]$_SDFFE_PN0P_  (.CLK(clknet_leaf_73_clk_p2c),
    .RESET_B(net1675),
    .D(_00899_),
    .Q_N(_06068_),
    .Q(\shift_storage.storage[277] ));
 sg13g2_dfrbp_1 \shift_storage.storage[278]$_SDFFE_PN0P_  (.CLK(clknet_leaf_73_clk_p2c),
    .RESET_B(net1676),
    .D(_00900_),
    .Q_N(_06067_),
    .Q(\shift_storage.storage[278] ));
 sg13g2_dfrbp_1 \shift_storage.storage[279]$_SDFFE_PN0P_  (.CLK(clknet_leaf_75_clk_p2c),
    .RESET_B(net1677),
    .D(_00901_),
    .Q_N(_06066_),
    .Q(\shift_storage.storage[279] ));
 sg13g2_dfrbp_1 \shift_storage.storage[27]$_SDFFE_PN0P_  (.CLK(clknet_leaf_49_clk_p2c),
    .RESET_B(net1678),
    .D(_00902_),
    .Q_N(_06065_),
    .Q(\shift_storage.storage[27] ));
 sg13g2_dfrbp_1 \shift_storage.storage[280]$_SDFFE_PN0P_  (.CLK(clknet_leaf_74_clk_p2c),
    .RESET_B(net1679),
    .D(_00903_),
    .Q_N(_06064_),
    .Q(\shift_storage.storage[280] ));
 sg13g2_dfrbp_1 \shift_storage.storage[281]$_SDFFE_PN0P_  (.CLK(clknet_leaf_74_clk_p2c),
    .RESET_B(net1680),
    .D(_00904_),
    .Q_N(_06063_),
    .Q(\shift_storage.storage[281] ));
 sg13g2_dfrbp_1 \shift_storage.storage[282]$_SDFFE_PN0P_  (.CLK(clknet_leaf_74_clk_p2c),
    .RESET_B(net1681),
    .D(_00905_),
    .Q_N(_06062_),
    .Q(\shift_storage.storage[282] ));
 sg13g2_dfrbp_1 \shift_storage.storage[283]$_SDFFE_PN0P_  (.CLK(clknet_leaf_74_clk_p2c),
    .RESET_B(net1682),
    .D(_00906_),
    .Q_N(_06061_),
    .Q(\shift_storage.storage[283] ));
 sg13g2_dfrbp_1 \shift_storage.storage[284]$_SDFFE_PN0P_  (.CLK(clknet_leaf_70_clk_p2c),
    .RESET_B(net1683),
    .D(_00907_),
    .Q_N(_06060_),
    .Q(\shift_storage.storage[284] ));
 sg13g2_dfrbp_1 \shift_storage.storage[285]$_SDFFE_PN0P_  (.CLK(clknet_leaf_69_clk_p2c),
    .RESET_B(net1684),
    .D(_00908_),
    .Q_N(_06059_),
    .Q(\shift_storage.storage[285] ));
 sg13g2_dfrbp_1 \shift_storage.storage[286]$_SDFFE_PN0P_  (.CLK(clknet_leaf_81_clk_p2c),
    .RESET_B(net1685),
    .D(_00909_),
    .Q_N(_06058_),
    .Q(\shift_storage.storage[286] ));
 sg13g2_dfrbp_1 \shift_storage.storage[287]$_SDFFE_PN0P_  (.CLK(clknet_leaf_81_clk_p2c),
    .RESET_B(net1686),
    .D(_00910_),
    .Q_N(_06057_),
    .Q(\shift_storage.storage[287] ));
 sg13g2_dfrbp_1 \shift_storage.storage[288]$_SDFFE_PN0P_  (.CLK(clknet_leaf_81_clk_p2c),
    .RESET_B(net1687),
    .D(_00911_),
    .Q_N(_06056_),
    .Q(\shift_storage.storage[288] ));
 sg13g2_dfrbp_1 \shift_storage.storage[289]$_SDFFE_PN0P_  (.CLK(clknet_leaf_81_clk_p2c),
    .RESET_B(net1688),
    .D(_00912_),
    .Q_N(_06055_),
    .Q(\shift_storage.storage[289] ));
 sg13g2_dfrbp_1 \shift_storage.storage[28]$_SDFFE_PN0P_  (.CLK(clknet_leaf_48_clk_p2c),
    .RESET_B(net1689),
    .D(_00913_),
    .Q_N(_06054_),
    .Q(\shift_storage.storage[28] ));
 sg13g2_dfrbp_1 \shift_storage.storage[290]$_SDFFE_PN0P_  (.CLK(clknet_leaf_81_clk_p2c),
    .RESET_B(net1690),
    .D(_00914_),
    .Q_N(_06053_),
    .Q(\shift_storage.storage[290] ));
 sg13g2_dfrbp_1 \shift_storage.storage[291]$_SDFFE_PN0P_  (.CLK(clknet_leaf_82_clk_p2c),
    .RESET_B(net1691),
    .D(_00915_),
    .Q_N(_06052_),
    .Q(\shift_storage.storage[291] ));
 sg13g2_dfrbp_1 \shift_storage.storage[292]$_SDFFE_PN0P_  (.CLK(clknet_leaf_82_clk_p2c),
    .RESET_B(net1692),
    .D(_00916_),
    .Q_N(_06051_),
    .Q(\shift_storage.storage[292] ));
 sg13g2_dfrbp_1 \shift_storage.storage[293]$_SDFFE_PN0P_  (.CLK(clknet_leaf_82_clk_p2c),
    .RESET_B(net1693),
    .D(_00917_),
    .Q_N(_06050_),
    .Q(\shift_storage.storage[293] ));
 sg13g2_dfrbp_1 \shift_storage.storage[294]$_SDFFE_PN0P_  (.CLK(clknet_leaf_82_clk_p2c),
    .RESET_B(net1694),
    .D(_00918_),
    .Q_N(_06049_),
    .Q(\shift_storage.storage[294] ));
 sg13g2_dfrbp_1 \shift_storage.storage[295]$_SDFFE_PN0P_  (.CLK(clknet_leaf_81_clk_p2c),
    .RESET_B(net1695),
    .D(_00919_),
    .Q_N(_06048_),
    .Q(\shift_storage.storage[295] ));
 sg13g2_dfrbp_1 \shift_storage.storage[296]$_SDFFE_PN0P_  (.CLK(clknet_leaf_69_clk_p2c),
    .RESET_B(net1696),
    .D(_00920_),
    .Q_N(_06047_),
    .Q(\shift_storage.storage[296] ));
 sg13g2_dfrbp_1 \shift_storage.storage[297]$_SDFFE_PN0P_  (.CLK(clknet_leaf_69_clk_p2c),
    .RESET_B(net1697),
    .D(_00921_),
    .Q_N(_06046_),
    .Q(\shift_storage.storage[297] ));
 sg13g2_dfrbp_1 \shift_storage.storage[298]$_SDFFE_PN0P_  (.CLK(clknet_leaf_69_clk_p2c),
    .RESET_B(net1698),
    .D(_00922_),
    .Q_N(_06045_),
    .Q(\shift_storage.storage[298] ));
 sg13g2_dfrbp_1 \shift_storage.storage[299]$_SDFFE_PN0P_  (.CLK(clknet_leaf_69_clk_p2c),
    .RESET_B(net1699),
    .D(_00923_),
    .Q_N(_06044_),
    .Q(\shift_storage.storage[299] ));
 sg13g2_dfrbp_1 \shift_storage.storage[29]$_SDFFE_PN0P_  (.CLK(clknet_leaf_48_clk_p2c),
    .RESET_B(net1700),
    .D(_00924_),
    .Q_N(_06043_),
    .Q(\shift_storage.storage[29] ));
 sg13g2_dfrbp_1 \shift_storage.storage[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_76_clk_p2c),
    .RESET_B(net1701),
    .D(_00925_),
    .Q_N(_06042_),
    .Q(\shift_storage.storage[2] ));
 sg13g2_dfrbp_1 \shift_storage.storage[300]$_SDFFE_PN0P_  (.CLK(clknet_leaf_71_clk_p2c),
    .RESET_B(net1702),
    .D(_00926_),
    .Q_N(_06041_),
    .Q(\shift_storage.storage[300] ));
 sg13g2_dfrbp_1 \shift_storage.storage[301]$_SDFFE_PN0P_  (.CLK(clknet_leaf_71_clk_p2c),
    .RESET_B(net1703),
    .D(_00927_),
    .Q_N(_06040_),
    .Q(\shift_storage.storage[301] ));
 sg13g2_dfrbp_1 \shift_storage.storage[302]$_SDFFE_PN0P_  (.CLK(clknet_leaf_71_clk_p2c),
    .RESET_B(net1704),
    .D(_00928_),
    .Q_N(_06039_),
    .Q(\shift_storage.storage[302] ));
 sg13g2_dfrbp_1 \shift_storage.storage[303]$_SDFFE_PN0P_  (.CLK(clknet_leaf_68_clk_p2c),
    .RESET_B(net1705),
    .D(_00929_),
    .Q_N(_06038_),
    .Q(\shift_storage.storage[303] ));
 sg13g2_dfrbp_1 \shift_storage.storage[304]$_SDFFE_PN0P_  (.CLK(clknet_leaf_68_clk_p2c),
    .RESET_B(net1706),
    .D(_00930_),
    .Q_N(_06037_),
    .Q(\shift_storage.storage[304] ));
 sg13g2_dfrbp_1 \shift_storage.storage[305]$_SDFFE_PN0P_  (.CLK(clknet_leaf_67_clk_p2c),
    .RESET_B(net1707),
    .D(_00931_),
    .Q_N(_06036_),
    .Q(\shift_storage.storage[305] ));
 sg13g2_dfrbp_1 \shift_storage.storage[306]$_SDFFE_PN0P_  (.CLK(clknet_leaf_66_clk_p2c),
    .RESET_B(net1708),
    .D(_00932_),
    .Q_N(_06035_),
    .Q(\shift_storage.storage[306] ));
 sg13g2_dfrbp_1 \shift_storage.storage[307]$_SDFFE_PN0P_  (.CLK(clknet_leaf_66_clk_p2c),
    .RESET_B(net1709),
    .D(_00933_),
    .Q_N(_06034_),
    .Q(\shift_storage.storage[307] ));
 sg13g2_dfrbp_1 \shift_storage.storage[308]$_SDFFE_PN0P_  (.CLK(clknet_leaf_66_clk_p2c),
    .RESET_B(net1710),
    .D(_00934_),
    .Q_N(_06033_),
    .Q(\shift_storage.storage[308] ));
 sg13g2_dfrbp_1 \shift_storage.storage[309]$_SDFFE_PN0P_  (.CLK(clknet_leaf_66_clk_p2c),
    .RESET_B(net1711),
    .D(_00935_),
    .Q_N(_06032_),
    .Q(\shift_storage.storage[309] ));
 sg13g2_dfrbp_1 \shift_storage.storage[30]$_SDFFE_PN0P_  (.CLK(clknet_leaf_48_clk_p2c),
    .RESET_B(net1712),
    .D(_00936_),
    .Q_N(_06031_),
    .Q(\shift_storage.storage[30] ));
 sg13g2_dfrbp_1 \shift_storage.storage[310]$_SDFFE_PN0P_  (.CLK(clknet_leaf_66_clk_p2c),
    .RESET_B(net1713),
    .D(_00937_),
    .Q_N(_06030_),
    .Q(\shift_storage.storage[310] ));
 sg13g2_dfrbp_1 \shift_storage.storage[311]$_SDFFE_PN0P_  (.CLK(clknet_leaf_65_clk_p2c),
    .RESET_B(net1714),
    .D(_00938_),
    .Q_N(_06029_),
    .Q(\shift_storage.storage[311] ));
 sg13g2_dfrbp_1 \shift_storage.storage[312]$_SDFFE_PN0P_  (.CLK(clknet_leaf_50_clk_p2c),
    .RESET_B(net1715),
    .D(_00939_),
    .Q_N(_06028_),
    .Q(\shift_storage.storage[312] ));
 sg13g2_dfrbp_1 \shift_storage.storage[313]$_SDFFE_PN0P_  (.CLK(clknet_leaf_65_clk_p2c),
    .RESET_B(net1716),
    .D(_00940_),
    .Q_N(_06027_),
    .Q(\shift_storage.storage[313] ));
 sg13g2_dfrbp_1 \shift_storage.storage[314]$_SDFFE_PN0P_  (.CLK(clknet_leaf_65_clk_p2c),
    .RESET_B(net1717),
    .D(_00941_),
    .Q_N(_06026_),
    .Q(\shift_storage.storage[314] ));
 sg13g2_dfrbp_1 \shift_storage.storage[315]$_SDFFE_PN0P_  (.CLK(clknet_leaf_50_clk_p2c),
    .RESET_B(net1718),
    .D(_00942_),
    .Q_N(_06025_),
    .Q(\shift_storage.storage[315] ));
 sg13g2_dfrbp_1 \shift_storage.storage[316]$_SDFFE_PN0P_  (.CLK(clknet_leaf_56_clk_p2c),
    .RESET_B(net1719),
    .D(_00943_),
    .Q_N(_06024_),
    .Q(\shift_storage.storage[316] ));
 sg13g2_dfrbp_1 \shift_storage.storage[317]$_SDFFE_PN0P_  (.CLK(clknet_leaf_56_clk_p2c),
    .RESET_B(net1720),
    .D(_00944_),
    .Q_N(_06023_),
    .Q(\shift_storage.storage[317] ));
 sg13g2_dfrbp_1 \shift_storage.storage[318]$_SDFFE_PN0P_  (.CLK(clknet_leaf_56_clk_p2c),
    .RESET_B(net1721),
    .D(_00945_),
    .Q_N(_06022_),
    .Q(\shift_storage.storage[318] ));
 sg13g2_dfrbp_1 \shift_storage.storage[319]$_SDFFE_PN0P_  (.CLK(clknet_leaf_56_clk_p2c),
    .RESET_B(net1722),
    .D(_00946_),
    .Q_N(_06021_),
    .Q(\shift_storage.storage[319] ));
 sg13g2_dfrbp_1 \shift_storage.storage[31]$_SDFFE_PN0P_  (.CLK(clknet_leaf_49_clk_p2c),
    .RESET_B(net1723),
    .D(_00947_),
    .Q_N(_06020_),
    .Q(\shift_storage.storage[31] ));
 sg13g2_dfrbp_1 \shift_storage.storage[320]$_SDFFE_PN0P_  (.CLK(clknet_leaf_55_clk_p2c),
    .RESET_B(net1724),
    .D(_00948_),
    .Q_N(_06019_),
    .Q(\shift_storage.storage[320] ));
 sg13g2_dfrbp_1 \shift_storage.storage[321]$_SDFFE_PN0P_  (.CLK(clknet_leaf_55_clk_p2c),
    .RESET_B(net1725),
    .D(_00949_),
    .Q_N(_06018_),
    .Q(\shift_storage.storage[321] ));
 sg13g2_dfrbp_1 \shift_storage.storage[322]$_SDFFE_PN0P_  (.CLK(clknet_leaf_55_clk_p2c),
    .RESET_B(net1726),
    .D(_00950_),
    .Q_N(_06017_),
    .Q(\shift_storage.storage[322] ));
 sg13g2_dfrbp_1 \shift_storage.storage[323]$_SDFFE_PN0P_  (.CLK(clknet_leaf_55_clk_p2c),
    .RESET_B(net1727),
    .D(_00951_),
    .Q_N(_06016_),
    .Q(\shift_storage.storage[323] ));
 sg13g2_dfrbp_1 \shift_storage.storage[324]$_SDFFE_PN0P_  (.CLK(clknet_leaf_57_clk_p2c),
    .RESET_B(net1728),
    .D(_00952_),
    .Q_N(_06015_),
    .Q(\shift_storage.storage[324] ));
 sg13g2_dfrbp_1 \shift_storage.storage[325]$_SDFFE_PN0P_  (.CLK(clknet_leaf_57_clk_p2c),
    .RESET_B(net1729),
    .D(_00953_),
    .Q_N(_06014_),
    .Q(\shift_storage.storage[325] ));
 sg13g2_dfrbp_1 \shift_storage.storage[326]$_SDFFE_PN0P_  (.CLK(clknet_leaf_57_clk_p2c),
    .RESET_B(net1730),
    .D(_00954_),
    .Q_N(_06013_),
    .Q(\shift_storage.storage[326] ));
 sg13g2_dfrbp_1 \shift_storage.storage[327]$_SDFFE_PN0P_  (.CLK(clknet_leaf_16_clk_p2c),
    .RESET_B(net1731),
    .D(_00955_),
    .Q_N(_06012_),
    .Q(\shift_storage.storage[327] ));
 sg13g2_dfrbp_1 \shift_storage.storage[328]$_SDFFE_PN0P_  (.CLK(clknet_leaf_15_clk_p2c),
    .RESET_B(net1732),
    .D(_00956_),
    .Q_N(_06011_),
    .Q(\shift_storage.storage[328] ));
 sg13g2_dfrbp_1 \shift_storage.storage[329]$_SDFFE_PN0P_  (.CLK(clknet_leaf_16_clk_p2c),
    .RESET_B(net1733),
    .D(_00957_),
    .Q_N(_06010_),
    .Q(\shift_storage.storage[329] ));
 sg13g2_dfrbp_1 \shift_storage.storage[32]$_SDFFE_PN0P_  (.CLK(clknet_leaf_47_clk_p2c),
    .RESET_B(net1734),
    .D(_00958_),
    .Q_N(_06009_),
    .Q(\shift_storage.storage[32] ));
 sg13g2_dfrbp_1 \shift_storage.storage[330]$_SDFFE_PN0P_  (.CLK(clknet_leaf_16_clk_p2c),
    .RESET_B(net1735),
    .D(_00959_),
    .Q_N(_06008_),
    .Q(\shift_storage.storage[330] ));
 sg13g2_dfrbp_1 \shift_storage.storage[331]$_SDFFE_PN0P_  (.CLK(clknet_leaf_18_clk_p2c),
    .RESET_B(net1736),
    .D(_00960_),
    .Q_N(_06007_),
    .Q(\shift_storage.storage[331] ));
 sg13g2_dfrbp_1 \shift_storage.storage[332]$_SDFFE_PN0P_  (.CLK(clknet_leaf_18_clk_p2c),
    .RESET_B(net1737),
    .D(_00961_),
    .Q_N(_06006_),
    .Q(\shift_storage.storage[332] ));
 sg13g2_dfrbp_1 \shift_storage.storage[333]$_SDFFE_PN0P_  (.CLK(clknet_leaf_18_clk_p2c),
    .RESET_B(net1738),
    .D(_00962_),
    .Q_N(_06005_),
    .Q(\shift_storage.storage[333] ));
 sg13g2_dfrbp_1 \shift_storage.storage[334]$_SDFFE_PN0P_  (.CLK(clknet_leaf_18_clk_p2c),
    .RESET_B(net1739),
    .D(_00963_),
    .Q_N(_06004_),
    .Q(\shift_storage.storage[334] ));
 sg13g2_dfrbp_1 \shift_storage.storage[335]$_SDFFE_PN0P_  (.CLK(clknet_leaf_18_clk_p2c),
    .RESET_B(net1740),
    .D(_00964_),
    .Q_N(_06003_),
    .Q(\shift_storage.storage[335] ));
 sg13g2_dfrbp_1 \shift_storage.storage[336]$_SDFFE_PN0P_  (.CLK(clknet_leaf_17_clk_p2c),
    .RESET_B(net1741),
    .D(_00965_),
    .Q_N(_06002_),
    .Q(\shift_storage.storage[336] ));
 sg13g2_dfrbp_1 \shift_storage.storage[337]$_SDFFE_PN0P_  (.CLK(clknet_leaf_17_clk_p2c),
    .RESET_B(net1742),
    .D(_00966_),
    .Q_N(_06001_),
    .Q(\shift_storage.storage[337] ));
 sg13g2_dfrbp_1 \shift_storage.storage[338]$_SDFFE_PN0P_  (.CLK(clknet_leaf_17_clk_p2c),
    .RESET_B(net1743),
    .D(_00967_),
    .Q_N(_06000_),
    .Q(\shift_storage.storage[338] ));
 sg13g2_dfrbp_1 \shift_storage.storage[339]$_SDFFE_PN0P_  (.CLK(clknet_leaf_17_clk_p2c),
    .RESET_B(net1744),
    .D(_00968_),
    .Q_N(_05999_),
    .Q(\shift_storage.storage[339] ));
 sg13g2_dfrbp_1 \shift_storage.storage[33]$_SDFFE_PN0P_  (.CLK(clknet_leaf_48_clk_p2c),
    .RESET_B(net1745),
    .D(_00969_),
    .Q_N(_05998_),
    .Q(\shift_storage.storage[33] ));
 sg13g2_dfrbp_1 \shift_storage.storage[340]$_SDFFE_PN0P_  (.CLK(clknet_leaf_17_clk_p2c),
    .RESET_B(net1746),
    .D(_00970_),
    .Q_N(_05997_),
    .Q(\shift_storage.storage[340] ));
 sg13g2_dfrbp_1 \shift_storage.storage[341]$_SDFFE_PN0P_  (.CLK(clknet_leaf_12_clk_p2c),
    .RESET_B(net1747),
    .D(_00971_),
    .Q_N(_05996_),
    .Q(\shift_storage.storage[341] ));
 sg13g2_dfrbp_1 \shift_storage.storage[342]$_SDFFE_PN0P_  (.CLK(clknet_leaf_12_clk_p2c),
    .RESET_B(net1748),
    .D(_00972_),
    .Q_N(_05995_),
    .Q(\shift_storage.storage[342] ));
 sg13g2_dfrbp_1 \shift_storage.storage[343]$_SDFFE_PN0P_  (.CLK(clknet_leaf_13_clk_p2c),
    .RESET_B(net1749),
    .D(_00973_),
    .Q_N(_05994_),
    .Q(\shift_storage.storage[343] ));
 sg13g2_dfrbp_1 \shift_storage.storage[344]$_SDFFE_PN0P_  (.CLK(clknet_leaf_13_clk_p2c),
    .RESET_B(net1750),
    .D(_00974_),
    .Q_N(_05993_),
    .Q(\shift_storage.storage[344] ));
 sg13g2_dfrbp_1 \shift_storage.storage[345]$_SDFFE_PN0P_  (.CLK(clknet_leaf_13_clk_p2c),
    .RESET_B(net1751),
    .D(_00975_),
    .Q_N(_05992_),
    .Q(\shift_storage.storage[345] ));
 sg13g2_dfrbp_1 \shift_storage.storage[346]$_SDFFE_PN0P_  (.CLK(clknet_leaf_11_clk_p2c),
    .RESET_B(net1752),
    .D(_00976_),
    .Q_N(_05991_),
    .Q(\shift_storage.storage[346] ));
 sg13g2_dfrbp_1 \shift_storage.storage[347]$_SDFFE_PN0P_  (.CLK(clknet_leaf_10_clk_p2c),
    .RESET_B(net1753),
    .D(_00977_),
    .Q_N(_05990_),
    .Q(\shift_storage.storage[347] ));
 sg13g2_dfrbp_1 \shift_storage.storage[348]$_SDFFE_PN0P_  (.CLK(clknet_leaf_10_clk_p2c),
    .RESET_B(net1754),
    .D(_00978_),
    .Q_N(_05989_),
    .Q(\shift_storage.storage[348] ));
 sg13g2_dfrbp_1 \shift_storage.storage[349]$_SDFFE_PN0P_  (.CLK(clknet_leaf_11_clk_p2c),
    .RESET_B(net1755),
    .D(_00979_),
    .Q_N(_05988_),
    .Q(\shift_storage.storage[349] ));
 sg13g2_dfrbp_1 \shift_storage.storage[34]$_SDFFE_PN0P_  (.CLK(clknet_leaf_97_clk_p2c),
    .RESET_B(net1756),
    .D(_00980_),
    .Q_N(_05987_),
    .Q(\shift_storage.storage[34] ));
 sg13g2_dfrbp_1 \shift_storage.storage[350]$_SDFFE_PN0P_  (.CLK(clknet_leaf_10_clk_p2c),
    .RESET_B(net1757),
    .D(_00981_),
    .Q_N(_05986_),
    .Q(\shift_storage.storage[350] ));
 sg13g2_dfrbp_1 \shift_storage.storage[351]$_SDFFE_PN0P_  (.CLK(clknet_leaf_10_clk_p2c),
    .RESET_B(net1758),
    .D(_00982_),
    .Q_N(_05985_),
    .Q(\shift_storage.storage[351] ));
 sg13g2_dfrbp_1 \shift_storage.storage[352]$_SDFFE_PN0P_  (.CLK(clknet_leaf_10_clk_p2c),
    .RESET_B(net1759),
    .D(_00983_),
    .Q_N(_05984_),
    .Q(\shift_storage.storage[352] ));
 sg13g2_dfrbp_1 \shift_storage.storage[353]$_SDFFE_PN0P_  (.CLK(clknet_leaf_10_clk_p2c),
    .RESET_B(net1760),
    .D(_00984_),
    .Q_N(_05983_),
    .Q(\shift_storage.storage[353] ));
 sg13g2_dfrbp_1 \shift_storage.storage[354]$_SDFFE_PN0P_  (.CLK(clknet_leaf_9_clk_p2c),
    .RESET_B(net1761),
    .D(_00985_),
    .Q_N(_05982_),
    .Q(\shift_storage.storage[354] ));
 sg13g2_dfrbp_1 \shift_storage.storage[355]$_SDFFE_PN0P_  (.CLK(clknet_leaf_9_clk_p2c),
    .RESET_B(net1762),
    .D(_00986_),
    .Q_N(_05981_),
    .Q(\shift_storage.storage[355] ));
 sg13g2_dfrbp_1 \shift_storage.storage[356]$_SDFFE_PN0P_  (.CLK(clknet_leaf_9_clk_p2c),
    .RESET_B(net1763),
    .D(_00987_),
    .Q_N(_05980_),
    .Q(\shift_storage.storage[356] ));
 sg13g2_dfrbp_1 \shift_storage.storage[357]$_SDFFE_PN0P_  (.CLK(clknet_leaf_9_clk_p2c),
    .RESET_B(net1764),
    .D(_00988_),
    .Q_N(_05979_),
    .Q(\shift_storage.storage[357] ));
 sg13g2_dfrbp_1 \shift_storage.storage[358]$_SDFFE_PN0P_  (.CLK(clknet_leaf_9_clk_p2c),
    .RESET_B(net1765),
    .D(_00989_),
    .Q_N(_05978_),
    .Q(\shift_storage.storage[358] ));
 sg13g2_dfrbp_1 \shift_storage.storage[359]$_SDFFE_PN0P_  (.CLK(clknet_leaf_9_clk_p2c),
    .RESET_B(net1766),
    .D(_00990_),
    .Q_N(_05977_),
    .Q(\shift_storage.storage[359] ));
 sg13g2_dfrbp_1 \shift_storage.storage[35]$_SDFFE_PN0P_  (.CLK(clknet_leaf_96_clk_p2c),
    .RESET_B(net1767),
    .D(_00991_),
    .Q_N(_05976_),
    .Q(\shift_storage.storage[35] ));
 sg13g2_dfrbp_1 \shift_storage.storage[360]$_SDFFE_PN0P_  (.CLK(clknet_leaf_8_clk_p2c),
    .RESET_B(net1768),
    .D(_00992_),
    .Q_N(_05975_),
    .Q(\shift_storage.storage[360] ));
 sg13g2_dfrbp_1 \shift_storage.storage[361]$_SDFFE_PN0P_  (.CLK(clknet_leaf_6_clk_p2c),
    .RESET_B(net1769),
    .D(_00993_),
    .Q_N(_05974_),
    .Q(\shift_storage.storage[361] ));
 sg13g2_dfrbp_1 \shift_storage.storage[362]$_SDFFE_PN0P_  (.CLK(clknet_leaf_6_clk_p2c),
    .RESET_B(net1770),
    .D(_00994_),
    .Q_N(_05973_),
    .Q(\shift_storage.storage[362] ));
 sg13g2_dfrbp_1 \shift_storage.storage[363]$_SDFFE_PN0P_  (.CLK(clknet_leaf_6_clk_p2c),
    .RESET_B(net1771),
    .D(_00995_),
    .Q_N(_05972_),
    .Q(\shift_storage.storage[363] ));
 sg13g2_dfrbp_1 \shift_storage.storage[364]$_SDFFE_PN0P_  (.CLK(clknet_leaf_6_clk_p2c),
    .RESET_B(net1772),
    .D(_00996_),
    .Q_N(_05971_),
    .Q(\shift_storage.storage[364] ));
 sg13g2_dfrbp_1 \shift_storage.storage[365]$_SDFFE_PN0P_  (.CLK(clknet_leaf_8_clk_p2c),
    .RESET_B(net1773),
    .D(_00997_),
    .Q_N(_05970_),
    .Q(\shift_storage.storage[365] ));
 sg13g2_dfrbp_1 \shift_storage.storage[366]$_SDFFE_PN0P_  (.CLK(clknet_leaf_8_clk_p2c),
    .RESET_B(net1774),
    .D(_00998_),
    .Q_N(_05969_),
    .Q(\shift_storage.storage[366] ));
 sg13g2_dfrbp_1 \shift_storage.storage[367]$_SDFFE_PN0P_  (.CLK(clknet_leaf_7_clk_p2c),
    .RESET_B(net1775),
    .D(_00999_),
    .Q_N(_05968_),
    .Q(\shift_storage.storage[367] ));
 sg13g2_dfrbp_1 \shift_storage.storage[368]$_SDFFE_PN0P_  (.CLK(clknet_leaf_8_clk_p2c),
    .RESET_B(net1776),
    .D(_01000_),
    .Q_N(_05967_),
    .Q(\shift_storage.storage[368] ));
 sg13g2_dfrbp_1 \shift_storage.storage[369]$_SDFFE_PN0P_  (.CLK(clknet_leaf_8_clk_p2c),
    .RESET_B(net1777),
    .D(_01001_),
    .Q_N(_05966_),
    .Q(\shift_storage.storage[369] ));
 sg13g2_dfrbp_1 \shift_storage.storage[36]$_SDFFE_PN0P_  (.CLK(clknet_leaf_96_clk_p2c),
    .RESET_B(net1778),
    .D(_01002_),
    .Q_N(_05965_),
    .Q(\shift_storage.storage[36] ));
 sg13g2_dfrbp_1 \shift_storage.storage[370]$_SDFFE_PN0P_  (.CLK(clknet_leaf_11_clk_p2c),
    .RESET_B(net1779),
    .D(_01003_),
    .Q_N(_05964_),
    .Q(\shift_storage.storage[370] ));
 sg13g2_dfrbp_1 \shift_storage.storage[371]$_SDFFE_PN0P_  (.CLK(clknet_leaf_11_clk_p2c),
    .RESET_B(net1780),
    .D(_01004_),
    .Q_N(_05963_),
    .Q(\shift_storage.storage[371] ));
 sg13g2_dfrbp_1 \shift_storage.storage[372]$_SDFFE_PN0P_  (.CLK(clknet_leaf_11_clk_p2c),
    .RESET_B(net1781),
    .D(_01005_),
    .Q_N(_05962_),
    .Q(\shift_storage.storage[372] ));
 sg13g2_dfrbp_1 \shift_storage.storage[373]$_SDFFE_PN0P_  (.CLK(clknet_leaf_11_clk_p2c),
    .RESET_B(net1782),
    .D(_01006_),
    .Q_N(_05961_),
    .Q(\shift_storage.storage[373] ));
 sg13g2_dfrbp_1 \shift_storage.storage[374]$_SDFFE_PN0P_  (.CLK(clknet_leaf_12_clk_p2c),
    .RESET_B(net1783),
    .D(_01007_),
    .Q_N(_05960_),
    .Q(\shift_storage.storage[374] ));
 sg13g2_dfrbp_1 \shift_storage.storage[375]$_SDFFE_PN0P_  (.CLK(clknet_leaf_12_clk_p2c),
    .RESET_B(net1784),
    .D(_01008_),
    .Q_N(_05959_),
    .Q(\shift_storage.storage[375] ));
 sg13g2_dfrbp_1 \shift_storage.storage[376]$_SDFFE_PN0P_  (.CLK(clknet_leaf_12_clk_p2c),
    .RESET_B(net1785),
    .D(_01009_),
    .Q_N(_05958_),
    .Q(\shift_storage.storage[376] ));
 sg13g2_dfrbp_1 \shift_storage.storage[377]$_SDFFE_PN0P_  (.CLK(clknet_leaf_12_clk_p2c),
    .RESET_B(net1786),
    .D(_01010_),
    .Q_N(_05957_),
    .Q(\shift_storage.storage[377] ));
 sg13g2_dfrbp_1 \shift_storage.storage[378]$_SDFFE_PN0P_  (.CLK(clknet_leaf_23_clk_p2c),
    .RESET_B(net1787),
    .D(_01011_),
    .Q_N(_05956_),
    .Q(\shift_storage.storage[378] ));
 sg13g2_dfrbp_1 \shift_storage.storage[379]$_SDFFE_PN0P_  (.CLK(clknet_leaf_22_clk_p2c),
    .RESET_B(net1788),
    .D(_01012_),
    .Q_N(_05955_),
    .Q(\shift_storage.storage[379] ));
 sg13g2_dfrbp_1 \shift_storage.storage[37]$_SDFFE_PN0P_  (.CLK(clknet_leaf_97_clk_p2c),
    .RESET_B(net1789),
    .D(_01013_),
    .Q_N(_05954_),
    .Q(\shift_storage.storage[37] ));
 sg13g2_dfrbp_1 \shift_storage.storage[380]$_SDFFE_PN0P_  (.CLK(clknet_leaf_23_clk_p2c),
    .RESET_B(net1790),
    .D(_01014_),
    .Q_N(_05953_),
    .Q(\shift_storage.storage[380] ));
 sg13g2_dfrbp_1 \shift_storage.storage[381]$_SDFFE_PN0P_  (.CLK(clknet_leaf_22_clk_p2c),
    .RESET_B(net1791),
    .D(_01015_),
    .Q_N(_05952_),
    .Q(\shift_storage.storage[381] ));
 sg13g2_dfrbp_1 \shift_storage.storage[382]$_SDFFE_PN0P_  (.CLK(clknet_leaf_22_clk_p2c),
    .RESET_B(net1792),
    .D(_01016_),
    .Q_N(_05951_),
    .Q(\shift_storage.storage[382] ));
 sg13g2_dfrbp_1 \shift_storage.storage[383]$_SDFFE_PN0P_  (.CLK(clknet_leaf_22_clk_p2c),
    .RESET_B(net1793),
    .D(_01017_),
    .Q_N(_05950_),
    .Q(\shift_storage.storage[383] ));
 sg13g2_dfrbp_1 \shift_storage.storage[384]$_SDFFE_PN0P_  (.CLK(clknet_leaf_22_clk_p2c),
    .RESET_B(net1794),
    .D(_01018_),
    .Q_N(_05949_),
    .Q(\shift_storage.storage[384] ));
 sg13g2_dfrbp_1 \shift_storage.storage[385]$_SDFFE_PN0P_  (.CLK(clknet_leaf_18_clk_p2c),
    .RESET_B(net1795),
    .D(_01019_),
    .Q_N(_05948_),
    .Q(\shift_storage.storage[385] ));
 sg13g2_dfrbp_1 \shift_storage.storage[386]$_SDFFE_PN0P_  (.CLK(clknet_leaf_21_clk_p2c),
    .RESET_B(net1796),
    .D(_01020_),
    .Q_N(_05947_),
    .Q(\shift_storage.storage[386] ));
 sg13g2_dfrbp_1 \shift_storage.storage[387]$_SDFFE_PN0P_  (.CLK(clknet_leaf_21_clk_p2c),
    .RESET_B(net1797),
    .D(_01021_),
    .Q_N(_05946_),
    .Q(\shift_storage.storage[387] ));
 sg13g2_dfrbp_1 \shift_storage.storage[388]$_SDFFE_PN0P_  (.CLK(clknet_leaf_20_clk_p2c),
    .RESET_B(net1798),
    .D(_01022_),
    .Q_N(_05945_),
    .Q(\shift_storage.storage[388] ));
 sg13g2_dfrbp_1 \shift_storage.storage[389]$_SDFFE_PN0P_  (.CLK(clknet_leaf_21_clk_p2c),
    .RESET_B(net1799),
    .D(_01023_),
    .Q_N(_05944_),
    .Q(\shift_storage.storage[389] ));
 sg13g2_dfrbp_1 \shift_storage.storage[38]$_SDFFE_PN0P_  (.CLK(clknet_leaf_97_clk_p2c),
    .RESET_B(net1800),
    .D(_01024_),
    .Q_N(_05943_),
    .Q(\shift_storage.storage[38] ));
 sg13g2_dfrbp_1 \shift_storage.storage[390]$_SDFFE_PN0P_  (.CLK(clknet_leaf_21_clk_p2c),
    .RESET_B(net1801),
    .D(_01025_),
    .Q_N(_05942_),
    .Q(\shift_storage.storage[390] ));
 sg13g2_dfrbp_1 \shift_storage.storage[391]$_SDFFE_PN0P_  (.CLK(clknet_leaf_21_clk_p2c),
    .RESET_B(net1802),
    .D(_01026_),
    .Q_N(_05941_),
    .Q(\shift_storage.storage[391] ));
 sg13g2_dfrbp_1 \shift_storage.storage[392]$_SDFFE_PN0P_  (.CLK(clknet_leaf_21_clk_p2c),
    .RESET_B(net1803),
    .D(_01027_),
    .Q_N(_05940_),
    .Q(\shift_storage.storage[392] ));
 sg13g2_dfrbp_1 \shift_storage.storage[393]$_SDFFE_PN0P_  (.CLK(clknet_leaf_21_clk_p2c),
    .RESET_B(net1804),
    .D(_01028_),
    .Q_N(_05939_),
    .Q(\shift_storage.storage[393] ));
 sg13g2_dfrbp_1 \shift_storage.storage[394]$_SDFFE_PN0P_  (.CLK(clknet_leaf_30_clk_p2c),
    .RESET_B(net1805),
    .D(_01029_),
    .Q_N(_05938_),
    .Q(\shift_storage.storage[394] ));
 sg13g2_dfrbp_1 \shift_storage.storage[395]$_SDFFE_PN0P_  (.CLK(clknet_leaf_29_clk_p2c),
    .RESET_B(net1806),
    .D(_01030_),
    .Q_N(_05937_),
    .Q(\shift_storage.storage[395] ));
 sg13g2_dfrbp_1 \shift_storage.storage[396]$_SDFFE_PN0P_  (.CLK(clknet_leaf_27_clk_p2c),
    .RESET_B(net1807),
    .D(_01031_),
    .Q_N(_05936_),
    .Q(\shift_storage.storage[396] ));
 sg13g2_dfrbp_1 \shift_storage.storage[397]$_SDFFE_PN0P_  (.CLK(clknet_leaf_27_clk_p2c),
    .RESET_B(net1808),
    .D(_01032_),
    .Q_N(_05935_),
    .Q(\shift_storage.storage[397] ));
 sg13g2_dfrbp_1 \shift_storage.storage[398]$_SDFFE_PN0P_  (.CLK(clknet_leaf_27_clk_p2c),
    .RESET_B(net1809),
    .D(_01033_),
    .Q_N(_05934_),
    .Q(\shift_storage.storage[398] ));
 sg13g2_dfrbp_1 \shift_storage.storage[399]$_SDFFE_PN0P_  (.CLK(clknet_leaf_27_clk_p2c),
    .RESET_B(net1810),
    .D(_01034_),
    .Q_N(_05933_),
    .Q(\shift_storage.storage[399] ));
 sg13g2_dfrbp_1 \shift_storage.storage[39]$_SDFFE_PN0P_  (.CLK(clknet_leaf_97_clk_p2c),
    .RESET_B(net1811),
    .D(_01035_),
    .Q_N(_05932_),
    .Q(\shift_storage.storage[39] ));
 sg13g2_dfrbp_1 \shift_storage.storage[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_76_clk_p2c),
    .RESET_B(net1812),
    .D(_01036_),
    .Q_N(_05931_),
    .Q(\shift_storage.storage[3] ));
 sg13g2_dfrbp_1 \shift_storage.storage[400]$_SDFFE_PN0P_  (.CLK(clknet_leaf_27_clk_p2c),
    .RESET_B(net1813),
    .D(_01037_),
    .Q_N(_05930_),
    .Q(\shift_storage.storage[400] ));
 sg13g2_dfrbp_1 \shift_storage.storage[401]$_SDFFE_PN0P_  (.CLK(clknet_leaf_29_clk_p2c),
    .RESET_B(net1814),
    .D(_01038_),
    .Q_N(_05929_),
    .Q(\shift_storage.storage[401] ));
 sg13g2_dfrbp_1 \shift_storage.storage[402]$_SDFFE_PN0P_  (.CLK(clknet_leaf_29_clk_p2c),
    .RESET_B(net1815),
    .D(_01039_),
    .Q_N(_05928_),
    .Q(\shift_storage.storage[402] ));
 sg13g2_dfrbp_1 \shift_storage.storage[403]$_SDFFE_PN0P_  (.CLK(clknet_leaf_28_clk_p2c),
    .RESET_B(net1816),
    .D(_01040_),
    .Q_N(_05927_),
    .Q(\shift_storage.storage[403] ));
 sg13g2_dfrbp_1 \shift_storage.storage[404]$_SDFFE_PN0P_  (.CLK(clknet_leaf_28_clk_p2c),
    .RESET_B(net1817),
    .D(_01041_),
    .Q_N(_05926_),
    .Q(\shift_storage.storage[404] ));
 sg13g2_dfrbp_1 \shift_storage.storage[405]$_SDFFE_PN0P_  (.CLK(clknet_leaf_28_clk_p2c),
    .RESET_B(net1818),
    .D(_01042_),
    .Q_N(_05925_),
    .Q(\shift_storage.storage[405] ));
 sg13g2_dfrbp_1 \shift_storage.storage[406]$_SDFFE_PN0P_  (.CLK(clknet_leaf_33_clk_p2c),
    .RESET_B(net1819),
    .D(_01043_),
    .Q_N(_05924_),
    .Q(\shift_storage.storage[406] ));
 sg13g2_dfrbp_1 \shift_storage.storage[407]$_SDFFE_PN0P_  (.CLK(clknet_leaf_33_clk_p2c),
    .RESET_B(net1820),
    .D(_01044_),
    .Q_N(_05923_),
    .Q(\shift_storage.storage[407] ));
 sg13g2_dfrbp_1 \shift_storage.storage[408]$_SDFFE_PN0P_  (.CLK(clknet_leaf_246_clk_p2c),
    .RESET_B(net1821),
    .D(_01045_),
    .Q_N(_05922_),
    .Q(\shift_storage.storage[408] ));
 sg13g2_dfrbp_1 \shift_storage.storage[409]$_SDFFE_PN0P_  (.CLK(clknet_leaf_246_clk_p2c),
    .RESET_B(net1822),
    .D(_01046_),
    .Q_N(_05921_),
    .Q(\shift_storage.storage[409] ));
 sg13g2_dfrbp_1 \shift_storage.storage[40]$_SDFFE_PN0P_  (.CLK(clknet_leaf_46_clk_p2c),
    .RESET_B(net1823),
    .D(_01047_),
    .Q_N(_05920_),
    .Q(\shift_storage.storage[40] ));
 sg13g2_dfrbp_1 \shift_storage.storage[410]$_SDFFE_PN0P_  (.CLK(clknet_leaf_33_clk_p2c),
    .RESET_B(net1824),
    .D(_01048_),
    .Q_N(_05919_),
    .Q(\shift_storage.storage[410] ));
 sg13g2_dfrbp_1 \shift_storage.storage[411]$_SDFFE_PN0P_  (.CLK(clknet_leaf_33_clk_p2c),
    .RESET_B(net1825),
    .D(_01049_),
    .Q_N(_05918_),
    .Q(\shift_storage.storage[411] ));
 sg13g2_dfrbp_1 \shift_storage.storage[412]$_SDFFE_PN0P_  (.CLK(clknet_leaf_246_clk_p2c),
    .RESET_B(net1826),
    .D(_01050_),
    .Q_N(_05917_),
    .Q(\shift_storage.storage[412] ));
 sg13g2_dfrbp_1 \shift_storage.storage[413]$_SDFFE_PN0P_  (.CLK(clknet_leaf_246_clk_p2c),
    .RESET_B(net1827),
    .D(_01051_),
    .Q_N(_05916_),
    .Q(\shift_storage.storage[413] ));
 sg13g2_dfrbp_1 \shift_storage.storage[414]$_SDFFE_PN0P_  (.CLK(clknet_leaf_245_clk_p2c),
    .RESET_B(net1828),
    .D(_01052_),
    .Q_N(_05915_),
    .Q(\shift_storage.storage[414] ));
 sg13g2_dfrbp_1 \shift_storage.storage[415]$_SDFFE_PN0P_  (.CLK(clknet_leaf_245_clk_p2c),
    .RESET_B(net1829),
    .D(_01053_),
    .Q_N(_05914_),
    .Q(\shift_storage.storage[415] ));
 sg13g2_dfrbp_1 \shift_storage.storage[416]$_SDFFE_PN0P_  (.CLK(clknet_leaf_245_clk_p2c),
    .RESET_B(net1830),
    .D(_01054_),
    .Q_N(_05913_),
    .Q(\shift_storage.storage[416] ));
 sg13g2_dfrbp_1 \shift_storage.storage[417]$_SDFFE_PN0P_  (.CLK(clknet_leaf_245_clk_p2c),
    .RESET_B(net1831),
    .D(_01055_),
    .Q_N(_05912_),
    .Q(\shift_storage.storage[417] ));
 sg13g2_dfrbp_1 \shift_storage.storage[418]$_SDFFE_PN0P_  (.CLK(clknet_leaf_245_clk_p2c),
    .RESET_B(net1832),
    .D(_01056_),
    .Q_N(_05911_),
    .Q(\shift_storage.storage[418] ));
 sg13g2_dfrbp_1 \shift_storage.storage[419]$_SDFFE_PN0P_  (.CLK(clknet_leaf_246_clk_p2c),
    .RESET_B(net1833),
    .D(_01057_),
    .Q_N(_05910_),
    .Q(\shift_storage.storage[419] ));
 sg13g2_dfrbp_1 \shift_storage.storage[41]$_SDFFE_PN0P_  (.CLK(clknet_leaf_46_clk_p2c),
    .RESET_B(net1834),
    .D(_01058_),
    .Q_N(_05909_),
    .Q(\shift_storage.storage[41] ));
 sg13g2_dfrbp_1 \shift_storage.storage[420]$_SDFFE_PN0P_  (.CLK(clknet_leaf_247_clk_p2c),
    .RESET_B(net1835),
    .D(_01059_),
    .Q_N(_05908_),
    .Q(\shift_storage.storage[420] ));
 sg13g2_dfrbp_1 \shift_storage.storage[421]$_SDFFE_PN0P_  (.CLK(clknet_leaf_247_clk_p2c),
    .RESET_B(net1836),
    .D(_01060_),
    .Q_N(_05907_),
    .Q(\shift_storage.storage[421] ));
 sg13g2_dfrbp_1 \shift_storage.storage[422]$_SDFFE_PN0P_  (.CLK(clknet_leaf_247_clk_p2c),
    .RESET_B(net1837),
    .D(_01061_),
    .Q_N(_05906_),
    .Q(\shift_storage.storage[422] ));
 sg13g2_dfrbp_1 \shift_storage.storage[423]$_SDFFE_PN0P_  (.CLK(clknet_leaf_251_clk_p2c),
    .RESET_B(net1838),
    .D(_01062_),
    .Q_N(_05905_),
    .Q(\shift_storage.storage[423] ));
 sg13g2_dfrbp_1 \shift_storage.storage[424]$_SDFFE_PN0P_  (.CLK(clknet_leaf_252_clk_p2c),
    .RESET_B(net1839),
    .D(_01063_),
    .Q_N(_05904_),
    .Q(\shift_storage.storage[424] ));
 sg13g2_dfrbp_1 \shift_storage.storage[425]$_SDFFE_PN0P_  (.CLK(clknet_leaf_252_clk_p2c),
    .RESET_B(net1840),
    .D(_01064_),
    .Q_N(_05903_),
    .Q(\shift_storage.storage[425] ));
 sg13g2_dfrbp_1 \shift_storage.storage[426]$_SDFFE_PN0P_  (.CLK(clknet_leaf_251_clk_p2c),
    .RESET_B(net1841),
    .D(_01065_),
    .Q_N(_05902_),
    .Q(\shift_storage.storage[426] ));
 sg13g2_dfrbp_1 \shift_storage.storage[427]$_SDFFE_PN0P_  (.CLK(clknet_leaf_252_clk_p2c),
    .RESET_B(net1842),
    .D(_01066_),
    .Q_N(_05901_),
    .Q(\shift_storage.storage[427] ));
 sg13g2_dfrbp_1 \shift_storage.storage[428]$_SDFFE_PN0P_  (.CLK(clknet_leaf_252_clk_p2c),
    .RESET_B(net1843),
    .D(_01067_),
    .Q_N(_05900_),
    .Q(\shift_storage.storage[428] ));
 sg13g2_dfrbp_1 \shift_storage.storage[429]$_SDFFE_PN0P_  (.CLK(clknet_leaf_252_clk_p2c),
    .RESET_B(net1844),
    .D(_01068_),
    .Q_N(_05899_),
    .Q(\shift_storage.storage[429] ));
 sg13g2_dfrbp_1 \shift_storage.storage[42]$_SDFFE_PN0P_  (.CLK(clknet_leaf_45_clk_p2c),
    .RESET_B(net1845),
    .D(_01069_),
    .Q_N(_05898_),
    .Q(\shift_storage.storage[42] ));
 sg13g2_dfrbp_1 \shift_storage.storage[430]$_SDFFE_PN0P_  (.CLK(clknet_leaf_253_clk_p2c),
    .RESET_B(net1846),
    .D(_01070_),
    .Q_N(_05897_),
    .Q(\shift_storage.storage[430] ));
 sg13g2_dfrbp_1 \shift_storage.storage[431]$_SDFFE_PN0P_  (.CLK(clknet_leaf_254_clk_p2c),
    .RESET_B(net1847),
    .D(_01071_),
    .Q_N(_05896_),
    .Q(\shift_storage.storage[431] ));
 sg13g2_dfrbp_1 \shift_storage.storage[432]$_SDFFE_PN0P_  (.CLK(clknet_leaf_252_clk_p2c),
    .RESET_B(net1848),
    .D(_01072_),
    .Q_N(_05895_),
    .Q(\shift_storage.storage[432] ));
 sg13g2_dfrbp_1 \shift_storage.storage[433]$_SDFFE_PN0P_  (.CLK(clknet_leaf_28_clk_p2c),
    .RESET_B(net1849),
    .D(_01073_),
    .Q_N(_05894_),
    .Q(\shift_storage.storage[433] ));
 sg13g2_dfrbp_1 \shift_storage.storage[434]$_SDFFE_PN0P_  (.CLK(clknet_leaf_26_clk_p2c),
    .RESET_B(net1850),
    .D(_01074_),
    .Q_N(_05893_),
    .Q(\shift_storage.storage[434] ));
 sg13g2_dfrbp_1 \shift_storage.storage[435]$_SDFFE_PN0P_  (.CLK(clknet_leaf_26_clk_p2c),
    .RESET_B(net1851),
    .D(_01075_),
    .Q_N(_05892_),
    .Q(\shift_storage.storage[435] ));
 sg13g2_dfrbp_1 \shift_storage.storage[436]$_SDFFE_PN0P_  (.CLK(clknet_leaf_26_clk_p2c),
    .RESET_B(net1852),
    .D(_01076_),
    .Q_N(_05891_),
    .Q(\shift_storage.storage[436] ));
 sg13g2_dfrbp_1 \shift_storage.storage[437]$_SDFFE_PN0P_  (.CLK(clknet_leaf_26_clk_p2c),
    .RESET_B(net1853),
    .D(_01077_),
    .Q_N(_05890_),
    .Q(\shift_storage.storage[437] ));
 sg13g2_dfrbp_1 \shift_storage.storage[438]$_SDFFE_PN0P_  (.CLK(clknet_leaf_26_clk_p2c),
    .RESET_B(net1854),
    .D(_01078_),
    .Q_N(_05889_),
    .Q(\shift_storage.storage[438] ));
 sg13g2_dfrbp_1 \shift_storage.storage[439]$_SDFFE_PN0P_  (.CLK(clknet_leaf_25_clk_p2c),
    .RESET_B(net1855),
    .D(_01079_),
    .Q_N(_05888_),
    .Q(\shift_storage.storage[439] ));
 sg13g2_dfrbp_1 \shift_storage.storage[43]$_SDFFE_PN0P_  (.CLK(clknet_leaf_46_clk_p2c),
    .RESET_B(net1856),
    .D(_01080_),
    .Q_N(_05887_),
    .Q(\shift_storage.storage[43] ));
 sg13g2_dfrbp_1 \shift_storage.storage[440]$_SDFFE_PN0P_  (.CLK(clknet_leaf_24_clk_p2c),
    .RESET_B(net1857),
    .D(_01081_),
    .Q_N(_05886_),
    .Q(\shift_storage.storage[440] ));
 sg13g2_dfrbp_1 \shift_storage.storage[441]$_SDFFE_PN0P_  (.CLK(clknet_leaf_24_clk_p2c),
    .RESET_B(net1858),
    .D(_01082_),
    .Q_N(_05885_),
    .Q(\shift_storage.storage[441] ));
 sg13g2_dfrbp_1 \shift_storage.storage[442]$_SDFFE_PN0P_  (.CLK(clknet_leaf_24_clk_p2c),
    .RESET_B(net1859),
    .D(_01083_),
    .Q_N(_05884_),
    .Q(\shift_storage.storage[442] ));
 sg13g2_dfrbp_1 \shift_storage.storage[443]$_SDFFE_PN0P_  (.CLK(clknet_leaf_24_clk_p2c),
    .RESET_B(net1860),
    .D(_01084_),
    .Q_N(_05883_),
    .Q(\shift_storage.storage[443] ));
 sg13g2_dfrbp_1 \shift_storage.storage[444]$_SDFFE_PN0P_  (.CLK(clknet_leaf_24_clk_p2c),
    .RESET_B(net1861),
    .D(_01085_),
    .Q_N(_05882_),
    .Q(\shift_storage.storage[444] ));
 sg13g2_dfrbp_1 \shift_storage.storage[445]$_SDFFE_PN0P_  (.CLK(clknet_leaf_23_clk_p2c),
    .RESET_B(net1862),
    .D(_01086_),
    .Q_N(_05881_),
    .Q(\shift_storage.storage[445] ));
 sg13g2_dfrbp_1 \shift_storage.storage[446]$_SDFFE_PN0P_  (.CLK(clknet_leaf_23_clk_p2c),
    .RESET_B(net1863),
    .D(_01087_),
    .Q_N(_05880_),
    .Q(\shift_storage.storage[446] ));
 sg13g2_dfrbp_1 \shift_storage.storage[447]$_SDFFE_PN0P_  (.CLK(clknet_leaf_23_clk_p2c),
    .RESET_B(net1864),
    .D(_01088_),
    .Q_N(_05879_),
    .Q(\shift_storage.storage[447] ));
 sg13g2_dfrbp_1 \shift_storage.storage[448]$_SDFFE_PN0P_  (.CLK(clknet_leaf_23_clk_p2c),
    .RESET_B(net1865),
    .D(_01089_),
    .Q_N(_05878_),
    .Q(\shift_storage.storage[448] ));
 sg13g2_dfrbp_1 \shift_storage.storage[449]$_SDFFE_PN0P_  (.CLK(clknet_leaf_7_clk_p2c),
    .RESET_B(net1866),
    .D(_01090_),
    .Q_N(_05877_),
    .Q(\shift_storage.storage[449] ));
 sg13g2_dfrbp_1 \shift_storage.storage[44]$_SDFFE_PN0P_  (.CLK(clknet_leaf_44_clk_p2c),
    .RESET_B(net1867),
    .D(_01091_),
    .Q_N(_05876_),
    .Q(\shift_storage.storage[44] ));
 sg13g2_dfrbp_1 \shift_storage.storage[450]$_SDFFE_PN0P_  (.CLK(clknet_leaf_7_clk_p2c),
    .RESET_B(net1868),
    .D(_01092_),
    .Q_N(_05875_),
    .Q(\shift_storage.storage[450] ));
 sg13g2_dfrbp_1 \shift_storage.storage[451]$_SDFFE_PN0P_  (.CLK(clknet_leaf_7_clk_p2c),
    .RESET_B(net1869),
    .D(_01093_),
    .Q_N(_05874_),
    .Q(\shift_storage.storage[451] ));
 sg13g2_dfrbp_1 \shift_storage.storage[452]$_SDFFE_PN0P_  (.CLK(clknet_leaf_7_clk_p2c),
    .RESET_B(net1870),
    .D(_01094_),
    .Q_N(_05873_),
    .Q(\shift_storage.storage[452] ));
 sg13g2_dfrbp_1 \shift_storage.storage[453]$_SDFFE_PN0P_  (.CLK(clknet_leaf_7_clk_p2c),
    .RESET_B(net1871),
    .D(_01095_),
    .Q_N(_05872_),
    .Q(\shift_storage.storage[453] ));
 sg13g2_dfrbp_1 \shift_storage.storage[454]$_SDFFE_PN0P_  (.CLK(clknet_leaf_6_clk_p2c),
    .RESET_B(net1872),
    .D(_01096_),
    .Q_N(_05871_),
    .Q(\shift_storage.storage[454] ));
 sg13g2_dfrbp_1 \shift_storage.storage[455]$_SDFFE_PN0P_  (.CLK(clknet_leaf_5_clk_p2c),
    .RESET_B(net1873),
    .D(_01097_),
    .Q_N(_05870_),
    .Q(\shift_storage.storage[455] ));
 sg13g2_dfrbp_1 \shift_storage.storage[456]$_SDFFE_PN0P_  (.CLK(clknet_leaf_5_clk_p2c),
    .RESET_B(net1874),
    .D(_01098_),
    .Q_N(_05869_),
    .Q(\shift_storage.storage[456] ));
 sg13g2_dfrbp_1 \shift_storage.storage[457]$_SDFFE_PN0P_  (.CLK(clknet_leaf_5_clk_p2c),
    .RESET_B(net1875),
    .D(_01099_),
    .Q_N(_05868_),
    .Q(\shift_storage.storage[457] ));
 sg13g2_dfrbp_1 \shift_storage.storage[458]$_SDFFE_PN0P_  (.CLK(clknet_leaf_5_clk_p2c),
    .RESET_B(net1876),
    .D(_01100_),
    .Q_N(_05867_),
    .Q(\shift_storage.storage[458] ));
 sg13g2_dfrbp_1 \shift_storage.storage[459]$_SDFFE_PN0P_  (.CLK(clknet_leaf_5_clk_p2c),
    .RESET_B(net1877),
    .D(_01101_),
    .Q_N(_05866_),
    .Q(\shift_storage.storage[459] ));
 sg13g2_dfrbp_1 \shift_storage.storage[45]$_SDFFE_PN0P_  (.CLK(clknet_leaf_44_clk_p2c),
    .RESET_B(net1878),
    .D(_01102_),
    .Q_N(_05865_),
    .Q(\shift_storage.storage[45] ));
 sg13g2_dfrbp_1 \shift_storage.storage[460]$_SDFFE_PN0P_  (.CLK(clknet_leaf_25_clk_p2c),
    .RESET_B(net1879),
    .D(_01103_),
    .Q_N(_05864_),
    .Q(\shift_storage.storage[460] ));
 sg13g2_dfrbp_1 \shift_storage.storage[461]$_SDFFE_PN0P_  (.CLK(clknet_leaf_25_clk_p2c),
    .RESET_B(net1880),
    .D(_01104_),
    .Q_N(_05863_),
    .Q(\shift_storage.storage[461] ));
 sg13g2_dfrbp_1 \shift_storage.storage[462]$_SDFFE_PN0P_  (.CLK(clknet_leaf_25_clk_p2c),
    .RESET_B(net1881),
    .D(_01105_),
    .Q_N(_05862_),
    .Q(\shift_storage.storage[462] ));
 sg13g2_dfrbp_1 \shift_storage.storage[463]$_SDFFE_PN0P_  (.CLK(clknet_leaf_254_clk_p2c),
    .RESET_B(net1882),
    .D(_01106_),
    .Q_N(_05861_),
    .Q(\shift_storage.storage[463] ));
 sg13g2_dfrbp_1 \shift_storage.storage[464]$_SDFFE_PN0P_  (.CLK(clknet_leaf_254_clk_p2c),
    .RESET_B(net1883),
    .D(_01107_),
    .Q_N(_05860_),
    .Q(\shift_storage.storage[464] ));
 sg13g2_dfrbp_1 \shift_storage.storage[465]$_SDFFE_PN0P_  (.CLK(clknet_leaf_254_clk_p2c),
    .RESET_B(net1884),
    .D(_01108_),
    .Q_N(_05859_),
    .Q(\shift_storage.storage[465] ));
 sg13g2_dfrbp_1 \shift_storage.storage[466]$_SDFFE_PN0P_  (.CLK(clknet_leaf_254_clk_p2c),
    .RESET_B(net1885),
    .D(_01109_),
    .Q_N(_05858_),
    .Q(\shift_storage.storage[466] ));
 sg13g2_dfrbp_1 \shift_storage.storage[467]$_SDFFE_PN0P_  (.CLK(clknet_leaf_253_clk_p2c),
    .RESET_B(net1886),
    .D(_01110_),
    .Q_N(_05857_),
    .Q(\shift_storage.storage[467] ));
 sg13g2_dfrbp_1 \shift_storage.storage[468]$_SDFFE_PN0P_  (.CLK(clknet_leaf_253_clk_p2c),
    .RESET_B(net1887),
    .D(_01111_),
    .Q_N(_05856_),
    .Q(\shift_storage.storage[468] ));
 sg13g2_dfrbp_1 \shift_storage.storage[469]$_SDFFE_PN0P_  (.CLK(clknet_leaf_253_clk_p2c),
    .RESET_B(net1888),
    .D(_01112_),
    .Q_N(_05855_),
    .Q(\shift_storage.storage[469] ));
 sg13g2_dfrbp_1 \shift_storage.storage[46]$_SDFFE_PN0P_  (.CLK(clknet_leaf_44_clk_p2c),
    .RESET_B(net1889),
    .D(_01113_),
    .Q_N(_05854_),
    .Q(\shift_storage.storage[46] ));
 sg13g2_dfrbp_1 \shift_storage.storage[470]$_SDFFE_PN0P_  (.CLK(clknet_leaf_253_clk_p2c),
    .RESET_B(net1890),
    .D(_01114_),
    .Q_N(_05853_),
    .Q(\shift_storage.storage[470] ));
 sg13g2_dfrbp_1 \shift_storage.storage[471]$_SDFFE_PN0P_  (.CLK(clknet_leaf_255_clk_p2c),
    .RESET_B(net1891),
    .D(_01115_),
    .Q_N(_05852_),
    .Q(\shift_storage.storage[471] ));
 sg13g2_dfrbp_1 \shift_storage.storage[472]$_SDFFE_PN0P_  (.CLK(clknet_leaf_259_clk_p2c),
    .RESET_B(net1892),
    .D(_01116_),
    .Q_N(_05851_),
    .Q(\shift_storage.storage[472] ));
 sg13g2_dfrbp_1 \shift_storage.storage[473]$_SDFFE_PN0P_  (.CLK(clknet_leaf_250_clk_p2c),
    .RESET_B(net1893),
    .D(_01117_),
    .Q_N(_05850_),
    .Q(\shift_storage.storage[473] ));
 sg13g2_dfrbp_1 \shift_storage.storage[474]$_SDFFE_PN0P_  (.CLK(clknet_leaf_250_clk_p2c),
    .RESET_B(net1894),
    .D(_01118_),
    .Q_N(_05849_),
    .Q(\shift_storage.storage[474] ));
 sg13g2_dfrbp_1 \shift_storage.storage[475]$_SDFFE_PN0P_  (.CLK(clknet_leaf_250_clk_p2c),
    .RESET_B(net1895),
    .D(_01119_),
    .Q_N(_05848_),
    .Q(\shift_storage.storage[475] ));
 sg13g2_dfrbp_1 \shift_storage.storage[476]$_SDFFE_PN0P_  (.CLK(clknet_leaf_250_clk_p2c),
    .RESET_B(net1896),
    .D(_01120_),
    .Q_N(_05847_),
    .Q(\shift_storage.storage[476] ));
 sg13g2_dfrbp_1 \shift_storage.storage[477]$_SDFFE_PN0P_  (.CLK(clknet_leaf_251_clk_p2c),
    .RESET_B(net1897),
    .D(_01121_),
    .Q_N(_05846_),
    .Q(\shift_storage.storage[477] ));
 sg13g2_dfrbp_1 \shift_storage.storage[478]$_SDFFE_PN0P_  (.CLK(clknet_leaf_251_clk_p2c),
    .RESET_B(net1898),
    .D(_01122_),
    .Q_N(_05845_),
    .Q(\shift_storage.storage[478] ));
 sg13g2_dfrbp_1 \shift_storage.storage[479]$_SDFFE_PN0P_  (.CLK(clknet_leaf_251_clk_p2c),
    .RESET_B(net1899),
    .D(_01123_),
    .Q_N(_05844_),
    .Q(\shift_storage.storage[479] ));
 sg13g2_dfrbp_1 \shift_storage.storage[47]$_SDFFE_PN0P_  (.CLK(clknet_leaf_45_clk_p2c),
    .RESET_B(net1900),
    .D(_01124_),
    .Q_N(_05843_),
    .Q(\shift_storage.storage[47] ));
 sg13g2_dfrbp_1 \shift_storage.storage[480]$_SDFFE_PN0P_  (.CLK(clknet_leaf_251_clk_p2c),
    .RESET_B(net1901),
    .D(_01125_),
    .Q_N(_05842_),
    .Q(\shift_storage.storage[480] ));
 sg13g2_dfrbp_1 \shift_storage.storage[481]$_SDFFE_PN0P_  (.CLK(clknet_leaf_248_clk_p2c),
    .RESET_B(net1902),
    .D(_01126_),
    .Q_N(_05841_),
    .Q(\shift_storage.storage[481] ));
 sg13g2_dfrbp_1 \shift_storage.storage[482]$_SDFFE_PN0P_  (.CLK(clknet_leaf_247_clk_p2c),
    .RESET_B(net1903),
    .D(_01127_),
    .Q_N(_05840_),
    .Q(\shift_storage.storage[482] ));
 sg13g2_dfrbp_1 \shift_storage.storage[483]$_SDFFE_PN0P_  (.CLK(clknet_leaf_247_clk_p2c),
    .RESET_B(net1904),
    .D(_01128_),
    .Q_N(_05839_),
    .Q(\shift_storage.storage[483] ));
 sg13g2_dfrbp_1 \shift_storage.storage[484]$_SDFFE_PN0P_  (.CLK(clknet_leaf_247_clk_p2c),
    .RESET_B(net1905),
    .D(_01129_),
    .Q_N(_05838_),
    .Q(\shift_storage.storage[484] ));
 sg13g2_dfrbp_1 \shift_storage.storage[485]$_SDFFE_PN0P_  (.CLK(clknet_leaf_248_clk_p2c),
    .RESET_B(net1906),
    .D(_01130_),
    .Q_N(_05837_),
    .Q(\shift_storage.storage[485] ));
 sg13g2_dfrbp_1 \shift_storage.storage[486]$_SDFFE_PN0P_  (.CLK(clknet_leaf_248_clk_p2c),
    .RESET_B(net1907),
    .D(_01131_),
    .Q_N(_05836_),
    .Q(\shift_storage.storage[486] ));
 sg13g2_dfrbp_1 \shift_storage.storage[487]$_SDFFE_PN0P_  (.CLK(clknet_leaf_239_clk_p2c),
    .RESET_B(net1908),
    .D(_01132_),
    .Q_N(_05835_),
    .Q(\shift_storage.storage[487] ));
 sg13g2_dfrbp_1 \shift_storage.storage[488]$_SDFFE_PN0P_  (.CLK(clknet_leaf_238_clk_p2c),
    .RESET_B(net1909),
    .D(_01133_),
    .Q_N(_05834_),
    .Q(\shift_storage.storage[488] ));
 sg13g2_dfrbp_1 \shift_storage.storage[489]$_SDFFE_PN0P_  (.CLK(clknet_leaf_248_clk_p2c),
    .RESET_B(net1910),
    .D(_01134_),
    .Q_N(_05833_),
    .Q(\shift_storage.storage[489] ));
 sg13g2_dfrbp_1 \shift_storage.storage[48]$_SDFFE_PN0P_  (.CLK(clknet_leaf_39_clk_p2c),
    .RESET_B(net1911),
    .D(_01135_),
    .Q_N(_05832_),
    .Q(\shift_storage.storage[48] ));
 sg13g2_dfrbp_1 \shift_storage.storage[490]$_SDFFE_PN0P_  (.CLK(clknet_leaf_248_clk_p2c),
    .RESET_B(net1912),
    .D(_01136_),
    .Q_N(_05831_),
    .Q(\shift_storage.storage[490] ));
 sg13g2_dfrbp_1 \shift_storage.storage[491]$_SDFFE_PN0P_  (.CLK(clknet_leaf_249_clk_p2c),
    .RESET_B(net1913),
    .D(_01137_),
    .Q_N(_05830_),
    .Q(\shift_storage.storage[491] ));
 sg13g2_dfrbp_1 \shift_storage.storage[492]$_SDFFE_PN0P_  (.CLK(clknet_leaf_249_clk_p2c),
    .RESET_B(net1914),
    .D(_01138_),
    .Q_N(_05829_),
    .Q(\shift_storage.storage[492] ));
 sg13g2_dfrbp_1 \shift_storage.storage[493]$_SDFFE_PN0P_  (.CLK(clknet_leaf_249_clk_p2c),
    .RESET_B(net1915),
    .D(_01139_),
    .Q_N(_05828_),
    .Q(\shift_storage.storage[493] ));
 sg13g2_dfrbp_1 \shift_storage.storage[494]$_SDFFE_PN0P_  (.CLK(clknet_leaf_249_clk_p2c),
    .RESET_B(net1916),
    .D(_01140_),
    .Q_N(_05827_),
    .Q(\shift_storage.storage[494] ));
 sg13g2_dfrbp_1 \shift_storage.storage[495]$_SDFFE_PN0P_  (.CLK(clknet_leaf_249_clk_p2c),
    .RESET_B(net1917),
    .D(_01141_),
    .Q_N(_05826_),
    .Q(\shift_storage.storage[495] ));
 sg13g2_dfrbp_1 \shift_storage.storage[496]$_SDFFE_PN0P_  (.CLK(clknet_leaf_249_clk_p2c),
    .RESET_B(net1918),
    .D(_01142_),
    .Q_N(_05825_),
    .Q(\shift_storage.storage[496] ));
 sg13g2_dfrbp_1 \shift_storage.storage[497]$_SDFFE_PN0P_  (.CLK(clknet_leaf_250_clk_p2c),
    .RESET_B(net1919),
    .D(_01143_),
    .Q_N(_05824_),
    .Q(\shift_storage.storage[497] ));
 sg13g2_dfrbp_1 \shift_storage.storage[498]$_SDFFE_PN0P_  (.CLK(clknet_leaf_250_clk_p2c),
    .RESET_B(net1920),
    .D(_01144_),
    .Q_N(_05823_),
    .Q(\shift_storage.storage[498] ));
 sg13g2_dfrbp_1 \shift_storage.storage[499]$_SDFFE_PN0P_  (.CLK(clknet_leaf_250_clk_p2c),
    .RESET_B(net1921),
    .D(_01145_),
    .Q_N(_05822_),
    .Q(\shift_storage.storage[499] ));
 sg13g2_dfrbp_1 \shift_storage.storage[49]$_SDFFE_PN0P_  (.CLK(clknet_leaf_39_clk_p2c),
    .RESET_B(net1922),
    .D(_01146_),
    .Q_N(_05821_),
    .Q(\shift_storage.storage[49] ));
 sg13g2_dfrbp_1 \shift_storage.storage[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_75_clk_p2c),
    .RESET_B(net1923),
    .D(_01147_),
    .Q_N(_05820_),
    .Q(\shift_storage.storage[4] ));
 sg13g2_dfrbp_1 \shift_storage.storage[500]$_SDFFE_PN0P_  (.CLK(clknet_leaf_259_clk_p2c),
    .RESET_B(net1924),
    .D(_01148_),
    .Q_N(_05819_),
    .Q(\shift_storage.storage[500] ));
 sg13g2_dfrbp_1 \shift_storage.storage[501]$_SDFFE_PN0P_  (.CLK(clknet_leaf_259_clk_p2c),
    .RESET_B(net1925),
    .D(_01149_),
    .Q_N(_05818_),
    .Q(\shift_storage.storage[501] ));
 sg13g2_dfrbp_1 \shift_storage.storage[502]$_SDFFE_PN0P_  (.CLK(clknet_leaf_258_clk_p2c),
    .RESET_B(net1926),
    .D(_01150_),
    .Q_N(_05817_),
    .Q(\shift_storage.storage[502] ));
 sg13g2_dfrbp_1 \shift_storage.storage[503]$_SDFFE_PN0P_  (.CLK(clknet_leaf_258_clk_p2c),
    .RESET_B(net1927),
    .D(_01151_),
    .Q_N(_05816_),
    .Q(\shift_storage.storage[503] ));
 sg13g2_dfrbp_1 \shift_storage.storage[504]$_SDFFE_PN0P_  (.CLK(clknet_leaf_258_clk_p2c),
    .RESET_B(net1928),
    .D(_01152_),
    .Q_N(_05815_),
    .Q(\shift_storage.storage[504] ));
 sg13g2_dfrbp_1 \shift_storage.storage[505]$_SDFFE_PN0P_  (.CLK(clknet_leaf_258_clk_p2c),
    .RESET_B(net1929),
    .D(_01153_),
    .Q_N(_05814_),
    .Q(\shift_storage.storage[505] ));
 sg13g2_dfrbp_1 \shift_storage.storage[506]$_SDFFE_PN0P_  (.CLK(clknet_leaf_256_clk_p2c),
    .RESET_B(net1930),
    .D(_01154_),
    .Q_N(_05813_),
    .Q(\shift_storage.storage[506] ));
 sg13g2_dfrbp_1 \shift_storage.storage[507]$_SDFFE_PN0P_  (.CLK(clknet_leaf_256_clk_p2c),
    .RESET_B(net1931),
    .D(_01155_),
    .Q_N(_05812_),
    .Q(\shift_storage.storage[507] ));
 sg13g2_dfrbp_1 \shift_storage.storage[508]$_SDFFE_PN0P_  (.CLK(clknet_leaf_256_clk_p2c),
    .RESET_B(net1932),
    .D(_01156_),
    .Q_N(_05811_),
    .Q(\shift_storage.storage[508] ));
 sg13g2_dfrbp_1 \shift_storage.storage[509]$_SDFFE_PN0P_  (.CLK(clknet_leaf_256_clk_p2c),
    .RESET_B(net1933),
    .D(_01157_),
    .Q_N(_05810_),
    .Q(\shift_storage.storage[509] ));
 sg13g2_dfrbp_1 \shift_storage.storage[50]$_SDFFE_PN0P_  (.CLK(clknet_leaf_39_clk_p2c),
    .RESET_B(net1934),
    .D(_01158_),
    .Q_N(_05809_),
    .Q(\shift_storage.storage[50] ));
 sg13g2_dfrbp_1 \shift_storage.storage[510]$_SDFFE_PN0P_  (.CLK(clknet_leaf_255_clk_p2c),
    .RESET_B(net1935),
    .D(_01159_),
    .Q_N(_05808_),
    .Q(\shift_storage.storage[510] ));
 sg13g2_dfrbp_1 \shift_storage.storage[511]$_SDFFE_PN0P_  (.CLK(clknet_leaf_255_clk_p2c),
    .RESET_B(net1936),
    .D(_01160_),
    .Q_N(_05807_),
    .Q(\shift_storage.storage[511] ));
 sg13g2_dfrbp_1 \shift_storage.storage[512]$_SDFFE_PN0P_  (.CLK(clknet_leaf_255_clk_p2c),
    .RESET_B(net1937),
    .D(_01161_),
    .Q_N(_05806_),
    .Q(\shift_storage.storage[512] ));
 sg13g2_dfrbp_1 \shift_storage.storage[513]$_SDFFE_PN0P_  (.CLK(clknet_leaf_255_clk_p2c),
    .RESET_B(net1938),
    .D(_01162_),
    .Q_N(_05805_),
    .Q(\shift_storage.storage[513] ));
 sg13g2_dfrbp_1 \shift_storage.storage[514]$_SDFFE_PN0P_  (.CLK(clknet_leaf_255_clk_p2c),
    .RESET_B(net1939),
    .D(_01163_),
    .Q_N(_05804_),
    .Q(\shift_storage.storage[514] ));
 sg13g2_dfrbp_1 \shift_storage.storage[515]$_SDFFE_PN0P_  (.CLK(clknet_leaf_277_clk_p2c),
    .RESET_B(net1940),
    .D(_01164_),
    .Q_N(_05803_),
    .Q(\shift_storage.storage[515] ));
 sg13g2_dfrbp_1 \shift_storage.storage[516]$_SDFFE_PN0P_  (.CLK(clknet_leaf_277_clk_p2c),
    .RESET_B(net1941),
    .D(_01165_),
    .Q_N(_05802_),
    .Q(\shift_storage.storage[516] ));
 sg13g2_dfrbp_1 \shift_storage.storage[517]$_SDFFE_PN0P_  (.CLK(clknet_leaf_277_clk_p2c),
    .RESET_B(net1942),
    .D(_01166_),
    .Q_N(_05801_),
    .Q(\shift_storage.storage[517] ));
 sg13g2_dfrbp_1 \shift_storage.storage[518]$_SDFFE_PN0P_  (.CLK(clknet_leaf_278_clk_p2c),
    .RESET_B(net1943),
    .D(_01167_),
    .Q_N(_05800_),
    .Q(\shift_storage.storage[518] ));
 sg13g2_dfrbp_1 \shift_storage.storage[519]$_SDFFE_PN0P_  (.CLK(clknet_leaf_278_clk_p2c),
    .RESET_B(net1944),
    .D(_01168_),
    .Q_N(_05799_),
    .Q(\shift_storage.storage[519] ));
 sg13g2_dfrbp_1 \shift_storage.storage[51]$_SDFFE_PN0P_  (.CLK(clknet_leaf_40_clk_p2c),
    .RESET_B(net1945),
    .D(_01169_),
    .Q_N(_05798_),
    .Q(\shift_storage.storage[51] ));
 sg13g2_dfrbp_1 \shift_storage.storage[520]$_SDFFE_PN0P_  (.CLK(clknet_leaf_278_clk_p2c),
    .RESET_B(net1946),
    .D(_01170_),
    .Q_N(_05797_),
    .Q(\shift_storage.storage[520] ));
 sg13g2_dfrbp_1 \shift_storage.storage[521]$_SDFFE_PN0P_  (.CLK(clknet_leaf_278_clk_p2c),
    .RESET_B(net1947),
    .D(_01171_),
    .Q_N(_05796_),
    .Q(\shift_storage.storage[521] ));
 sg13g2_dfrbp_1 \shift_storage.storage[522]$_SDFFE_PN0P_  (.CLK(clknet_leaf_4_clk_p2c),
    .RESET_B(net1948),
    .D(_01172_),
    .Q_N(_05795_),
    .Q(\shift_storage.storage[522] ));
 sg13g2_dfrbp_1 \shift_storage.storage[523]$_SDFFE_PN0P_  (.CLK(clknet_leaf_278_clk_p2c),
    .RESET_B(net1949),
    .D(_01173_),
    .Q_N(_05794_),
    .Q(\shift_storage.storage[523] ));
 sg13g2_dfrbp_1 \shift_storage.storage[524]$_SDFFE_PN0P_  (.CLK(clknet_leaf_3_clk_p2c),
    .RESET_B(net1950),
    .D(_01174_),
    .Q_N(_05793_),
    .Q(\shift_storage.storage[524] ));
 sg13g2_dfrbp_1 \shift_storage.storage[525]$_SDFFE_PN0P_  (.CLK(clknet_leaf_4_clk_p2c),
    .RESET_B(net1951),
    .D(_01175_),
    .Q_N(_05792_),
    .Q(\shift_storage.storage[525] ));
 sg13g2_dfrbp_1 \shift_storage.storage[526]$_SDFFE_PN0P_  (.CLK(clknet_leaf_4_clk_p2c),
    .RESET_B(net1952),
    .D(_01176_),
    .Q_N(_05791_),
    .Q(\shift_storage.storage[526] ));
 sg13g2_dfrbp_1 \shift_storage.storage[527]$_SDFFE_PN0P_  (.CLK(clknet_leaf_4_clk_p2c),
    .RESET_B(net1953),
    .D(_01177_),
    .Q_N(_05790_),
    .Q(\shift_storage.storage[527] ));
 sg13g2_dfrbp_1 \shift_storage.storage[528]$_SDFFE_PN0P_  (.CLK(clknet_leaf_5_clk_p2c),
    .RESET_B(net1954),
    .D(_01178_),
    .Q_N(_05789_),
    .Q(\shift_storage.storage[528] ));
 sg13g2_dfrbp_1 \shift_storage.storage[529]$_SDFFE_PN0P_  (.CLK(clknet_leaf_4_clk_p2c),
    .RESET_B(net1955),
    .D(_01179_),
    .Q_N(_05788_),
    .Q(\shift_storage.storage[529] ));
 sg13g2_dfrbp_1 \shift_storage.storage[52]$_SDFFE_PN0P_  (.CLK(clknet_leaf_40_clk_p2c),
    .RESET_B(net1956),
    .D(_01180_),
    .Q_N(_05787_),
    .Q(\shift_storage.storage[52] ));
 sg13g2_dfrbp_1 \shift_storage.storage[530]$_SDFFE_PN0P_  (.CLK(clknet_leaf_4_clk_p2c),
    .RESET_B(net1957),
    .D(_01181_),
    .Q_N(_05786_),
    .Q(\shift_storage.storage[530] ));
 sg13g2_dfrbp_1 \shift_storage.storage[531]$_SDFFE_PN0P_  (.CLK(clknet_leaf_3_clk_p2c),
    .RESET_B(net1958),
    .D(_01182_),
    .Q_N(_05785_),
    .Q(\shift_storage.storage[531] ));
 sg13g2_dfrbp_1 \shift_storage.storage[532]$_SDFFE_PN0P_  (.CLK(clknet_leaf_1_clk_p2c),
    .RESET_B(net1959),
    .D(_01183_),
    .Q_N(_05784_),
    .Q(\shift_storage.storage[532] ));
 sg13g2_dfrbp_1 \shift_storage.storage[533]$_SDFFE_PN0P_  (.CLK(clknet_leaf_1_clk_p2c),
    .RESET_B(net1960),
    .D(_01184_),
    .Q_N(_05783_),
    .Q(\shift_storage.storage[533] ));
 sg13g2_dfrbp_1 \shift_storage.storage[534]$_SDFFE_PN0P_  (.CLK(clknet_leaf_1_clk_p2c),
    .RESET_B(net1961),
    .D(_01185_),
    .Q_N(_05782_),
    .Q(\shift_storage.storage[534] ));
 sg13g2_dfrbp_1 \shift_storage.storage[535]$_SDFFE_PN0P_  (.CLK(clknet_leaf_1_clk_p2c),
    .RESET_B(net1962),
    .D(_01186_),
    .Q_N(_05781_),
    .Q(\shift_storage.storage[535] ));
 sg13g2_dfrbp_1 \shift_storage.storage[536]$_SDFFE_PN0P_  (.CLK(clknet_leaf_1_clk_p2c),
    .RESET_B(net1963),
    .D(_01187_),
    .Q_N(_05780_),
    .Q(\shift_storage.storage[536] ));
 sg13g2_dfrbp_1 \shift_storage.storage[537]$_SDFFE_PN0P_  (.CLK(clknet_leaf_1_clk_p2c),
    .RESET_B(net1964),
    .D(_01188_),
    .Q_N(_05779_),
    .Q(\shift_storage.storage[537] ));
 sg13g2_dfrbp_1 \shift_storage.storage[538]$_SDFFE_PN0P_  (.CLK(clknet_leaf_0_clk_p2c),
    .RESET_B(net1965),
    .D(_01189_),
    .Q_N(_05778_),
    .Q(\shift_storage.storage[538] ));
 sg13g2_dfrbp_1 \shift_storage.storage[539]$_SDFFE_PN0P_  (.CLK(clknet_leaf_0_clk_p2c),
    .RESET_B(net1966),
    .D(_01190_),
    .Q_N(_05777_),
    .Q(\shift_storage.storage[539] ));
 sg13g2_dfrbp_1 \shift_storage.storage[53]$_SDFFE_PN0P_  (.CLK(clknet_leaf_40_clk_p2c),
    .RESET_B(net1967),
    .D(_01191_),
    .Q_N(_05776_),
    .Q(\shift_storage.storage[53] ));
 sg13g2_dfrbp_1 \shift_storage.storage[540]$_SDFFE_PN0P_  (.CLK(clknet_leaf_0_clk_p2c),
    .RESET_B(net1968),
    .D(_01192_),
    .Q_N(_05775_),
    .Q(\shift_storage.storage[540] ));
 sg13g2_dfrbp_1 \shift_storage.storage[541]$_SDFFE_PN0P_  (.CLK(clknet_leaf_0_clk_p2c),
    .RESET_B(net1969),
    .D(_01193_),
    .Q_N(_05774_),
    .Q(\shift_storage.storage[541] ));
 sg13g2_dfrbp_1 \shift_storage.storage[542]$_SDFFE_PN0P_  (.CLK(clknet_leaf_0_clk_p2c),
    .RESET_B(net1970),
    .D(_01194_),
    .Q_N(_05773_),
    .Q(\shift_storage.storage[542] ));
 sg13g2_dfrbp_1 \shift_storage.storage[543]$_SDFFE_PN0P_  (.CLK(clknet_leaf_0_clk_p2c),
    .RESET_B(net1971),
    .D(_01195_),
    .Q_N(_05772_),
    .Q(\shift_storage.storage[543] ));
 sg13g2_dfrbp_1 \shift_storage.storage[544]$_SDFFE_PN0P_  (.CLK(clknet_leaf_0_clk_p2c),
    .RESET_B(net1972),
    .D(_01196_),
    .Q_N(_05771_),
    .Q(\shift_storage.storage[544] ));
 sg13g2_dfrbp_1 \shift_storage.storage[545]$_SDFFE_PN0P_  (.CLK(clknet_leaf_1_clk_p2c),
    .RESET_B(net1973),
    .D(_01197_),
    .Q_N(_05770_),
    .Q(\shift_storage.storage[545] ));
 sg13g2_dfrbp_1 \shift_storage.storage[546]$_SDFFE_PN0P_  (.CLK(clknet_leaf_293_clk_p2c),
    .RESET_B(net1974),
    .D(_01198_),
    .Q_N(_05769_),
    .Q(\shift_storage.storage[546] ));
 sg13g2_dfrbp_1 \shift_storage.storage[547]$_SDFFE_PN0P_  (.CLK(clknet_leaf_293_clk_p2c),
    .RESET_B(net1975),
    .D(_01199_),
    .Q_N(_05768_),
    .Q(\shift_storage.storage[547] ));
 sg13g2_dfrbp_1 \shift_storage.storage[548]$_SDFFE_PN0P_  (.CLK(clknet_leaf_293_clk_p2c),
    .RESET_B(net1976),
    .D(_01200_),
    .Q_N(_05767_),
    .Q(\shift_storage.storage[548] ));
 sg13g2_dfrbp_1 \shift_storage.storage[549]$_SDFFE_PN0P_  (.CLK(clknet_leaf_292_clk_p2c),
    .RESET_B(net1977),
    .D(_01201_),
    .Q_N(_05766_),
    .Q(\shift_storage.storage[549] ));
 sg13g2_dfrbp_1 \shift_storage.storage[54]$_SDFFE_PN0P_  (.CLK(clknet_leaf_37_clk_p2c),
    .RESET_B(net1978),
    .D(_01202_),
    .Q_N(_05765_),
    .Q(\shift_storage.storage[54] ));
 sg13g2_dfrbp_1 \shift_storage.storage[550]$_SDFFE_PN0P_  (.CLK(clknet_leaf_292_clk_p2c),
    .RESET_B(net1979),
    .D(_01203_),
    .Q_N(_05764_),
    .Q(\shift_storage.storage[550] ));
 sg13g2_dfrbp_1 \shift_storage.storage[551]$_SDFFE_PN0P_  (.CLK(clknet_leaf_292_clk_p2c),
    .RESET_B(net1980),
    .D(_01204_),
    .Q_N(_05763_),
    .Q(\shift_storage.storage[551] ));
 sg13g2_dfrbp_1 \shift_storage.storage[552]$_SDFFE_PN0P_  (.CLK(clknet_leaf_293_clk_p2c),
    .RESET_B(net1981),
    .D(_01205_),
    .Q_N(_05762_),
    .Q(\shift_storage.storage[552] ));
 sg13g2_dfrbp_1 \shift_storage.storage[553]$_SDFFE_PN0P_  (.CLK(clknet_leaf_293_clk_p2c),
    .RESET_B(net1982),
    .D(_01206_),
    .Q_N(_05761_),
    .Q(\shift_storage.storage[553] ));
 sg13g2_dfrbp_1 \shift_storage.storage[554]$_SDFFE_PN0P_  (.CLK(clknet_leaf_293_clk_p2c),
    .RESET_B(net1983),
    .D(_01207_),
    .Q_N(_05760_),
    .Q(\shift_storage.storage[554] ));
 sg13g2_dfrbp_1 \shift_storage.storage[555]$_SDFFE_PN0P_  (.CLK(clknet_leaf_2_clk_p2c),
    .RESET_B(net1984),
    .D(_01208_),
    .Q_N(_05759_),
    .Q(\shift_storage.storage[555] ));
 sg13g2_dfrbp_1 \shift_storage.storage[556]$_SDFFE_PN0P_  (.CLK(clknet_leaf_2_clk_p2c),
    .RESET_B(net1985),
    .D(_01209_),
    .Q_N(_05758_),
    .Q(\shift_storage.storage[556] ));
 sg13g2_dfrbp_1 \shift_storage.storage[557]$_SDFFE_PN0P_  (.CLK(clknet_leaf_2_clk_p2c),
    .RESET_B(net1986),
    .D(_01210_),
    .Q_N(_05757_),
    .Q(\shift_storage.storage[557] ));
 sg13g2_dfrbp_1 \shift_storage.storage[558]$_SDFFE_PN0P_  (.CLK(clknet_leaf_2_clk_p2c),
    .RESET_B(net1987),
    .D(_01211_),
    .Q_N(_05756_),
    .Q(\shift_storage.storage[558] ));
 sg13g2_dfrbp_1 \shift_storage.storage[559]$_SDFFE_PN0P_  (.CLK(clknet_leaf_3_clk_p2c),
    .RESET_B(net1988),
    .D(_01212_),
    .Q_N(_05755_),
    .Q(\shift_storage.storage[559] ));
 sg13g2_dfrbp_1 \shift_storage.storage[55]$_SDFFE_PN0P_  (.CLK(clknet_leaf_37_clk_p2c),
    .RESET_B(net1989),
    .D(_01213_),
    .Q_N(_05754_),
    .Q(\shift_storage.storage[55] ));
 sg13g2_dfrbp_1 \shift_storage.storage[560]$_SDFFE_PN0P_  (.CLK(clknet_leaf_2_clk_p2c),
    .RESET_B(net1990),
    .D(_01214_),
    .Q_N(_05753_),
    .Q(\shift_storage.storage[560] ));
 sg13g2_dfrbp_1 \shift_storage.storage[561]$_SDFFE_PN0P_  (.CLK(clknet_leaf_3_clk_p2c),
    .RESET_B(net1991),
    .D(_01215_),
    .Q_N(_05752_),
    .Q(\shift_storage.storage[561] ));
 sg13g2_dfrbp_1 \shift_storage.storage[562]$_SDFFE_PN0P_  (.CLK(clknet_leaf_2_clk_p2c),
    .RESET_B(net1992),
    .D(_01216_),
    .Q_N(_05751_),
    .Q(\shift_storage.storage[562] ));
 sg13g2_dfrbp_1 \shift_storage.storage[563]$_SDFFE_PN0P_  (.CLK(clknet_leaf_3_clk_p2c),
    .RESET_B(net1993),
    .D(_01217_),
    .Q_N(_05750_),
    .Q(\shift_storage.storage[563] ));
 sg13g2_dfrbp_1 \shift_storage.storage[564]$_SDFFE_PN0P_  (.CLK(clknet_leaf_280_clk_p2c),
    .RESET_B(net1994),
    .D(_01218_),
    .Q_N(_05749_),
    .Q(\shift_storage.storage[564] ));
 sg13g2_dfrbp_1 \shift_storage.storage[565]$_SDFFE_PN0P_  (.CLK(clknet_leaf_280_clk_p2c),
    .RESET_B(net1995),
    .D(_01219_),
    .Q_N(_05748_),
    .Q(\shift_storage.storage[565] ));
 sg13g2_dfrbp_1 \shift_storage.storage[566]$_SDFFE_PN0P_  (.CLK(clknet_leaf_280_clk_p2c),
    .RESET_B(net1996),
    .D(_01220_),
    .Q_N(_05747_),
    .Q(\shift_storage.storage[566] ));
 sg13g2_dfrbp_1 \shift_storage.storage[567]$_SDFFE_PN0P_  (.CLK(clknet_leaf_280_clk_p2c),
    .RESET_B(net1997),
    .D(_01221_),
    .Q_N(_05746_),
    .Q(\shift_storage.storage[567] ));
 sg13g2_dfrbp_1 \shift_storage.storage[568]$_SDFFE_PN0P_  (.CLK(clknet_leaf_280_clk_p2c),
    .RESET_B(net1998),
    .D(_01222_),
    .Q_N(_05745_),
    .Q(\shift_storage.storage[568] ));
 sg13g2_dfrbp_1 \shift_storage.storage[569]$_SDFFE_PN0P_  (.CLK(clknet_leaf_280_clk_p2c),
    .RESET_B(net1999),
    .D(_01223_),
    .Q_N(_05744_),
    .Q(\shift_storage.storage[569] ));
 sg13g2_dfrbp_1 \shift_storage.storage[56]$_SDFFE_PN0P_  (.CLK(clknet_leaf_38_clk_p2c),
    .RESET_B(net2000),
    .D(_01224_),
    .Q_N(_05743_),
    .Q(\shift_storage.storage[56] ));
 sg13g2_dfrbp_1 \shift_storage.storage[570]$_SDFFE_PN0P_  (.CLK(clknet_leaf_286_clk_p2c),
    .RESET_B(net2001),
    .D(_01225_),
    .Q_N(_05742_),
    .Q(\shift_storage.storage[570] ));
 sg13g2_dfrbp_1 \shift_storage.storage[571]$_SDFFE_PN0P_  (.CLK(clknet_leaf_286_clk_p2c),
    .RESET_B(net2002),
    .D(_01226_),
    .Q_N(_05741_),
    .Q(\shift_storage.storage[571] ));
 sg13g2_dfrbp_1 \shift_storage.storage[572]$_SDFFE_PN0P_  (.CLK(clknet_leaf_286_clk_p2c),
    .RESET_B(net2003),
    .D(_01227_),
    .Q_N(_05740_),
    .Q(\shift_storage.storage[572] ));
 sg13g2_dfrbp_1 \shift_storage.storage[573]$_SDFFE_PN0P_  (.CLK(clknet_leaf_285_clk_p2c),
    .RESET_B(net2004),
    .D(_01228_),
    .Q_N(_05739_),
    .Q(\shift_storage.storage[573] ));
 sg13g2_dfrbp_1 \shift_storage.storage[574]$_SDFFE_PN0P_  (.CLK(clknet_leaf_285_clk_p2c),
    .RESET_B(net2005),
    .D(_01229_),
    .Q_N(_05738_),
    .Q(\shift_storage.storage[574] ));
 sg13g2_dfrbp_1 \shift_storage.storage[575]$_SDFFE_PN0P_  (.CLK(clknet_leaf_287_clk_p2c),
    .RESET_B(net2006),
    .D(_01230_),
    .Q_N(_05737_),
    .Q(\shift_storage.storage[575] ));
 sg13g2_dfrbp_1 \shift_storage.storage[576]$_SDFFE_PN0P_  (.CLK(clknet_leaf_287_clk_p2c),
    .RESET_B(net2007),
    .D(_01231_),
    .Q_N(_05736_),
    .Q(\shift_storage.storage[576] ));
 sg13g2_dfrbp_1 \shift_storage.storage[577]$_SDFFE_PN0P_  (.CLK(clknet_leaf_287_clk_p2c),
    .RESET_B(net2008),
    .D(_01232_),
    .Q_N(_05735_),
    .Q(\shift_storage.storage[577] ));
 sg13g2_dfrbp_1 \shift_storage.storage[578]$_SDFFE_PN0P_  (.CLK(clknet_leaf_286_clk_p2c),
    .RESET_B(net2009),
    .D(_01233_),
    .Q_N(_05734_),
    .Q(\shift_storage.storage[578] ));
 sg13g2_dfrbp_1 \shift_storage.storage[579]$_SDFFE_PN0P_  (.CLK(clknet_leaf_286_clk_p2c),
    .RESET_B(net2010),
    .D(_01234_),
    .Q_N(_05733_),
    .Q(\shift_storage.storage[579] ));
 sg13g2_dfrbp_1 \shift_storage.storage[57]$_SDFFE_PN0P_  (.CLK(clknet_leaf_38_clk_p2c),
    .RESET_B(net2011),
    .D(_01235_),
    .Q_N(_05732_),
    .Q(\shift_storage.storage[57] ));
 sg13g2_dfrbp_1 \shift_storage.storage[580]$_SDFFE_PN0P_  (.CLK(clknet_leaf_286_clk_p2c),
    .RESET_B(net2012),
    .D(_01236_),
    .Q_N(_05731_),
    .Q(\shift_storage.storage[580] ));
 sg13g2_dfrbp_1 \shift_storage.storage[581]$_SDFFE_PN0P_  (.CLK(clknet_leaf_286_clk_p2c),
    .RESET_B(net2013),
    .D(_01237_),
    .Q_N(_05730_),
    .Q(\shift_storage.storage[581] ));
 sg13g2_dfrbp_1 \shift_storage.storage[582]$_SDFFE_PN0P_  (.CLK(clknet_leaf_292_clk_p2c),
    .RESET_B(net2014),
    .D(_01238_),
    .Q_N(_05729_),
    .Q(\shift_storage.storage[582] ));
 sg13g2_dfrbp_1 \shift_storage.storage[583]$_SDFFE_PN0P_  (.CLK(clknet_leaf_292_clk_p2c),
    .RESET_B(net2015),
    .D(_01239_),
    .Q_N(_05728_),
    .Q(\shift_storage.storage[583] ));
 sg13g2_dfrbp_1 \shift_storage.storage[584]$_SDFFE_PN0P_  (.CLK(clknet_leaf_292_clk_p2c),
    .RESET_B(net2016),
    .D(_01240_),
    .Q_N(_05727_),
    .Q(\shift_storage.storage[584] ));
 sg13g2_dfrbp_1 \shift_storage.storage[585]$_SDFFE_PN0P_  (.CLK(clknet_leaf_291_clk_p2c),
    .RESET_B(net2017),
    .D(_01241_),
    .Q_N(_05726_),
    .Q(\shift_storage.storage[585] ));
 sg13g2_dfrbp_1 \shift_storage.storage[586]$_SDFFE_PN0P_  (.CLK(clknet_leaf_291_clk_p2c),
    .RESET_B(net2018),
    .D(_01242_),
    .Q_N(_05725_),
    .Q(\shift_storage.storage[586] ));
 sg13g2_dfrbp_1 \shift_storage.storage[587]$_SDFFE_PN0P_  (.CLK(clknet_leaf_291_clk_p2c),
    .RESET_B(net2019),
    .D(_01243_),
    .Q_N(_05724_),
    .Q(\shift_storage.storage[587] ));
 sg13g2_dfrbp_1 \shift_storage.storage[588]$_SDFFE_PN0P_  (.CLK(clknet_leaf_291_clk_p2c),
    .RESET_B(net2020),
    .D(_01244_),
    .Q_N(_05723_),
    .Q(\shift_storage.storage[588] ));
 sg13g2_dfrbp_1 \shift_storage.storage[589]$_SDFFE_PN0P_  (.CLK(clknet_leaf_291_clk_p2c),
    .RESET_B(net2021),
    .D(_01245_),
    .Q_N(_05722_),
    .Q(\shift_storage.storage[589] ));
 sg13g2_dfrbp_1 \shift_storage.storage[58]$_SDFFE_PN0P_  (.CLK(clknet_leaf_105_clk_p2c),
    .RESET_B(net2022),
    .D(_01246_),
    .Q_N(_05721_),
    .Q(\shift_storage.storage[58] ));
 sg13g2_dfrbp_1 \shift_storage.storage[590]$_SDFFE_PN0P_  (.CLK(clknet_leaf_290_clk_p2c),
    .RESET_B(net2023),
    .D(_01247_),
    .Q_N(_05720_),
    .Q(\shift_storage.storage[590] ));
 sg13g2_dfrbp_1 \shift_storage.storage[591]$_SDFFE_PN0P_  (.CLK(clknet_leaf_290_clk_p2c),
    .RESET_B(net2024),
    .D(_01248_),
    .Q_N(_05719_),
    .Q(\shift_storage.storage[591] ));
 sg13g2_dfrbp_1 \shift_storage.storage[592]$_SDFFE_PN0P_  (.CLK(clknet_leaf_290_clk_p2c),
    .RESET_B(net2025),
    .D(_01249_),
    .Q_N(_05718_),
    .Q(\shift_storage.storage[592] ));
 sg13g2_dfrbp_1 \shift_storage.storage[593]$_SDFFE_PN0P_  (.CLK(clknet_leaf_289_clk_p2c),
    .RESET_B(net2026),
    .D(_01250_),
    .Q_N(_05717_),
    .Q(\shift_storage.storage[593] ));
 sg13g2_dfrbp_1 \shift_storage.storage[594]$_SDFFE_PN0P_  (.CLK(clknet_leaf_289_clk_p2c),
    .RESET_B(net2027),
    .D(_01251_),
    .Q_N(_05716_),
    .Q(\shift_storage.storage[594] ));
 sg13g2_dfrbp_1 \shift_storage.storage[595]$_SDFFE_PN0P_  (.CLK(clknet_leaf_289_clk_p2c),
    .RESET_B(net2028),
    .D(_01252_),
    .Q_N(_05715_),
    .Q(\shift_storage.storage[595] ));
 sg13g2_dfrbp_1 \shift_storage.storage[596]$_SDFFE_PN0P_  (.CLK(clknet_leaf_289_clk_p2c),
    .RESET_B(net2029),
    .D(_01253_),
    .Q_N(_05714_),
    .Q(\shift_storage.storage[596] ));
 sg13g2_dfrbp_1 \shift_storage.storage[597]$_SDFFE_PN0P_  (.CLK(clknet_leaf_289_clk_p2c),
    .RESET_B(net2030),
    .D(_01254_),
    .Q_N(_05713_),
    .Q(\shift_storage.storage[597] ));
 sg13g2_dfrbp_1 \shift_storage.storage[598]$_SDFFE_PN0P_  (.CLK(clknet_leaf_289_clk_p2c),
    .RESET_B(net2031),
    .D(_01255_),
    .Q_N(_05712_),
    .Q(\shift_storage.storage[598] ));
 sg13g2_dfrbp_1 \shift_storage.storage[599]$_SDFFE_PN0P_  (.CLK(clknet_leaf_290_clk_p2c),
    .RESET_B(net2032),
    .D(_01256_),
    .Q_N(_05711_),
    .Q(\shift_storage.storage[599] ));
 sg13g2_dfrbp_1 \shift_storage.storage[59]$_SDFFE_PN0P_  (.CLK(clknet_leaf_38_clk_p2c),
    .RESET_B(net2033),
    .D(_01257_),
    .Q_N(_05710_),
    .Q(\shift_storage.storage[59] ));
 sg13g2_dfrbp_1 \shift_storage.storage[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_76_clk_p2c),
    .RESET_B(net2034),
    .D(_01258_),
    .Q_N(_05709_),
    .Q(\shift_storage.storage[5] ));
 sg13g2_dfrbp_1 \shift_storage.storage[600]$_SDFFE_PN0P_  (.CLK(clknet_leaf_290_clk_p2c),
    .RESET_B(net2035),
    .D(_01259_),
    .Q_N(_05708_),
    .Q(\shift_storage.storage[600] ));
 sg13g2_dfrbp_1 \shift_storage.storage[601]$_SDFFE_PN0P_  (.CLK(clknet_leaf_290_clk_p2c),
    .RESET_B(net2036),
    .D(_01260_),
    .Q_N(_05707_),
    .Q(\shift_storage.storage[601] ));
 sg13g2_dfrbp_1 \shift_storage.storage[602]$_SDFFE_PN0P_  (.CLK(clknet_leaf_287_clk_p2c),
    .RESET_B(net2037),
    .D(_01261_),
    .Q_N(_05706_),
    .Q(\shift_storage.storage[602] ));
 sg13g2_dfrbp_1 \shift_storage.storage[603]$_SDFFE_PN0P_  (.CLK(clknet_leaf_287_clk_p2c),
    .RESET_B(net2038),
    .D(_01262_),
    .Q_N(_05705_),
    .Q(\shift_storage.storage[603] ));
 sg13g2_dfrbp_1 \shift_storage.storage[604]$_SDFFE_PN0P_  (.CLK(clknet_leaf_288_clk_p2c),
    .RESET_B(net2039),
    .D(_01263_),
    .Q_N(_05704_),
    .Q(\shift_storage.storage[604] ));
 sg13g2_dfrbp_1 \shift_storage.storage[605]$_SDFFE_PN0P_  (.CLK(clknet_leaf_288_clk_p2c),
    .RESET_B(net2040),
    .D(_01264_),
    .Q_N(_05703_),
    .Q(\shift_storage.storage[605] ));
 sg13g2_dfrbp_1 \shift_storage.storage[606]$_SDFFE_PN0P_  (.CLK(clknet_leaf_288_clk_p2c),
    .RESET_B(net2041),
    .D(_01265_),
    .Q_N(_05702_),
    .Q(\shift_storage.storage[606] ));
 sg13g2_dfrbp_1 \shift_storage.storage[607]$_SDFFE_PN0P_  (.CLK(clknet_leaf_288_clk_p2c),
    .RESET_B(net2042),
    .D(_01266_),
    .Q_N(_05701_),
    .Q(\shift_storage.storage[607] ));
 sg13g2_dfrbp_1 \shift_storage.storage[608]$_SDFFE_PN0P_  (.CLK(clknet_leaf_288_clk_p2c),
    .RESET_B(net2043),
    .D(_01267_),
    .Q_N(_05700_),
    .Q(\shift_storage.storage[608] ));
 sg13g2_dfrbp_1 \shift_storage.storage[609]$_SDFFE_PN0P_  (.CLK(clknet_leaf_288_clk_p2c),
    .RESET_B(net2044),
    .D(_01268_),
    .Q_N(_05699_),
    .Q(\shift_storage.storage[609] ));
 sg13g2_dfrbp_1 \shift_storage.storage[60]$_SDFFE_PN0P_  (.CLK(clknet_leaf_38_clk_p2c),
    .RESET_B(net2045),
    .D(_01269_),
    .Q_N(_05698_),
    .Q(\shift_storage.storage[60] ));
 sg13g2_dfrbp_1 \shift_storage.storage[610]$_SDFFE_PN0P_  (.CLK(clknet_leaf_285_clk_p2c),
    .RESET_B(net2046),
    .D(_01270_),
    .Q_N(_05697_),
    .Q(\shift_storage.storage[610] ));
 sg13g2_dfrbp_1 \shift_storage.storage[611]$_SDFFE_PN0P_  (.CLK(clknet_leaf_285_clk_p2c),
    .RESET_B(net2047),
    .D(_01271_),
    .Q_N(_05696_),
    .Q(\shift_storage.storage[611] ));
 sg13g2_dfrbp_1 \shift_storage.storage[612]$_SDFFE_PN0P_  (.CLK(clknet_leaf_284_clk_p2c),
    .RESET_B(net2048),
    .D(_01272_),
    .Q_N(_05695_),
    .Q(\shift_storage.storage[612] ));
 sg13g2_dfrbp_1 \shift_storage.storage[613]$_SDFFE_PN0P_  (.CLK(clknet_leaf_284_clk_p2c),
    .RESET_B(net2049),
    .D(_01273_),
    .Q_N(_05694_),
    .Q(\shift_storage.storage[613] ));
 sg13g2_dfrbp_1 \shift_storage.storage[614]$_SDFFE_PN0P_  (.CLK(clknet_leaf_284_clk_p2c),
    .RESET_B(net2050),
    .D(_01274_),
    .Q_N(_05693_),
    .Q(\shift_storage.storage[614] ));
 sg13g2_dfrbp_1 \shift_storage.storage[615]$_SDFFE_PN0P_  (.CLK(clknet_leaf_284_clk_p2c),
    .RESET_B(net2051),
    .D(_01275_),
    .Q_N(_05692_),
    .Q(\shift_storage.storage[615] ));
 sg13g2_dfrbp_1 \shift_storage.storage[616]$_SDFFE_PN0P_  (.CLK(clknet_leaf_284_clk_p2c),
    .RESET_B(net2052),
    .D(_01276_),
    .Q_N(_05691_),
    .Q(\shift_storage.storage[616] ));
 sg13g2_dfrbp_1 \shift_storage.storage[617]$_SDFFE_PN0P_  (.CLK(clknet_leaf_284_clk_p2c),
    .RESET_B(net2053),
    .D(_01277_),
    .Q_N(_05690_),
    .Q(\shift_storage.storage[617] ));
 sg13g2_dfrbp_1 \shift_storage.storage[618]$_SDFFE_PN0P_  (.CLK(clknet_leaf_283_clk_p2c),
    .RESET_B(net2054),
    .D(_01278_),
    .Q_N(_05689_),
    .Q(\shift_storage.storage[618] ));
 sg13g2_dfrbp_1 \shift_storage.storage[619]$_SDFFE_PN0P_  (.CLK(clknet_leaf_282_clk_p2c),
    .RESET_B(net2055),
    .D(_01279_),
    .Q_N(_05688_),
    .Q(\shift_storage.storage[619] ));
 sg13g2_dfrbp_1 \shift_storage.storage[61]$_SDFFE_PN0P_  (.CLK(clknet_leaf_38_clk_p2c),
    .RESET_B(net2056),
    .D(_01280_),
    .Q_N(_05687_),
    .Q(\shift_storage.storage[61] ));
 sg13g2_dfrbp_1 \shift_storage.storage[620]$_SDFFE_PN0P_  (.CLK(clknet_leaf_285_clk_p2c),
    .RESET_B(net2057),
    .D(_01281_),
    .Q_N(_05686_),
    .Q(\shift_storage.storage[620] ));
 sg13g2_dfrbp_1 \shift_storage.storage[621]$_SDFFE_PN0P_  (.CLK(clknet_leaf_285_clk_p2c),
    .RESET_B(net2058),
    .D(_01282_),
    .Q_N(_05685_),
    .Q(\shift_storage.storage[621] ));
 sg13g2_dfrbp_1 \shift_storage.storage[622]$_SDFFE_PN0P_  (.CLK(clknet_leaf_281_clk_p2c),
    .RESET_B(net2059),
    .D(_01283_),
    .Q_N(_05684_),
    .Q(\shift_storage.storage[622] ));
 sg13g2_dfrbp_1 \shift_storage.storage[623]$_SDFFE_PN0P_  (.CLK(clknet_leaf_281_clk_p2c),
    .RESET_B(net2060),
    .D(_01284_),
    .Q_N(_05683_),
    .Q(\shift_storage.storage[623] ));
 sg13g2_dfrbp_1 \shift_storage.storage[624]$_SDFFE_PN0P_  (.CLK(clknet_leaf_281_clk_p2c),
    .RESET_B(net2061),
    .D(_01285_),
    .Q_N(_05682_),
    .Q(\shift_storage.storage[624] ));
 sg13g2_dfrbp_1 \shift_storage.storage[625]$_SDFFE_PN0P_  (.CLK(clknet_leaf_281_clk_p2c),
    .RESET_B(net2062),
    .D(_01286_),
    .Q_N(_05681_),
    .Q(\shift_storage.storage[625] ));
 sg13g2_dfrbp_1 \shift_storage.storage[626]$_SDFFE_PN0P_  (.CLK(clknet_leaf_281_clk_p2c),
    .RESET_B(net2063),
    .D(_01287_),
    .Q_N(_05680_),
    .Q(\shift_storage.storage[626] ));
 sg13g2_dfrbp_1 \shift_storage.storage[627]$_SDFFE_PN0P_  (.CLK(clknet_leaf_282_clk_p2c),
    .RESET_B(net2064),
    .D(_01288_),
    .Q_N(_05679_),
    .Q(\shift_storage.storage[627] ));
 sg13g2_dfrbp_1 \shift_storage.storage[628]$_SDFFE_PN0P_  (.CLK(clknet_leaf_282_clk_p2c),
    .RESET_B(net2065),
    .D(_01289_),
    .Q_N(_05678_),
    .Q(\shift_storage.storage[628] ));
 sg13g2_dfrbp_1 \shift_storage.storage[629]$_SDFFE_PN0P_  (.CLK(clknet_leaf_274_clk_p2c),
    .RESET_B(net2066),
    .D(_01290_),
    .Q_N(_05677_),
    .Q(\shift_storage.storage[629] ));
 sg13g2_dfrbp_1 \shift_storage.storage[62]$_SDFFE_PN0P_  (.CLK(clknet_leaf_39_clk_p2c),
    .RESET_B(net2067),
    .D(_01291_),
    .Q_N(_05676_),
    .Q(\shift_storage.storage[62] ));
 sg13g2_dfrbp_1 \shift_storage.storage[630]$_SDFFE_PN0P_  (.CLK(clknet_leaf_276_clk_p2c),
    .RESET_B(net2068),
    .D(_01292_),
    .Q_N(_05675_),
    .Q(\shift_storage.storage[630] ));
 sg13g2_dfrbp_1 \shift_storage.storage[631]$_SDFFE_PN0P_  (.CLK(clknet_leaf_276_clk_p2c),
    .RESET_B(net2069),
    .D(_01293_),
    .Q_N(_05674_),
    .Q(\shift_storage.storage[631] ));
 sg13g2_dfrbp_1 \shift_storage.storage[632]$_SDFFE_PN0P_  (.CLK(clknet_leaf_276_clk_p2c),
    .RESET_B(net2070),
    .D(_01294_),
    .Q_N(_05673_),
    .Q(\shift_storage.storage[632] ));
 sg13g2_dfrbp_1 \shift_storage.storage[633]$_SDFFE_PN0P_  (.CLK(clknet_leaf_279_clk_p2c),
    .RESET_B(net2071),
    .D(_01295_),
    .Q_N(_05672_),
    .Q(\shift_storage.storage[633] ));
 sg13g2_dfrbp_1 \shift_storage.storage[634]$_SDFFE_PN0P_  (.CLK(clknet_leaf_279_clk_p2c),
    .RESET_B(net2072),
    .D(_01296_),
    .Q_N(_05671_),
    .Q(\shift_storage.storage[634] ));
 sg13g2_dfrbp_1 \shift_storage.storage[635]$_SDFFE_PN0P_  (.CLK(clknet_leaf_279_clk_p2c),
    .RESET_B(net2073),
    .D(_01297_),
    .Q_N(_05670_),
    .Q(\shift_storage.storage[635] ));
 sg13g2_dfrbp_1 \shift_storage.storage[636]$_SDFFE_PN0P_  (.CLK(clknet_leaf_279_clk_p2c),
    .RESET_B(net2074),
    .D(_01298_),
    .Q_N(_05669_),
    .Q(\shift_storage.storage[636] ));
 sg13g2_dfrbp_1 \shift_storage.storage[637]$_SDFFE_PN0P_  (.CLK(clknet_leaf_278_clk_p2c),
    .RESET_B(net2075),
    .D(_01299_),
    .Q_N(_05668_),
    .Q(\shift_storage.storage[637] ));
 sg13g2_dfrbp_1 \shift_storage.storage[638]$_SDFFE_PN0P_  (.CLK(clknet_leaf_278_clk_p2c),
    .RESET_B(net2076),
    .D(_01300_),
    .Q_N(_05667_),
    .Q(\shift_storage.storage[638] ));
 sg13g2_dfrbp_1 \shift_storage.storage[639]$_SDFFE_PN0P_  (.CLK(clknet_leaf_279_clk_p2c),
    .RESET_B(net2077),
    .D(_01301_),
    .Q_N(_05666_),
    .Q(\shift_storage.storage[639] ));
 sg13g2_dfrbp_1 \shift_storage.storage[63]$_SDFFE_PN0P_  (.CLK(clknet_leaf_45_clk_p2c),
    .RESET_B(net2078),
    .D(_01302_),
    .Q_N(_05665_),
    .Q(\shift_storage.storage[63] ));
 sg13g2_dfrbp_1 \shift_storage.storage[640]$_SDFFE_PN0P_  (.CLK(clknet_leaf_279_clk_p2c),
    .RESET_B(net2079),
    .D(_01303_),
    .Q_N(_05664_),
    .Q(\shift_storage.storage[640] ));
 sg13g2_dfrbp_1 \shift_storage.storage[641]$_SDFFE_PN0P_  (.CLK(clknet_leaf_276_clk_p2c),
    .RESET_B(net2080),
    .D(_01304_),
    .Q_N(_05663_),
    .Q(\shift_storage.storage[641] ));
 sg13g2_dfrbp_1 \shift_storage.storage[642]$_SDFFE_PN0P_  (.CLK(clknet_leaf_277_clk_p2c),
    .RESET_B(net2081),
    .D(_01305_),
    .Q_N(_05662_),
    .Q(\shift_storage.storage[642] ));
 sg13g2_dfrbp_1 \shift_storage.storage[643]$_SDFFE_PN0P_  (.CLK(clknet_leaf_277_clk_p2c),
    .RESET_B(net2082),
    .D(_01306_),
    .Q_N(_05661_),
    .Q(\shift_storage.storage[643] ));
 sg13g2_dfrbp_1 \shift_storage.storage[644]$_SDFFE_PN0P_  (.CLK(clknet_leaf_277_clk_p2c),
    .RESET_B(net2083),
    .D(_01307_),
    .Q_N(_05660_),
    .Q(\shift_storage.storage[644] ));
 sg13g2_dfrbp_1 \shift_storage.storage[645]$_SDFFE_PN0P_  (.CLK(clknet_leaf_277_clk_p2c),
    .RESET_B(net2084),
    .D(_01308_),
    .Q_N(_05659_),
    .Q(\shift_storage.storage[645] ));
 sg13g2_dfrbp_1 \shift_storage.storage[646]$_SDFFE_PN0P_  (.CLK(clknet_leaf_276_clk_p2c),
    .RESET_B(net2085),
    .D(_01309_),
    .Q_N(_05658_),
    .Q(\shift_storage.storage[646] ));
 sg13g2_dfrbp_1 \shift_storage.storage[647]$_SDFFE_PN0P_  (.CLK(clknet_leaf_275_clk_p2c),
    .RESET_B(net2086),
    .D(_01310_),
    .Q_N(_05657_),
    .Q(\shift_storage.storage[647] ));
 sg13g2_dfrbp_1 \shift_storage.storage[648]$_SDFFE_PN0P_  (.CLK(clknet_leaf_256_clk_p2c),
    .RESET_B(net2087),
    .D(_01311_),
    .Q_N(_05656_),
    .Q(\shift_storage.storage[648] ));
 sg13g2_dfrbp_1 \shift_storage.storage[649]$_SDFFE_PN0P_  (.CLK(clknet_leaf_256_clk_p2c),
    .RESET_B(net2088),
    .D(_01312_),
    .Q_N(_05655_),
    .Q(\shift_storage.storage[649] ));
 sg13g2_dfrbp_1 \shift_storage.storage[64]$_SDFFE_PN0P_  (.CLK(clknet_leaf_45_clk_p2c),
    .RESET_B(net2089),
    .D(_01313_),
    .Q_N(_05654_),
    .Q(\shift_storage.storage[64] ));
 sg13g2_dfrbp_1 \shift_storage.storage[650]$_SDFFE_PN0P_  (.CLK(clknet_leaf_257_clk_p2c),
    .RESET_B(net2090),
    .D(_01314_),
    .Q_N(_05653_),
    .Q(\shift_storage.storage[650] ));
 sg13g2_dfrbp_1 \shift_storage.storage[651]$_SDFFE_PN0P_  (.CLK(clknet_leaf_257_clk_p2c),
    .RESET_B(net2091),
    .D(_01315_),
    .Q_N(_05652_),
    .Q(\shift_storage.storage[651] ));
 sg13g2_dfrbp_1 \shift_storage.storage[652]$_SDFFE_PN0P_  (.CLK(clknet_leaf_275_clk_p2c),
    .RESET_B(net2092),
    .D(_01316_),
    .Q_N(_05651_),
    .Q(\shift_storage.storage[652] ));
 sg13g2_dfrbp_1 \shift_storage.storage[653]$_SDFFE_PN0P_  (.CLK(clknet_leaf_257_clk_p2c),
    .RESET_B(net2093),
    .D(_01317_),
    .Q_N(_05650_),
    .Q(\shift_storage.storage[653] ));
 sg13g2_dfrbp_1 \shift_storage.storage[654]$_SDFFE_PN0P_  (.CLK(clknet_leaf_257_clk_p2c),
    .RESET_B(net2094),
    .D(_01318_),
    .Q_N(_05649_),
    .Q(\shift_storage.storage[654] ));
 sg13g2_dfrbp_1 \shift_storage.storage[655]$_SDFFE_PN0P_  (.CLK(clknet_leaf_257_clk_p2c),
    .RESET_B(net2095),
    .D(_01319_),
    .Q_N(_05648_),
    .Q(\shift_storage.storage[655] ));
 sg13g2_dfrbp_1 \shift_storage.storage[656]$_SDFFE_PN0P_  (.CLK(clknet_leaf_257_clk_p2c),
    .RESET_B(net2096),
    .D(_01320_),
    .Q_N(_05647_),
    .Q(\shift_storage.storage[656] ));
 sg13g2_dfrbp_1 \shift_storage.storage[657]$_SDFFE_PN0P_  (.CLK(clknet_leaf_258_clk_p2c),
    .RESET_B(net2097),
    .D(_01321_),
    .Q_N(_05646_),
    .Q(\shift_storage.storage[657] ));
 sg13g2_dfrbp_1 \shift_storage.storage[658]$_SDFFE_PN0P_  (.CLK(clknet_leaf_258_clk_p2c),
    .RESET_B(net2098),
    .D(_01322_),
    .Q_N(_05645_),
    .Q(\shift_storage.storage[658] ));
 sg13g2_dfrbp_1 \shift_storage.storage[659]$_SDFFE_PN0P_  (.CLK(clknet_leaf_263_clk_p2c),
    .RESET_B(net2099),
    .D(_01323_),
    .Q_N(_05644_),
    .Q(\shift_storage.storage[659] ));
 sg13g2_dfrbp_1 \shift_storage.storage[65]$_SDFFE_PN0P_  (.CLK(clknet_leaf_45_clk_p2c),
    .RESET_B(net2100),
    .D(_01324_),
    .Q_N(_05643_),
    .Q(\shift_storage.storage[65] ));
 sg13g2_dfrbp_1 \shift_storage.storage[660]$_SDFFE_PN0P_  (.CLK(clknet_leaf_263_clk_p2c),
    .RESET_B(net2101),
    .D(_01325_),
    .Q_N(_05642_),
    .Q(\shift_storage.storage[660] ));
 sg13g2_dfrbp_1 \shift_storage.storage[661]$_SDFFE_PN0P_  (.CLK(clknet_leaf_261_clk_p2c),
    .RESET_B(net2102),
    .D(_01326_),
    .Q_N(_05641_),
    .Q(\shift_storage.storage[661] ));
 sg13g2_dfrbp_1 \shift_storage.storage[662]$_SDFFE_PN0P_  (.CLK(clknet_leaf_261_clk_p2c),
    .RESET_B(net2103),
    .D(_01327_),
    .Q_N(_05640_),
    .Q(\shift_storage.storage[662] ));
 sg13g2_dfrbp_1 \shift_storage.storage[663]$_SDFFE_PN0P_  (.CLK(clknet_leaf_261_clk_p2c),
    .RESET_B(net2104),
    .D(_01328_),
    .Q_N(_05639_),
    .Q(\shift_storage.storage[663] ));
 sg13g2_dfrbp_1 \shift_storage.storage[664]$_SDFFE_PN0P_  (.CLK(clknet_leaf_263_clk_p2c),
    .RESET_B(net2105),
    .D(_01329_),
    .Q_N(_05638_),
    .Q(\shift_storage.storage[664] ));
 sg13g2_dfrbp_1 \shift_storage.storage[665]$_SDFFE_PN0P_  (.CLK(clknet_leaf_262_clk_p2c),
    .RESET_B(net2106),
    .D(_01330_),
    .Q_N(_05637_),
    .Q(\shift_storage.storage[665] ));
 sg13g2_dfrbp_1 \shift_storage.storage[666]$_SDFFE_PN0P_  (.CLK(clknet_leaf_263_clk_p2c),
    .RESET_B(net2107),
    .D(_01331_),
    .Q_N(_05636_),
    .Q(\shift_storage.storage[666] ));
 sg13g2_dfrbp_1 \shift_storage.storage[667]$_SDFFE_PN0P_  (.CLK(clknet_leaf_263_clk_p2c),
    .RESET_B(net2108),
    .D(_01332_),
    .Q_N(_05635_),
    .Q(\shift_storage.storage[667] ));
 sg13g2_dfrbp_1 \shift_storage.storage[668]$_SDFFE_PN0P_  (.CLK(clknet_leaf_264_clk_p2c),
    .RESET_B(net2109),
    .D(_01333_),
    .Q_N(_05634_),
    .Q(\shift_storage.storage[668] ));
 sg13g2_dfrbp_1 \shift_storage.storage[669]$_SDFFE_PN0P_  (.CLK(clknet_leaf_264_clk_p2c),
    .RESET_B(net2110),
    .D(_01334_),
    .Q_N(_05633_),
    .Q(\shift_storage.storage[669] ));
 sg13g2_dfrbp_1 \shift_storage.storage[66]$_SDFFE_PN0P_  (.CLK(clknet_leaf_39_clk_p2c),
    .RESET_B(net2111),
    .D(_01335_),
    .Q_N(_05632_),
    .Q(\shift_storage.storage[66] ));
 sg13g2_dfrbp_1 \shift_storage.storage[670]$_SDFFE_PN0P_  (.CLK(clknet_leaf_269_clk_p2c),
    .RESET_B(net2112),
    .D(_01336_),
    .Q_N(_05631_),
    .Q(\shift_storage.storage[670] ));
 sg13g2_dfrbp_1 \shift_storage.storage[671]$_SDFFE_PN0P_  (.CLK(clknet_leaf_269_clk_p2c),
    .RESET_B(net2113),
    .D(_01337_),
    .Q_N(_05630_),
    .Q(\shift_storage.storage[671] ));
 sg13g2_dfrbp_1 \shift_storage.storage[672]$_SDFFE_PN0P_  (.CLK(clknet_leaf_269_clk_p2c),
    .RESET_B(net2114),
    .D(_01338_),
    .Q_N(_05629_),
    .Q(\shift_storage.storage[672] ));
 sg13g2_dfrbp_1 \shift_storage.storage[673]$_SDFFE_PN0P_  (.CLK(clknet_leaf_275_clk_p2c),
    .RESET_B(net2115),
    .D(_01339_),
    .Q_N(_05628_),
    .Q(\shift_storage.storage[673] ));
 sg13g2_dfrbp_1 \shift_storage.storage[674]$_SDFFE_PN0P_  (.CLK(clknet_leaf_275_clk_p2c),
    .RESET_B(net2116),
    .D(_01340_),
    .Q_N(_05627_),
    .Q(\shift_storage.storage[674] ));
 sg13g2_dfrbp_1 \shift_storage.storage[675]$_SDFFE_PN0P_  (.CLK(clknet_leaf_275_clk_p2c),
    .RESET_B(net2117),
    .D(_01341_),
    .Q_N(_05626_),
    .Q(\shift_storage.storage[675] ));
 sg13g2_dfrbp_1 \shift_storage.storage[676]$_SDFFE_PN0P_  (.CLK(clknet_leaf_275_clk_p2c),
    .RESET_B(net2118),
    .D(_01342_),
    .Q_N(_05625_),
    .Q(\shift_storage.storage[676] ));
 sg13g2_dfrbp_1 \shift_storage.storage[677]$_SDFFE_PN0P_  (.CLK(clknet_leaf_276_clk_p2c),
    .RESET_B(net2119),
    .D(_01343_),
    .Q_N(_05624_),
    .Q(\shift_storage.storage[677] ));
 sg13g2_dfrbp_1 \shift_storage.storage[678]$_SDFFE_PN0P_  (.CLK(clknet_leaf_274_clk_p2c),
    .RESET_B(net2120),
    .D(_01344_),
    .Q_N(_05623_),
    .Q(\shift_storage.storage[678] ));
 sg13g2_dfrbp_1 \shift_storage.storage[679]$_SDFFE_PN0P_  (.CLK(clknet_leaf_274_clk_p2c),
    .RESET_B(net2121),
    .D(_01345_),
    .Q_N(_05622_),
    .Q(\shift_storage.storage[679] ));
 sg13g2_dfrbp_1 \shift_storage.storage[67]$_SDFFE_PN0P_  (.CLK(clknet_leaf_39_clk_p2c),
    .RESET_B(net2122),
    .D(_01346_),
    .Q_N(_05621_),
    .Q(\shift_storage.storage[67] ));
 sg13g2_dfrbp_1 \shift_storage.storage[680]$_SDFFE_PN0P_  (.CLK(clknet_leaf_274_clk_p2c),
    .RESET_B(net2123),
    .D(_01347_),
    .Q_N(_05620_),
    .Q(\shift_storage.storage[680] ));
 sg13g2_dfrbp_1 \shift_storage.storage[681]$_SDFFE_PN0P_  (.CLK(clknet_leaf_274_clk_p2c),
    .RESET_B(net2124),
    .D(_01348_),
    .Q_N(_05619_),
    .Q(\shift_storage.storage[681] ));
 sg13g2_dfrbp_1 \shift_storage.storage[682]$_SDFFE_PN0P_  (.CLK(clknet_leaf_270_clk_p2c),
    .RESET_B(net2125),
    .D(_01349_),
    .Q_N(_05618_),
    .Q(\shift_storage.storage[682] ));
 sg13g2_dfrbp_1 \shift_storage.storage[683]$_SDFFE_PN0P_  (.CLK(clknet_leaf_272_clk_p2c),
    .RESET_B(net2126),
    .D(_01350_),
    .Q_N(_05617_),
    .Q(\shift_storage.storage[683] ));
 sg13g2_dfrbp_1 \shift_storage.storage[684]$_SDFFE_PN0P_  (.CLK(clknet_leaf_272_clk_p2c),
    .RESET_B(net2127),
    .D(_01351_),
    .Q_N(_05616_),
    .Q(\shift_storage.storage[684] ));
 sg13g2_dfrbp_1 \shift_storage.storage[685]$_SDFFE_PN0P_  (.CLK(clknet_leaf_273_clk_p2c),
    .RESET_B(net2128),
    .D(_01352_),
    .Q_N(_05615_),
    .Q(\shift_storage.storage[685] ));
 sg13g2_dfrbp_1 \shift_storage.storage[686]$_SDFFE_PN0P_  (.CLK(clknet_leaf_273_clk_p2c),
    .RESET_B(net2129),
    .D(_01353_),
    .Q_N(_05614_),
    .Q(\shift_storage.storage[686] ));
 sg13g2_dfrbp_1 \shift_storage.storage[687]$_SDFFE_PN0P_  (.CLK(clknet_leaf_273_clk_p2c),
    .RESET_B(net2130),
    .D(_01354_),
    .Q_N(_05613_),
    .Q(\shift_storage.storage[687] ));
 sg13g2_dfrbp_1 \shift_storage.storage[688]$_SDFFE_PN0P_  (.CLK(clknet_leaf_274_clk_p2c),
    .RESET_B(net2131),
    .D(_01355_),
    .Q_N(_05612_),
    .Q(\shift_storage.storage[688] ));
 sg13g2_dfrbp_1 \shift_storage.storage[689]$_SDFFE_PN0P_  (.CLK(clknet_leaf_273_clk_p2c),
    .RESET_B(net2132),
    .D(_01356_),
    .Q_N(_05611_),
    .Q(\shift_storage.storage[689] ));
 sg13g2_dfrbp_1 \shift_storage.storage[68]$_SDFFE_PN0P_  (.CLK(clknet_leaf_98_clk_p2c),
    .RESET_B(net2133),
    .D(_01357_),
    .Q_N(_05610_),
    .Q(\shift_storage.storage[68] ));
 sg13g2_dfrbp_1 \shift_storage.storage[690]$_SDFFE_PN0P_  (.CLK(clknet_leaf_282_clk_p2c),
    .RESET_B(net2134),
    .D(_01358_),
    .Q_N(_05609_),
    .Q(\shift_storage.storage[690] ));
 sg13g2_dfrbp_1 \shift_storage.storage[691]$_SDFFE_PN0P_  (.CLK(clknet_leaf_282_clk_p2c),
    .RESET_B(net2135),
    .D(_01359_),
    .Q_N(_05608_),
    .Q(\shift_storage.storage[691] ));
 sg13g2_dfrbp_1 \shift_storage.storage[692]$_SDFFE_PN0P_  (.CLK(clknet_leaf_282_clk_p2c),
    .RESET_B(net2136),
    .D(_01360_),
    .Q_N(_05607_),
    .Q(\shift_storage.storage[692] ));
 sg13g2_dfrbp_1 \shift_storage.storage[693]$_SDFFE_PN0P_  (.CLK(clknet_leaf_283_clk_p2c),
    .RESET_B(net2137),
    .D(_01361_),
    .Q_N(_05606_),
    .Q(\shift_storage.storage[693] ));
 sg13g2_dfrbp_1 \shift_storage.storage[694]$_SDFFE_PN0P_  (.CLK(clknet_leaf_283_clk_p2c),
    .RESET_B(net2138),
    .D(_01362_),
    .Q_N(_05605_),
    .Q(\shift_storage.storage[694] ));
 sg13g2_dfrbp_1 \shift_storage.storage[695]$_SDFFE_PN0P_  (.CLK(clknet_leaf_283_clk_p2c),
    .RESET_B(net2139),
    .D(_01363_),
    .Q_N(_05604_),
    .Q(\shift_storage.storage[695] ));
 sg13g2_dfrbp_1 \shift_storage.storage[696]$_SDFFE_PN0P_  (.CLK(clknet_leaf_283_clk_p2c),
    .RESET_B(net2140),
    .D(_01364_),
    .Q_N(_05603_),
    .Q(\shift_storage.storage[696] ));
 sg13g2_dfrbp_1 \shift_storage.storage[697]$_SDFFE_PN0P_  (.CLK(clknet_leaf_283_clk_p2c),
    .RESET_B(net2141),
    .D(_01365_),
    .Q_N(_05602_),
    .Q(\shift_storage.storage[697] ));
 sg13g2_dfrbp_1 \shift_storage.storage[698]$_SDFFE_PN0P_  (.CLK(clknet_leaf_273_clk_p2c),
    .RESET_B(net2142),
    .D(_01366_),
    .Q_N(_05601_),
    .Q(\shift_storage.storage[698] ));
 sg13g2_dfrbp_1 \shift_storage.storage[699]$_SDFFE_PN0P_  (.CLK(clknet_leaf_272_clk_p2c),
    .RESET_B(net2143),
    .D(_01367_),
    .Q_N(_05600_),
    .Q(\shift_storage.storage[699] ));
 sg13g2_dfrbp_1 \shift_storage.storage[69]$_SDFFE_PN0P_  (.CLK(clknet_leaf_98_clk_p2c),
    .RESET_B(net2144),
    .D(_01368_),
    .Q_N(_05599_),
    .Q(\shift_storage.storage[69] ));
 sg13g2_dfrbp_1 \shift_storage.storage[6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_73_clk_p2c),
    .RESET_B(net2145),
    .D(_01369_),
    .Q_N(_05598_),
    .Q(\shift_storage.storage[6] ));
 sg13g2_dfrbp_1 \shift_storage.storage[700]$_SDFFE_PN0P_  (.CLK(clknet_leaf_272_clk_p2c),
    .RESET_B(net2146),
    .D(_01370_),
    .Q_N(_05597_),
    .Q(\shift_storage.storage[700] ));
 sg13g2_dfrbp_1 \shift_storage.storage[701]$_SDFFE_PN0P_  (.CLK(clknet_leaf_272_clk_p2c),
    .RESET_B(net2147),
    .D(_01371_),
    .Q_N(_05596_),
    .Q(\shift_storage.storage[701] ));
 sg13g2_dfrbp_1 \shift_storage.storage[702]$_SDFFE_PN0P_  (.CLK(clknet_leaf_272_clk_p2c),
    .RESET_B(net2148),
    .D(_01372_),
    .Q_N(_05595_),
    .Q(\shift_storage.storage[702] ));
 sg13g2_dfrbp_1 \shift_storage.storage[703]$_SDFFE_PN0P_  (.CLK(clknet_leaf_271_clk_p2c),
    .RESET_B(net2149),
    .D(_01373_),
    .Q_N(_05594_),
    .Q(\shift_storage.storage[703] ));
 sg13g2_dfrbp_1 \shift_storage.storage[704]$_SDFFE_PN0P_  (.CLK(clknet_leaf_271_clk_p2c),
    .RESET_B(net2150),
    .D(_01374_),
    .Q_N(_05593_),
    .Q(\shift_storage.storage[704] ));
 sg13g2_dfrbp_1 \shift_storage.storage[705]$_SDFFE_PN0P_  (.CLK(clknet_leaf_271_clk_p2c),
    .RESET_B(net2151),
    .D(_01375_),
    .Q_N(_05592_),
    .Q(\shift_storage.storage[705] ));
 sg13g2_dfrbp_1 \shift_storage.storage[706]$_SDFFE_PN0P_  (.CLK(clknet_leaf_271_clk_p2c),
    .RESET_B(net2152),
    .D(_01376_),
    .Q_N(_05591_),
    .Q(\shift_storage.storage[706] ));
 sg13g2_dfrbp_1 \shift_storage.storage[707]$_SDFFE_PN0P_  (.CLK(clknet_leaf_271_clk_p2c),
    .RESET_B(net2153),
    .D(_01377_),
    .Q_N(_05590_),
    .Q(\shift_storage.storage[707] ));
 sg13g2_dfrbp_1 \shift_storage.storage[708]$_SDFFE_PN0P_  (.CLK(clknet_leaf_271_clk_p2c),
    .RESET_B(net2154),
    .D(_01378_),
    .Q_N(_05589_),
    .Q(\shift_storage.storage[708] ));
 sg13g2_dfrbp_1 \shift_storage.storage[709]$_SDFFE_PN0P_  (.CLK(clknet_leaf_268_clk_p2c),
    .RESET_B(net2155),
    .D(_01379_),
    .Q_N(_05588_),
    .Q(\shift_storage.storage[709] ));
 sg13g2_dfrbp_1 \shift_storage.storage[70]$_SDFFE_PN0P_  (.CLK(clknet_leaf_98_clk_p2c),
    .RESET_B(net2156),
    .D(_01380_),
    .Q_N(_05587_),
    .Q(\shift_storage.storage[70] ));
 sg13g2_dfrbp_1 \shift_storage.storage[710]$_SDFFE_PN0P_  (.CLK(clknet_leaf_270_clk_p2c),
    .RESET_B(net2157),
    .D(_01381_),
    .Q_N(_05586_),
    .Q(\shift_storage.storage[710] ));
 sg13g2_dfrbp_1 \shift_storage.storage[711]$_SDFFE_PN0P_  (.CLK(clknet_leaf_270_clk_p2c),
    .RESET_B(net2158),
    .D(_01382_),
    .Q_N(_05585_),
    .Q(\shift_storage.storage[711] ));
 sg13g2_dfrbp_1 \shift_storage.storage[712]$_SDFFE_PN0P_  (.CLK(clknet_leaf_270_clk_p2c),
    .RESET_B(net2159),
    .D(_01383_),
    .Q_N(_05584_),
    .Q(\shift_storage.storage[712] ));
 sg13g2_dfrbp_1 \shift_storage.storage[713]$_SDFFE_PN0P_  (.CLK(clknet_leaf_270_clk_p2c),
    .RESET_B(net2160),
    .D(_01384_),
    .Q_N(_05583_),
    .Q(\shift_storage.storage[713] ));
 sg13g2_dfrbp_1 \shift_storage.storage[714]$_SDFFE_PN0P_  (.CLK(clknet_leaf_269_clk_p2c),
    .RESET_B(net2161),
    .D(_01385_),
    .Q_N(_05582_),
    .Q(\shift_storage.storage[714] ));
 sg13g2_dfrbp_1 \shift_storage.storage[715]$_SDFFE_PN0P_  (.CLK(clknet_leaf_269_clk_p2c),
    .RESET_B(net2162),
    .D(_01386_),
    .Q_N(_05581_),
    .Q(\shift_storage.storage[715] ));
 sg13g2_dfrbp_1 \shift_storage.storage[716]$_SDFFE_PN0P_  (.CLK(clknet_leaf_269_clk_p2c),
    .RESET_B(net2163),
    .D(_01387_),
    .Q_N(_05580_),
    .Q(\shift_storage.storage[716] ));
 sg13g2_dfrbp_1 \shift_storage.storage[717]$_SDFFE_PN0P_  (.CLK(clknet_leaf_269_clk_p2c),
    .RESET_B(net2164),
    .D(_01388_),
    .Q_N(_05579_),
    .Q(\shift_storage.storage[717] ));
 sg13g2_dfrbp_1 \shift_storage.storage[718]$_SDFFE_PN0P_  (.CLK(clknet_leaf_268_clk_p2c),
    .RESET_B(net2165),
    .D(_01389_),
    .Q_N(_05578_),
    .Q(\shift_storage.storage[718] ));
 sg13g2_dfrbp_1 \shift_storage.storage[719]$_SDFFE_PN0P_  (.CLK(clknet_leaf_268_clk_p2c),
    .RESET_B(net2166),
    .D(_01390_),
    .Q_N(_05577_),
    .Q(\shift_storage.storage[719] ));
 sg13g2_dfrbp_1 \shift_storage.storage[71]$_SDFFE_PN0P_  (.CLK(clknet_leaf_98_clk_p2c),
    .RESET_B(net2167),
    .D(_01391_),
    .Q_N(_05576_),
    .Q(\shift_storage.storage[71] ));
 sg13g2_dfrbp_1 \shift_storage.storage[720]$_SDFFE_PN0P_  (.CLK(clknet_leaf_267_clk_p2c),
    .RESET_B(net2168),
    .D(_01392_),
    .Q_N(_05575_),
    .Q(\shift_storage.storage[720] ));
 sg13g2_dfrbp_1 \shift_storage.storage[721]$_SDFFE_PN0P_  (.CLK(clknet_leaf_267_clk_p2c),
    .RESET_B(net2169),
    .D(_01393_),
    .Q_N(_05574_),
    .Q(\shift_storage.storage[721] ));
 sg13g2_dfrbp_1 \shift_storage.storage[722]$_SDFFE_PN0P_  (.CLK(clknet_leaf_268_clk_p2c),
    .RESET_B(net2170),
    .D(_01394_),
    .Q_N(_05573_),
    .Q(\shift_storage.storage[722] ));
 sg13g2_dfrbp_1 \shift_storage.storage[723]$_SDFFE_PN0P_  (.CLK(clknet_leaf_268_clk_p2c),
    .RESET_B(net2171),
    .D(_01395_),
    .Q_N(_05572_),
    .Q(\shift_storage.storage[723] ));
 sg13g2_dfrbp_1 \shift_storage.storage[724]$_SDFFE_PN0P_  (.CLK(clknet_leaf_267_clk_p2c),
    .RESET_B(net2172),
    .D(_01396_),
    .Q_N(_05571_),
    .Q(\shift_storage.storage[724] ));
 sg13g2_dfrbp_1 \shift_storage.storage[725]$_SDFFE_PN0P_  (.CLK(clknet_leaf_267_clk_p2c),
    .RESET_B(net2173),
    .D(_01397_),
    .Q_N(_05570_),
    .Q(\shift_storage.storage[725] ));
 sg13g2_dfrbp_1 \shift_storage.storage[726]$_SDFFE_PN0P_  (.CLK(clknet_leaf_267_clk_p2c),
    .RESET_B(net2174),
    .D(_01398_),
    .Q_N(_05569_),
    .Q(\shift_storage.storage[726] ));
 sg13g2_dfrbp_1 \shift_storage.storage[727]$_SDFFE_PN0P_  (.CLK(clknet_leaf_266_clk_p2c),
    .RESET_B(net2175),
    .D(_01399_),
    .Q_N(_05568_),
    .Q(\shift_storage.storage[727] ));
 sg13g2_dfrbp_1 \shift_storage.storage[728]$_SDFFE_PN0P_  (.CLK(clknet_leaf_266_clk_p2c),
    .RESET_B(net2176),
    .D(_01400_),
    .Q_N(_05567_),
    .Q(\shift_storage.storage[728] ));
 sg13g2_dfrbp_1 \shift_storage.storage[729]$_SDFFE_PN0P_  (.CLK(clknet_leaf_220_clk_p2c),
    .RESET_B(net2177),
    .D(_01401_),
    .Q_N(_05566_),
    .Q(\shift_storage.storage[729] ));
 sg13g2_dfrbp_1 \shift_storage.storage[72]$_SDFFE_PN0P_  (.CLK(clknet_leaf_97_clk_p2c),
    .RESET_B(net2178),
    .D(_01402_),
    .Q_N(_05565_),
    .Q(\shift_storage.storage[72] ));
 sg13g2_dfrbp_1 \shift_storage.storage[730]$_SDFFE_PN0P_  (.CLK(clknet_leaf_220_clk_p2c),
    .RESET_B(net2179),
    .D(_01403_),
    .Q_N(_05564_),
    .Q(\shift_storage.storage[730] ));
 sg13g2_dfrbp_1 \shift_storage.storage[731]$_SDFFE_PN0P_  (.CLK(clknet_leaf_266_clk_p2c),
    .RESET_B(net2180),
    .D(_01404_),
    .Q_N(_05563_),
    .Q(\shift_storage.storage[731] ));
 sg13g2_dfrbp_1 \shift_storage.storage[732]$_SDFFE_PN0P_  (.CLK(clknet_leaf_267_clk_p2c),
    .RESET_B(net2181),
    .D(_01405_),
    .Q_N(_05562_),
    .Q(\shift_storage.storage[732] ));
 sg13g2_dfrbp_1 \shift_storage.storage[733]$_SDFFE_PN0P_  (.CLK(clknet_leaf_265_clk_p2c),
    .RESET_B(net2182),
    .D(_01406_),
    .Q_N(_05561_),
    .Q(\shift_storage.storage[733] ));
 sg13g2_dfrbp_1 \shift_storage.storage[734]$_SDFFE_PN0P_  (.CLK(clknet_leaf_265_clk_p2c),
    .RESET_B(net2183),
    .D(_01407_),
    .Q_N(_05560_),
    .Q(\shift_storage.storage[734] ));
 sg13g2_dfrbp_1 \shift_storage.storage[735]$_SDFFE_PN0P_  (.CLK(clknet_leaf_265_clk_p2c),
    .RESET_B(net2184),
    .D(_01408_),
    .Q_N(_05559_),
    .Q(\shift_storage.storage[735] ));
 sg13g2_dfrbp_1 \shift_storage.storage[736]$_SDFFE_PN0P_  (.CLK(clknet_leaf_264_clk_p2c),
    .RESET_B(net2185),
    .D(_01409_),
    .Q_N(_05558_),
    .Q(\shift_storage.storage[736] ));
 sg13g2_dfrbp_1 \shift_storage.storage[737]$_SDFFE_PN0P_  (.CLK(clknet_leaf_264_clk_p2c),
    .RESET_B(net2186),
    .D(_01410_),
    .Q_N(_05557_),
    .Q(\shift_storage.storage[737] ));
 sg13g2_dfrbp_1 \shift_storage.storage[738]$_SDFFE_PN0P_  (.CLK(clknet_leaf_264_clk_p2c),
    .RESET_B(net2187),
    .D(_01411_),
    .Q_N(_05556_),
    .Q(\shift_storage.storage[738] ));
 sg13g2_dfrbp_1 \shift_storage.storage[739]$_SDFFE_PN0P_  (.CLK(clknet_leaf_264_clk_p2c),
    .RESET_B(net2188),
    .D(_01412_),
    .Q_N(_05555_),
    .Q(\shift_storage.storage[739] ));
 sg13g2_dfrbp_1 \shift_storage.storage[73]$_SDFFE_PN0P_  (.CLK(clknet_leaf_97_clk_p2c),
    .RESET_B(net2189),
    .D(_01413_),
    .Q_N(_05554_),
    .Q(\shift_storage.storage[73] ));
 sg13g2_dfrbp_1 \shift_storage.storage[740]$_SDFFE_PN0P_  (.CLK(clknet_leaf_265_clk_p2c),
    .RESET_B(net2190),
    .D(_01414_),
    .Q_N(_05553_),
    .Q(\shift_storage.storage[740] ));
 sg13g2_dfrbp_1 \shift_storage.storage[741]$_SDFFE_PN0P_  (.CLK(clknet_leaf_262_clk_p2c),
    .RESET_B(net2191),
    .D(_01415_),
    .Q_N(_05552_),
    .Q(\shift_storage.storage[741] ));
 sg13g2_dfrbp_1 \shift_storage.storage[742]$_SDFFE_PN0P_  (.CLK(clknet_leaf_262_clk_p2c),
    .RESET_B(net2192),
    .D(_01416_),
    .Q_N(_05551_),
    .Q(\shift_storage.storage[742] ));
 sg13g2_dfrbp_1 \shift_storage.storage[743]$_SDFFE_PN0P_  (.CLK(clknet_leaf_262_clk_p2c),
    .RESET_B(net2193),
    .D(_01417_),
    .Q_N(_05550_),
    .Q(\shift_storage.storage[743] ));
 sg13g2_dfrbp_1 \shift_storage.storage[744]$_SDFFE_PN0P_  (.CLK(clknet_leaf_262_clk_p2c),
    .RESET_B(net2194),
    .D(_01418_),
    .Q_N(_05549_),
    .Q(\shift_storage.storage[744] ));
 sg13g2_dfrbp_1 \shift_storage.storage[745]$_SDFFE_PN0P_  (.CLK(clknet_leaf_225_clk_p2c),
    .RESET_B(net2195),
    .D(_01419_),
    .Q_N(_05548_),
    .Q(\shift_storage.storage[745] ));
 sg13g2_dfrbp_1 \shift_storage.storage[746]$_SDFFE_PN0P_  (.CLK(clknet_leaf_225_clk_p2c),
    .RESET_B(net2196),
    .D(_01420_),
    .Q_N(_05547_),
    .Q(\shift_storage.storage[746] ));
 sg13g2_dfrbp_1 \shift_storage.storage[747]$_SDFFE_PN0P_  (.CLK(clknet_leaf_225_clk_p2c),
    .RESET_B(net2197),
    .D(_01421_),
    .Q_N(_05546_),
    .Q(\shift_storage.storage[747] ));
 sg13g2_dfrbp_1 \shift_storage.storage[748]$_SDFFE_PN0P_  (.CLK(clknet_leaf_225_clk_p2c),
    .RESET_B(net2198),
    .D(_01422_),
    .Q_N(_05545_),
    .Q(\shift_storage.storage[748] ));
 sg13g2_dfrbp_1 \shift_storage.storage[749]$_SDFFE_PN0P_  (.CLK(clknet_leaf_225_clk_p2c),
    .RESET_B(net2199),
    .D(_01423_),
    .Q_N(_05544_),
    .Q(\shift_storage.storage[749] ));
 sg13g2_dfrbp_1 \shift_storage.storage[74]$_SDFFE_PN0P_  (.CLK(clknet_leaf_98_clk_p2c),
    .RESET_B(net2200),
    .D(_01424_),
    .Q_N(_05543_),
    .Q(\shift_storage.storage[74] ));
 sg13g2_dfrbp_1 \shift_storage.storage[750]$_SDFFE_PN0P_  (.CLK(clknet_leaf_226_clk_p2c),
    .RESET_B(net2201),
    .D(_01425_),
    .Q_N(_05542_),
    .Q(\shift_storage.storage[750] ));
 sg13g2_dfrbp_1 \shift_storage.storage[751]$_SDFFE_PN0P_  (.CLK(clknet_leaf_224_clk_p2c),
    .RESET_B(net2202),
    .D(_01426_),
    .Q_N(_05541_),
    .Q(\shift_storage.storage[751] ));
 sg13g2_dfrbp_1 \shift_storage.storage[752]$_SDFFE_PN0P_  (.CLK(clknet_leaf_224_clk_p2c),
    .RESET_B(net2203),
    .D(_01427_),
    .Q_N(_05540_),
    .Q(\shift_storage.storage[752] ));
 sg13g2_dfrbp_1 \shift_storage.storage[753]$_SDFFE_PN0P_  (.CLK(clknet_leaf_224_clk_p2c),
    .RESET_B(net2204),
    .D(_01428_),
    .Q_N(_05539_),
    .Q(\shift_storage.storage[753] ));
 sg13g2_dfrbp_1 \shift_storage.storage[754]$_SDFFE_PN0P_  (.CLK(clknet_leaf_222_clk_p2c),
    .RESET_B(net2205),
    .D(_01429_),
    .Q_N(_05538_),
    .Q(\shift_storage.storage[754] ));
 sg13g2_dfrbp_1 \shift_storage.storage[755]$_SDFFE_PN0P_  (.CLK(clknet_leaf_222_clk_p2c),
    .RESET_B(net2206),
    .D(_01430_),
    .Q_N(_05537_),
    .Q(\shift_storage.storage[755] ));
 sg13g2_dfrbp_1 \shift_storage.storage[756]$_SDFFE_PN0P_  (.CLK(clknet_leaf_222_clk_p2c),
    .RESET_B(net2207),
    .D(_01431_),
    .Q_N(_05536_),
    .Q(\shift_storage.storage[756] ));
 sg13g2_dfrbp_1 \shift_storage.storage[757]$_SDFFE_PN0P_  (.CLK(clknet_leaf_222_clk_p2c),
    .RESET_B(net2208),
    .D(_01432_),
    .Q_N(_05535_),
    .Q(\shift_storage.storage[757] ));
 sg13g2_dfrbp_1 \shift_storage.storage[758]$_SDFFE_PN0P_  (.CLK(clknet_leaf_221_clk_p2c),
    .RESET_B(net2209),
    .D(_01433_),
    .Q_N(_05534_),
    .Q(\shift_storage.storage[758] ));
 sg13g2_dfrbp_1 \shift_storage.storage[759]$_SDFFE_PN0P_  (.CLK(clknet_leaf_222_clk_p2c),
    .RESET_B(net2210),
    .D(_01434_),
    .Q_N(_05533_),
    .Q(\shift_storage.storage[759] ));
 sg13g2_dfrbp_1 \shift_storage.storage[75]$_SDFFE_PN0P_  (.CLK(clknet_leaf_99_clk_p2c),
    .RESET_B(net2211),
    .D(_01435_),
    .Q_N(_05532_),
    .Q(\shift_storage.storage[75] ));
 sg13g2_dfrbp_1 \shift_storage.storage[760]$_SDFFE_PN0P_  (.CLK(clknet_leaf_265_clk_p2c),
    .RESET_B(net2212),
    .D(_01436_),
    .Q_N(_05531_),
    .Q(\shift_storage.storage[760] ));
 sg13g2_dfrbp_1 \shift_storage.storage[761]$_SDFFE_PN0P_  (.CLK(clknet_leaf_265_clk_p2c),
    .RESET_B(net2213),
    .D(_01437_),
    .Q_N(_05530_),
    .Q(\shift_storage.storage[761] ));
 sg13g2_dfrbp_1 \shift_storage.storage[762]$_SDFFE_PN0P_  (.CLK(clknet_leaf_266_clk_p2c),
    .RESET_B(net2214),
    .D(_01438_),
    .Q_N(_05529_),
    .Q(\shift_storage.storage[762] ));
 sg13g2_dfrbp_1 \shift_storage.storage[763]$_SDFFE_PN0P_  (.CLK(clknet_leaf_266_clk_p2c),
    .RESET_B(net2215),
    .D(_01439_),
    .Q_N(_05528_),
    .Q(\shift_storage.storage[763] ));
 sg13g2_dfrbp_1 \shift_storage.storage[764]$_SDFFE_PN0P_  (.CLK(clknet_leaf_220_clk_p2c),
    .RESET_B(net2216),
    .D(_01440_),
    .Q_N(_05527_),
    .Q(\shift_storage.storage[764] ));
 sg13g2_dfrbp_1 \shift_storage.storage[765]$_SDFFE_PN0P_  (.CLK(clknet_leaf_221_clk_p2c),
    .RESET_B(net2217),
    .D(_01441_),
    .Q_N(_05526_),
    .Q(\shift_storage.storage[765] ));
 sg13g2_dfrbp_1 \shift_storage.storage[766]$_SDFFE_PN0P_  (.CLK(clknet_leaf_221_clk_p2c),
    .RESET_B(net2218),
    .D(_01442_),
    .Q_N(_05525_),
    .Q(\shift_storage.storage[766] ));
 sg13g2_dfrbp_1 \shift_storage.storage[767]$_SDFFE_PN0P_  (.CLK(clknet_leaf_221_clk_p2c),
    .RESET_B(net2219),
    .D(_01443_),
    .Q_N(_05524_),
    .Q(\shift_storage.storage[767] ));
 sg13g2_dfrbp_1 \shift_storage.storage[768]$_SDFFE_PN0P_  (.CLK(clknet_leaf_221_clk_p2c),
    .RESET_B(net2220),
    .D(_01444_),
    .Q_N(_05523_),
    .Q(\shift_storage.storage[768] ));
 sg13g2_dfrbp_1 \shift_storage.storage[769]$_SDFFE_PN0P_  (.CLK(clknet_leaf_221_clk_p2c),
    .RESET_B(net2221),
    .D(_01445_),
    .Q_N(_05522_),
    .Q(\shift_storage.storage[769] ));
 sg13g2_dfrbp_1 \shift_storage.storage[76]$_SDFFE_PN0P_  (.CLK(clknet_leaf_100_clk_p2c),
    .RESET_B(net2222),
    .D(_01446_),
    .Q_N(_05521_),
    .Q(\shift_storage.storage[76] ));
 sg13g2_dfrbp_1 \shift_storage.storage[770]$_SDFFE_PN0P_  (.CLK(clknet_leaf_223_clk_p2c),
    .RESET_B(net2223),
    .D(_01447_),
    .Q_N(_05520_),
    .Q(\shift_storage.storage[770] ));
 sg13g2_dfrbp_1 \shift_storage.storage[771]$_SDFFE_PN0P_  (.CLK(clknet_leaf_223_clk_p2c),
    .RESET_B(net2224),
    .D(_01448_),
    .Q_N(_05519_),
    .Q(\shift_storage.storage[771] ));
 sg13g2_dfrbp_1 \shift_storage.storage[772]$_SDFFE_PN0P_  (.CLK(clknet_leaf_220_clk_p2c),
    .RESET_B(net2225),
    .D(_01449_),
    .Q_N(_05518_),
    .Q(\shift_storage.storage[772] ));
 sg13g2_dfrbp_1 \shift_storage.storage[773]$_SDFFE_PN0P_  (.CLK(clknet_leaf_220_clk_p2c),
    .RESET_B(net2226),
    .D(_01450_),
    .Q_N(_05517_),
    .Q(\shift_storage.storage[773] ));
 sg13g2_dfrbp_1 \shift_storage.storage[774]$_SDFFE_PN0P_  (.CLK(clknet_leaf_219_clk_p2c),
    .RESET_B(net2227),
    .D(_01451_),
    .Q_N(_05516_),
    .Q(\shift_storage.storage[774] ));
 sg13g2_dfrbp_1 \shift_storage.storage[775]$_SDFFE_PN0P_  (.CLK(clknet_leaf_219_clk_p2c),
    .RESET_B(net2228),
    .D(_01452_),
    .Q_N(_05515_),
    .Q(\shift_storage.storage[775] ));
 sg13g2_dfrbp_1 \shift_storage.storage[776]$_SDFFE_PN0P_  (.CLK(clknet_leaf_219_clk_p2c),
    .RESET_B(net2229),
    .D(_01453_),
    .Q_N(_05514_),
    .Q(\shift_storage.storage[776] ));
 sg13g2_dfrbp_1 \shift_storage.storage[777]$_SDFFE_PN0P_  (.CLK(clknet_leaf_215_clk_p2c),
    .RESET_B(net2230),
    .D(_01454_),
    .Q_N(_05513_),
    .Q(\shift_storage.storage[777] ));
 sg13g2_dfrbp_1 \shift_storage.storage[778]$_SDFFE_PN0P_  (.CLK(clknet_leaf_215_clk_p2c),
    .RESET_B(net2231),
    .D(_01455_),
    .Q_N(_05512_),
    .Q(\shift_storage.storage[778] ));
 sg13g2_dfrbp_1 \shift_storage.storage[779]$_SDFFE_PN0P_  (.CLK(clknet_leaf_215_clk_p2c),
    .RESET_B(net2232),
    .D(_01456_),
    .Q_N(_05511_),
    .Q(\shift_storage.storage[779] ));
 sg13g2_dfrbp_1 \shift_storage.storage[77]$_SDFFE_PN0P_  (.CLK(clknet_leaf_100_clk_p2c),
    .RESET_B(net2233),
    .D(_01457_),
    .Q_N(_05510_),
    .Q(\shift_storage.storage[77] ));
 sg13g2_dfrbp_1 \shift_storage.storage[780]$_SDFFE_PN0P_  (.CLK(clknet_leaf_215_clk_p2c),
    .RESET_B(net2234),
    .D(_01458_),
    .Q_N(_05509_),
    .Q(\shift_storage.storage[780] ));
 sg13g2_dfrbp_1 \shift_storage.storage[781]$_SDFFE_PN0P_  (.CLK(clknet_leaf_215_clk_p2c),
    .RESET_B(net2235),
    .D(_01459_),
    .Q_N(_05508_),
    .Q(\shift_storage.storage[781] ));
 sg13g2_dfrbp_1 \shift_storage.storage[782]$_SDFFE_PN0P_  (.CLK(clknet_leaf_229_clk_p2c),
    .RESET_B(net2236),
    .D(_01460_),
    .Q_N(_05507_),
    .Q(\shift_storage.storage[782] ));
 sg13g2_dfrbp_1 \shift_storage.storage[783]$_SDFFE_PN0P_  (.CLK(clknet_leaf_215_clk_p2c),
    .RESET_B(net2237),
    .D(_01461_),
    .Q_N(_05506_),
    .Q(\shift_storage.storage[783] ));
 sg13g2_dfrbp_1 \shift_storage.storage[784]$_SDFFE_PN0P_  (.CLK(clknet_leaf_229_clk_p2c),
    .RESET_B(net2238),
    .D(_01462_),
    .Q_N(_05505_),
    .Q(\shift_storage.storage[784] ));
 sg13g2_dfrbp_1 \shift_storage.storage[785]$_SDFFE_PN0P_  (.CLK(clknet_leaf_229_clk_p2c),
    .RESET_B(net2239),
    .D(_01463_),
    .Q_N(_05504_),
    .Q(\shift_storage.storage[785] ));
 sg13g2_dfrbp_1 \shift_storage.storage[786]$_SDFFE_PN0P_  (.CLK(clknet_leaf_215_clk_p2c),
    .RESET_B(net2240),
    .D(_01464_),
    .Q_N(_05503_),
    .Q(\shift_storage.storage[786] ));
 sg13g2_dfrbp_1 \shift_storage.storage[787]$_SDFFE_PN0P_  (.CLK(clknet_leaf_223_clk_p2c),
    .RESET_B(net2241),
    .D(_01465_),
    .Q_N(_05502_),
    .Q(\shift_storage.storage[787] ));
 sg13g2_dfrbp_1 \shift_storage.storage[788]$_SDFFE_PN0P_  (.CLK(clknet_leaf_223_clk_p2c),
    .RESET_B(net2242),
    .D(_01466_),
    .Q_N(_05501_),
    .Q(\shift_storage.storage[788] ));
 sg13g2_dfrbp_1 \shift_storage.storage[789]$_SDFFE_PN0P_  (.CLK(clknet_leaf_223_clk_p2c),
    .RESET_B(net2243),
    .D(_01467_),
    .Q_N(_05500_),
    .Q(\shift_storage.storage[789] ));
 sg13g2_dfrbp_1 \shift_storage.storage[78]$_SDFFE_PN0P_  (.CLK(clknet_leaf_97_clk_p2c),
    .RESET_B(net2244),
    .D(_01468_),
    .Q_N(_05499_),
    .Q(\shift_storage.storage[78] ));
 sg13g2_dfrbp_1 \shift_storage.storage[790]$_SDFFE_PN0P_  (.CLK(clknet_leaf_223_clk_p2c),
    .RESET_B(net2245),
    .D(_01469_),
    .Q_N(_05498_),
    .Q(\shift_storage.storage[790] ));
 sg13g2_dfrbp_1 \shift_storage.storage[791]$_SDFFE_PN0P_  (.CLK(clknet_leaf_224_clk_p2c),
    .RESET_B(net2246),
    .D(_01470_),
    .Q_N(_05497_),
    .Q(\shift_storage.storage[791] ));
 sg13g2_dfrbp_1 \shift_storage.storage[792]$_SDFFE_PN0P_  (.CLK(clknet_leaf_224_clk_p2c),
    .RESET_B(net2247),
    .D(_01471_),
    .Q_N(_05496_),
    .Q(\shift_storage.storage[792] ));
 sg13g2_dfrbp_1 \shift_storage.storage[793]$_SDFFE_PN0P_  (.CLK(clknet_leaf_224_clk_p2c),
    .RESET_B(net2248),
    .D(_01472_),
    .Q_N(_05495_),
    .Q(\shift_storage.storage[793] ));
 sg13g2_dfrbp_1 \shift_storage.storage[794]$_SDFFE_PN0P_  (.CLK(clknet_leaf_228_clk_p2c),
    .RESET_B(net2249),
    .D(_01473_),
    .Q_N(_05494_),
    .Q(\shift_storage.storage[794] ));
 sg13g2_dfrbp_1 \shift_storage.storage[795]$_SDFFE_PN0P_  (.CLK(clknet_leaf_228_clk_p2c),
    .RESET_B(net2250),
    .D(_01474_),
    .Q_N(_05493_),
    .Q(\shift_storage.storage[795] ));
 sg13g2_dfrbp_1 \shift_storage.storage[796]$_SDFFE_PN0P_  (.CLK(clknet_leaf_228_clk_p2c),
    .RESET_B(net2251),
    .D(_01475_),
    .Q_N(_05492_),
    .Q(\shift_storage.storage[796] ));
 sg13g2_dfrbp_1 \shift_storage.storage[797]$_SDFFE_PN0P_  (.CLK(clknet_leaf_227_clk_p2c),
    .RESET_B(net2252),
    .D(_01476_),
    .Q_N(_05491_),
    .Q(\shift_storage.storage[797] ));
 sg13g2_dfrbp_1 \shift_storage.storage[798]$_SDFFE_PN0P_  (.CLK(clknet_leaf_227_clk_p2c),
    .RESET_B(net2253),
    .D(_01477_),
    .Q_N(_05490_),
    .Q(\shift_storage.storage[798] ));
 sg13g2_dfrbp_1 \shift_storage.storage[799]$_SDFFE_PN0P_  (.CLK(clknet_leaf_227_clk_p2c),
    .RESET_B(net2254),
    .D(_01478_),
    .Q_N(_05489_),
    .Q(\shift_storage.storage[799] ));
 sg13g2_dfrbp_1 \shift_storage.storage[79]$_SDFFE_PN0P_  (.CLK(clknet_leaf_94_clk_p2c),
    .RESET_B(net2255),
    .D(_01479_),
    .Q_N(_05488_),
    .Q(\shift_storage.storage[79] ));
 sg13g2_dfrbp_1 \shift_storage.storage[7]$_SDFFE_PN0P_  (.CLK(clknet_leaf_73_clk_p2c),
    .RESET_B(net2256),
    .D(_01480_),
    .Q_N(_05487_),
    .Q(\shift_storage.storage[7] ));
 sg13g2_dfrbp_1 \shift_storage.storage[800]$_SDFFE_PN0P_  (.CLK(clknet_leaf_226_clk_p2c),
    .RESET_B(net2257),
    .D(_01481_),
    .Q_N(_05486_),
    .Q(\shift_storage.storage[800] ));
 sg13g2_dfrbp_1 \shift_storage.storage[801]$_SDFFE_PN0P_  (.CLK(clknet_leaf_226_clk_p2c),
    .RESET_B(net2258),
    .D(_01482_),
    .Q_N(_05485_),
    .Q(\shift_storage.storage[801] ));
 sg13g2_dfrbp_1 \shift_storage.storage[802]$_SDFFE_PN0P_  (.CLK(clknet_leaf_226_clk_p2c),
    .RESET_B(net2259),
    .D(_01483_),
    .Q_N(_05484_),
    .Q(\shift_storage.storage[802] ));
 sg13g2_dfrbp_1 \shift_storage.storage[803]$_SDFFE_PN0P_  (.CLK(clknet_leaf_226_clk_p2c),
    .RESET_B(net2260),
    .D(_01484_),
    .Q_N(_05483_),
    .Q(\shift_storage.storage[803] ));
 sg13g2_dfrbp_1 \shift_storage.storage[804]$_SDFFE_PN0P_  (.CLK(clknet_leaf_226_clk_p2c),
    .RESET_B(net2261),
    .D(_01485_),
    .Q_N(_05482_),
    .Q(\shift_storage.storage[804] ));
 sg13g2_dfrbp_1 \shift_storage.storage[805]$_SDFFE_PN0P_  (.CLK(clknet_leaf_261_clk_p2c),
    .RESET_B(net2262),
    .D(_01486_),
    .Q_N(_05481_),
    .Q(\shift_storage.storage[805] ));
 sg13g2_dfrbp_1 \shift_storage.storage[806]$_SDFFE_PN0P_  (.CLK(clknet_leaf_261_clk_p2c),
    .RESET_B(net2263),
    .D(_01487_),
    .Q_N(_05480_),
    .Q(\shift_storage.storage[806] ));
 sg13g2_dfrbp_1 \shift_storage.storage[807]$_SDFFE_PN0P_  (.CLK(clknet_leaf_261_clk_p2c),
    .RESET_B(net2264),
    .D(_01488_),
    .Q_N(_05479_),
    .Q(\shift_storage.storage[807] ));
 sg13g2_dfrbp_1 \shift_storage.storage[808]$_SDFFE_PN0P_  (.CLK(clknet_leaf_260_clk_p2c),
    .RESET_B(net2265),
    .D(_01489_),
    .Q_N(_05478_),
    .Q(\shift_storage.storage[808] ));
 sg13g2_dfrbp_1 \shift_storage.storage[809]$_SDFFE_PN0P_  (.CLK(clknet_leaf_259_clk_p2c),
    .RESET_B(net2266),
    .D(_01490_),
    .Q_N(_05477_),
    .Q(\shift_storage.storage[809] ));
 sg13g2_dfrbp_1 \shift_storage.storage[80]$_SDFFE_PN0P_  (.CLK(clknet_leaf_94_clk_p2c),
    .RESET_B(net2267),
    .D(_01491_),
    .Q_N(_05476_),
    .Q(\shift_storage.storage[80] ));
 sg13g2_dfrbp_1 \shift_storage.storage[810]$_SDFFE_PN0P_  (.CLK(clknet_leaf_259_clk_p2c),
    .RESET_B(net2268),
    .D(_01492_),
    .Q_N(_05475_),
    .Q(\shift_storage.storage[810] ));
 sg13g2_dfrbp_1 \shift_storage.storage[811]$_SDFFE_PN0P_  (.CLK(clknet_leaf_260_clk_p2c),
    .RESET_B(net2269),
    .D(_01493_),
    .Q_N(_05474_),
    .Q(\shift_storage.storage[811] ));
 sg13g2_dfrbp_1 \shift_storage.storage[812]$_SDFFE_PN0P_  (.CLK(clknet_leaf_260_clk_p2c),
    .RESET_B(net2270),
    .D(_01494_),
    .Q_N(_05473_),
    .Q(\shift_storage.storage[812] ));
 sg13g2_dfrbp_1 \shift_storage.storage[813]$_SDFFE_PN0P_  (.CLK(clknet_leaf_249_clk_p2c),
    .RESET_B(net2271),
    .D(_01495_),
    .Q_N(_05472_),
    .Q(\shift_storage.storage[813] ));
 sg13g2_dfrbp_1 \shift_storage.storage[814]$_SDFFE_PN0P_  (.CLK(clknet_leaf_260_clk_p2c),
    .RESET_B(net2272),
    .D(_01496_),
    .Q_N(_05471_),
    .Q(\shift_storage.storage[814] ));
 sg13g2_dfrbp_1 \shift_storage.storage[815]$_SDFFE_PN0P_  (.CLK(clknet_leaf_260_clk_p2c),
    .RESET_B(net2273),
    .D(_01497_),
    .Q_N(_05470_),
    .Q(\shift_storage.storage[815] ));
 sg13g2_dfrbp_1 \shift_storage.storage[816]$_SDFFE_PN0P_  (.CLK(clknet_leaf_226_clk_p2c),
    .RESET_B(net2274),
    .D(_01498_),
    .Q_N(_05469_),
    .Q(\shift_storage.storage[816] ));
 sg13g2_dfrbp_1 \shift_storage.storage[817]$_SDFFE_PN0P_  (.CLK(clknet_leaf_237_clk_p2c),
    .RESET_B(net2275),
    .D(_01499_),
    .Q_N(_05468_),
    .Q(\shift_storage.storage[817] ));
 sg13g2_dfrbp_1 \shift_storage.storage[818]$_SDFFE_PN0P_  (.CLK(clknet_leaf_237_clk_p2c),
    .RESET_B(net2276),
    .D(_01500_),
    .Q_N(_05467_),
    .Q(\shift_storage.storage[818] ));
 sg13g2_dfrbp_1 \shift_storage.storage[819]$_SDFFE_PN0P_  (.CLK(clknet_leaf_238_clk_p2c),
    .RESET_B(net2277),
    .D(_01501_),
    .Q_N(_05466_),
    .Q(\shift_storage.storage[819] ));
 sg13g2_dfrbp_1 \shift_storage.storage[81]$_SDFFE_PN0P_  (.CLK(clknet_leaf_96_clk_p2c),
    .RESET_B(net2278),
    .D(_01502_),
    .Q_N(_05465_),
    .Q(\shift_storage.storage[81] ));
 sg13g2_dfrbp_1 \shift_storage.storage[820]$_SDFFE_PN0P_  (.CLK(clknet_leaf_238_clk_p2c),
    .RESET_B(net2279),
    .D(_01503_),
    .Q_N(_05464_),
    .Q(\shift_storage.storage[820] ));
 sg13g2_dfrbp_1 \shift_storage.storage[821]$_SDFFE_PN0P_  (.CLK(clknet_leaf_238_clk_p2c),
    .RESET_B(net2280),
    .D(_01504_),
    .Q_N(_05463_),
    .Q(\shift_storage.storage[821] ));
 sg13g2_dfrbp_1 \shift_storage.storage[822]$_SDFFE_PN0P_  (.CLK(clknet_leaf_238_clk_p2c),
    .RESET_B(net2281),
    .D(_01505_),
    .Q_N(_05462_),
    .Q(\shift_storage.storage[822] ));
 sg13g2_dfrbp_1 \shift_storage.storage[823]$_SDFFE_PN0P_  (.CLK(clknet_leaf_238_clk_p2c),
    .RESET_B(net2282),
    .D(_01506_),
    .Q_N(_05461_),
    .Q(\shift_storage.storage[823] ));
 sg13g2_dfrbp_1 \shift_storage.storage[824]$_SDFFE_PN0P_  (.CLK(clknet_leaf_236_clk_p2c),
    .RESET_B(net2283),
    .D(_01507_),
    .Q_N(_05460_),
    .Q(\shift_storage.storage[824] ));
 sg13g2_dfrbp_1 \shift_storage.storage[825]$_SDFFE_PN0P_  (.CLK(clknet_leaf_237_clk_p2c),
    .RESET_B(net2284),
    .D(_01508_),
    .Q_N(_05459_),
    .Q(\shift_storage.storage[825] ));
 sg13g2_dfrbp_1 \shift_storage.storage[826]$_SDFFE_PN0P_  (.CLK(clknet_leaf_237_clk_p2c),
    .RESET_B(net2285),
    .D(_01509_),
    .Q_N(_05458_),
    .Q(\shift_storage.storage[826] ));
 sg13g2_dfrbp_1 \shift_storage.storage[827]$_SDFFE_PN0P_  (.CLK(clknet_leaf_237_clk_p2c),
    .RESET_B(net2286),
    .D(_01510_),
    .Q_N(_05457_),
    .Q(\shift_storage.storage[827] ));
 sg13g2_dfrbp_1 \shift_storage.storage[828]$_SDFFE_PN0P_  (.CLK(clknet_leaf_237_clk_p2c),
    .RESET_B(net2287),
    .D(_01511_),
    .Q_N(_05456_),
    .Q(\shift_storage.storage[828] ));
 sg13g2_dfrbp_1 \shift_storage.storage[829]$_SDFFE_PN0P_  (.CLK(clknet_leaf_236_clk_p2c),
    .RESET_B(net2288),
    .D(_01512_),
    .Q_N(_05455_),
    .Q(\shift_storage.storage[829] ));
 sg13g2_dfrbp_1 \shift_storage.storage[82]$_SDFFE_PN0P_  (.CLK(clknet_leaf_96_clk_p2c),
    .RESET_B(net2289),
    .D(_01513_),
    .Q_N(_05454_),
    .Q(\shift_storage.storage[82] ));
 sg13g2_dfrbp_1 \shift_storage.storage[830]$_SDFFE_PN0P_  (.CLK(clknet_leaf_236_clk_p2c),
    .RESET_B(net2290),
    .D(_01514_),
    .Q_N(_05453_),
    .Q(\shift_storage.storage[830] ));
 sg13g2_dfrbp_1 \shift_storage.storage[831]$_SDFFE_PN0P_  (.CLK(clknet_leaf_236_clk_p2c),
    .RESET_B(net2291),
    .D(_01515_),
    .Q_N(_05452_),
    .Q(\shift_storage.storage[831] ));
 sg13g2_dfrbp_1 \shift_storage.storage[832]$_SDFFE_PN0P_  (.CLK(clknet_leaf_236_clk_p2c),
    .RESET_B(net2292),
    .D(_01516_),
    .Q_N(_05451_),
    .Q(\shift_storage.storage[832] ));
 sg13g2_dfrbp_1 \shift_storage.storage[833]$_SDFFE_PN0P_  (.CLK(clknet_leaf_235_clk_p2c),
    .RESET_B(net2293),
    .D(_01517_),
    .Q_N(_05450_),
    .Q(\shift_storage.storage[833] ));
 sg13g2_dfrbp_1 \shift_storage.storage[834]$_SDFFE_PN0P_  (.CLK(clknet_leaf_233_clk_p2c),
    .RESET_B(net2294),
    .D(_01518_),
    .Q_N(_05449_),
    .Q(\shift_storage.storage[834] ));
 sg13g2_dfrbp_1 \shift_storage.storage[835]$_SDFFE_PN0P_  (.CLK(clknet_leaf_233_clk_p2c),
    .RESET_B(net2295),
    .D(_01519_),
    .Q_N(_05448_),
    .Q(\shift_storage.storage[835] ));
 sg13g2_dfrbp_1 \shift_storage.storage[836]$_SDFFE_PN0P_  (.CLK(clknet_leaf_232_clk_p2c),
    .RESET_B(net2296),
    .D(_01520_),
    .Q_N(_05447_),
    .Q(\shift_storage.storage[836] ));
 sg13g2_dfrbp_1 \shift_storage.storage[837]$_SDFFE_PN0P_  (.CLK(clknet_leaf_232_clk_p2c),
    .RESET_B(net2297),
    .D(_01521_),
    .Q_N(_05446_),
    .Q(\shift_storage.storage[837] ));
 sg13g2_dfrbp_1 \shift_storage.storage[838]$_SDFFE_PN0P_  (.CLK(clknet_leaf_230_clk_p2c),
    .RESET_B(net2298),
    .D(_01522_),
    .Q_N(_05445_),
    .Q(\shift_storage.storage[838] ));
 sg13g2_dfrbp_1 \shift_storage.storage[839]$_SDFFE_PN0P_  (.CLK(clknet_leaf_230_clk_p2c),
    .RESET_B(net2299),
    .D(_01523_),
    .Q_N(_05444_),
    .Q(\shift_storage.storage[839] ));
 sg13g2_dfrbp_1 \shift_storage.storage[83]$_SDFFE_PN0P_  (.CLK(clknet_leaf_96_clk_p2c),
    .RESET_B(net2300),
    .D(_01524_),
    .Q_N(_05443_),
    .Q(\shift_storage.storage[83] ));
 sg13g2_dfrbp_1 \shift_storage.storage[840]$_SDFFE_PN0P_  (.CLK(clknet_leaf_230_clk_p2c),
    .RESET_B(net2301),
    .D(_01525_),
    .Q_N(_05442_),
    .Q(\shift_storage.storage[840] ));
 sg13g2_dfrbp_1 \shift_storage.storage[841]$_SDFFE_PN0P_  (.CLK(clknet_leaf_227_clk_p2c),
    .RESET_B(net2302),
    .D(_01526_),
    .Q_N(_05441_),
    .Q(\shift_storage.storage[841] ));
 sg13g2_dfrbp_1 \shift_storage.storage[842]$_SDFFE_PN0P_  (.CLK(clknet_leaf_227_clk_p2c),
    .RESET_B(net2303),
    .D(_01527_),
    .Q_N(_05440_),
    .Q(\shift_storage.storage[842] ));
 sg13g2_dfrbp_1 \shift_storage.storage[843]$_SDFFE_PN0P_  (.CLK(clknet_leaf_227_clk_p2c),
    .RESET_B(net2304),
    .D(_01528_),
    .Q_N(_05439_),
    .Q(\shift_storage.storage[843] ));
 sg13g2_dfrbp_1 \shift_storage.storage[844]$_SDFFE_PN0P_  (.CLK(clknet_leaf_227_clk_p2c),
    .RESET_B(net2305),
    .D(_01529_),
    .Q_N(_05438_),
    .Q(\shift_storage.storage[844] ));
 sg13g2_dfrbp_1 \shift_storage.storage[845]$_SDFFE_PN0P_  (.CLK(clknet_leaf_228_clk_p2c),
    .RESET_B(net2306),
    .D(_01530_),
    .Q_N(_05437_),
    .Q(\shift_storage.storage[845] ));
 sg13g2_dfrbp_1 \shift_storage.storage[846]$_SDFFE_PN0P_  (.CLK(clknet_leaf_228_clk_p2c),
    .RESET_B(net2307),
    .D(_01531_),
    .Q_N(_05436_),
    .Q(\shift_storage.storage[846] ));
 sg13g2_dfrbp_1 \shift_storage.storage[847]$_SDFFE_PN0P_  (.CLK(clknet_leaf_229_clk_p2c),
    .RESET_B(net2308),
    .D(_01532_),
    .Q_N(_05435_),
    .Q(\shift_storage.storage[847] ));
 sg13g2_dfrbp_1 \shift_storage.storage[848]$_SDFFE_PN0P_  (.CLK(clknet_leaf_230_clk_p2c),
    .RESET_B(net2309),
    .D(_01533_),
    .Q_N(_05434_),
    .Q(\shift_storage.storage[848] ));
 sg13g2_dfrbp_1 \shift_storage.storage[849]$_SDFFE_PN0P_  (.CLK(clknet_leaf_230_clk_p2c),
    .RESET_B(net2310),
    .D(_01534_),
    .Q_N(_05433_),
    .Q(\shift_storage.storage[849] ));
 sg13g2_dfrbp_1 \shift_storage.storage[84]$_SDFFE_PN0P_  (.CLK(clknet_leaf_95_clk_p2c),
    .RESET_B(net2311),
    .D(_01535_),
    .Q_N(_05432_),
    .Q(\shift_storage.storage[84] ));
 sg13g2_dfrbp_1 \shift_storage.storage[850]$_SDFFE_PN0P_  (.CLK(clknet_leaf_229_clk_p2c),
    .RESET_B(net2312),
    .D(_01536_),
    .Q_N(_05431_),
    .Q(\shift_storage.storage[850] ));
 sg13g2_dfrbp_1 \shift_storage.storage[851]$_SDFFE_PN0P_  (.CLK(clknet_leaf_229_clk_p2c),
    .RESET_B(net2313),
    .D(_01537_),
    .Q_N(_05430_),
    .Q(\shift_storage.storage[851] ));
 sg13g2_dfrbp_1 \shift_storage.storage[852]$_SDFFE_PN0P_  (.CLK(clknet_leaf_214_clk_p2c),
    .RESET_B(net2314),
    .D(_01538_),
    .Q_N(_05429_),
    .Q(\shift_storage.storage[852] ));
 sg13g2_dfrbp_1 \shift_storage.storage[853]$_SDFFE_PN0P_  (.CLK(clknet_leaf_214_clk_p2c),
    .RESET_B(net2315),
    .D(_01539_),
    .Q_N(_05428_),
    .Q(\shift_storage.storage[853] ));
 sg13g2_dfrbp_1 \shift_storage.storage[854]$_SDFFE_PN0P_  (.CLK(clknet_leaf_214_clk_p2c),
    .RESET_B(net2316),
    .D(_01540_),
    .Q_N(_05427_),
    .Q(\shift_storage.storage[854] ));
 sg13g2_dfrbp_1 \shift_storage.storage[855]$_SDFFE_PN0P_  (.CLK(clknet_leaf_214_clk_p2c),
    .RESET_B(net2317),
    .D(_01541_),
    .Q_N(_05426_),
    .Q(\shift_storage.storage[855] ));
 sg13g2_dfrbp_1 \shift_storage.storage[856]$_SDFFE_PN0P_  (.CLK(clknet_leaf_214_clk_p2c),
    .RESET_B(net2318),
    .D(_01542_),
    .Q_N(_05425_),
    .Q(\shift_storage.storage[856] ));
 sg13g2_dfrbp_1 \shift_storage.storage[857]$_SDFFE_PN0P_  (.CLK(clknet_leaf_212_clk_p2c),
    .RESET_B(net2319),
    .D(_01543_),
    .Q_N(_05424_),
    .Q(\shift_storage.storage[857] ));
 sg13g2_dfrbp_1 \shift_storage.storage[858]$_SDFFE_PN0P_  (.CLK(clknet_leaf_214_clk_p2c),
    .RESET_B(net2320),
    .D(_01544_),
    .Q_N(_05423_),
    .Q(\shift_storage.storage[858] ));
 sg13g2_dfrbp_1 \shift_storage.storage[859]$_SDFFE_PN0P_  (.CLK(clknet_leaf_213_clk_p2c),
    .RESET_B(net2321),
    .D(_01545_),
    .Q_N(_05422_),
    .Q(\shift_storage.storage[859] ));
 sg13g2_dfrbp_1 \shift_storage.storage[85]$_SDFFE_PN0P_  (.CLK(clknet_leaf_96_clk_p2c),
    .RESET_B(net2322),
    .D(_01546_),
    .Q_N(_05421_),
    .Q(\shift_storage.storage[85] ));
 sg13g2_dfrbp_1 \shift_storage.storage[860]$_SDFFE_PN0P_  (.CLK(clknet_leaf_212_clk_p2c),
    .RESET_B(net2323),
    .D(_01547_),
    .Q_N(_05420_),
    .Q(\shift_storage.storage[860] ));
 sg13g2_dfrbp_1 \shift_storage.storage[861]$_SDFFE_PN0P_  (.CLK(clknet_leaf_212_clk_p2c),
    .RESET_B(net2324),
    .D(_01548_),
    .Q_N(_05419_),
    .Q(\shift_storage.storage[861] ));
 sg13g2_dfrbp_1 \shift_storage.storage[862]$_SDFFE_PN0P_  (.CLK(clknet_leaf_212_clk_p2c),
    .RESET_B(net2325),
    .D(_01549_),
    .Q_N(_05418_),
    .Q(\shift_storage.storage[862] ));
 sg13g2_dfrbp_1 \shift_storage.storage[863]$_SDFFE_PN0P_  (.CLK(clknet_leaf_212_clk_p2c),
    .RESET_B(net2326),
    .D(_01550_),
    .Q_N(_05417_),
    .Q(\shift_storage.storage[863] ));
 sg13g2_dfrbp_1 \shift_storage.storage[864]$_SDFFE_PN0P_  (.CLK(clknet_leaf_195_clk_p2c),
    .RESET_B(net2327),
    .D(_01551_),
    .Q_N(_05416_),
    .Q(\shift_storage.storage[864] ));
 sg13g2_dfrbp_1 \shift_storage.storage[865]$_SDFFE_PN0P_  (.CLK(clknet_leaf_195_clk_p2c),
    .RESET_B(net2328),
    .D(_01552_),
    .Q_N(_05415_),
    .Q(\shift_storage.storage[865] ));
 sg13g2_dfrbp_1 \shift_storage.storage[866]$_SDFFE_PN0P_  (.CLK(clknet_leaf_195_clk_p2c),
    .RESET_B(net2329),
    .D(_01553_),
    .Q_N(_05414_),
    .Q(\shift_storage.storage[866] ));
 sg13g2_dfrbp_1 \shift_storage.storage[867]$_SDFFE_PN0P_  (.CLK(clknet_leaf_211_clk_p2c),
    .RESET_B(net2330),
    .D(_01554_),
    .Q_N(_05413_),
    .Q(\shift_storage.storage[867] ));
 sg13g2_dfrbp_1 \shift_storage.storage[868]$_SDFFE_PN0P_  (.CLK(clknet_leaf_211_clk_p2c),
    .RESET_B(net2331),
    .D(_01555_),
    .Q_N(_05412_),
    .Q(\shift_storage.storage[868] ));
 sg13g2_dfrbp_1 \shift_storage.storage[869]$_SDFFE_PN0P_  (.CLK(clknet_leaf_209_clk_p2c),
    .RESET_B(net2332),
    .D(_01556_),
    .Q_N(_05411_),
    .Q(\shift_storage.storage[869] ));
 sg13g2_dfrbp_1 \shift_storage.storage[86]$_SDFFE_PN0P_  (.CLK(clknet_leaf_95_clk_p2c),
    .RESET_B(net2333),
    .D(_01557_),
    .Q_N(_05410_),
    .Q(\shift_storage.storage[86] ));
 sg13g2_dfrbp_1 \shift_storage.storage[870]$_SDFFE_PN0P_  (.CLK(clknet_leaf_209_clk_p2c),
    .RESET_B(net2334),
    .D(_01558_),
    .Q_N(_05409_),
    .Q(\shift_storage.storage[870] ));
 sg13g2_dfrbp_1 \shift_storage.storage[871]$_SDFFE_PN0P_  (.CLK(clknet_leaf_208_clk_p2c),
    .RESET_B(net2335),
    .D(_01559_),
    .Q_N(_05408_),
    .Q(\shift_storage.storage[871] ));
 sg13g2_dfrbp_1 \shift_storage.storage[872]$_SDFFE_PN0P_  (.CLK(clknet_leaf_208_clk_p2c),
    .RESET_B(net2336),
    .D(_01560_),
    .Q_N(_05407_),
    .Q(\shift_storage.storage[872] ));
 sg13g2_dfrbp_1 \shift_storage.storage[873]$_SDFFE_PN0P_  (.CLK(clknet_leaf_208_clk_p2c),
    .RESET_B(net2337),
    .D(_01561_),
    .Q_N(_05406_),
    .Q(\shift_storage.storage[873] ));
 sg13g2_dfrbp_1 \shift_storage.storage[874]$_SDFFE_PN0P_  (.CLK(clknet_leaf_208_clk_p2c),
    .RESET_B(net2338),
    .D(_01562_),
    .Q_N(_05405_),
    .Q(\shift_storage.storage[874] ));
 sg13g2_dfrbp_1 \shift_storage.storage[875]$_SDFFE_PN0P_  (.CLK(clknet_leaf_217_clk_p2c),
    .RESET_B(net2339),
    .D(_01563_),
    .Q_N(_05404_),
    .Q(\shift_storage.storage[875] ));
 sg13g2_dfrbp_1 \shift_storage.storage[876]$_SDFFE_PN0P_  (.CLK(clknet_leaf_217_clk_p2c),
    .RESET_B(net2340),
    .D(_01564_),
    .Q_N(_05403_),
    .Q(\shift_storage.storage[876] ));
 sg13g2_dfrbp_1 \shift_storage.storage[877]$_SDFFE_PN0P_  (.CLK(clknet_leaf_217_clk_p2c),
    .RESET_B(net2341),
    .D(_01565_),
    .Q_N(_05402_),
    .Q(\shift_storage.storage[877] ));
 sg13g2_dfrbp_1 \shift_storage.storage[878]$_SDFFE_PN0P_  (.CLK(clknet_leaf_217_clk_p2c),
    .RESET_B(net2342),
    .D(_01566_),
    .Q_N(_05401_),
    .Q(\shift_storage.storage[878] ));
 sg13g2_dfrbp_1 \shift_storage.storage[879]$_SDFFE_PN0P_  (.CLK(clknet_leaf_218_clk_p2c),
    .RESET_B(net2343),
    .D(_01567_),
    .Q_N(_05400_),
    .Q(\shift_storage.storage[879] ));
 sg13g2_dfrbp_1 \shift_storage.storage[87]$_SDFFE_PN0P_  (.CLK(clknet_leaf_95_clk_p2c),
    .RESET_B(net2344),
    .D(_01568_),
    .Q_N(_05399_),
    .Q(\shift_storage.storage[87] ));
 sg13g2_dfrbp_1 \shift_storage.storage[880]$_SDFFE_PN0P_  (.CLK(clknet_leaf_218_clk_p2c),
    .RESET_B(net2345),
    .D(_01569_),
    .Q_N(_05398_),
    .Q(\shift_storage.storage[880] ));
 sg13g2_dfrbp_1 \shift_storage.storage[881]$_SDFFE_PN0P_  (.CLK(clknet_leaf_218_clk_p2c),
    .RESET_B(net2346),
    .D(_01570_),
    .Q_N(_05397_),
    .Q(\shift_storage.storage[881] ));
 sg13g2_dfrbp_1 \shift_storage.storage[882]$_SDFFE_PN0P_  (.CLK(clknet_leaf_218_clk_p2c),
    .RESET_B(net2347),
    .D(_01571_),
    .Q_N(_05396_),
    .Q(\shift_storage.storage[882] ));
 sg13g2_dfrbp_1 \shift_storage.storage[883]$_SDFFE_PN0P_  (.CLK(clknet_leaf_218_clk_p2c),
    .RESET_B(net2348),
    .D(_01572_),
    .Q_N(_05395_),
    .Q(\shift_storage.storage[883] ));
 sg13g2_dfrbp_1 \shift_storage.storage[884]$_SDFFE_PN0P_  (.CLK(clknet_leaf_219_clk_p2c),
    .RESET_B(net2349),
    .D(_01573_),
    .Q_N(_05394_),
    .Q(\shift_storage.storage[884] ));
 sg13g2_dfrbp_1 \shift_storage.storage[885]$_SDFFE_PN0P_  (.CLK(clknet_leaf_219_clk_p2c),
    .RESET_B(net2350),
    .D(_01574_),
    .Q_N(_05393_),
    .Q(\shift_storage.storage[885] ));
 sg13g2_dfrbp_1 \shift_storage.storage[886]$_SDFFE_PN0P_  (.CLK(clknet_leaf_219_clk_p2c),
    .RESET_B(net2351),
    .D(_01575_),
    .Q_N(_05392_),
    .Q(\shift_storage.storage[886] ));
 sg13g2_dfrbp_1 \shift_storage.storage[887]$_SDFFE_PN0P_  (.CLK(clknet_leaf_216_clk_p2c),
    .RESET_B(net2352),
    .D(_01576_),
    .Q_N(_05391_),
    .Q(\shift_storage.storage[887] ));
 sg13g2_dfrbp_1 \shift_storage.storage[888]$_SDFFE_PN0P_  (.CLK(clknet_leaf_216_clk_p2c),
    .RESET_B(net2353),
    .D(_01577_),
    .Q_N(_05390_),
    .Q(\shift_storage.storage[888] ));
 sg13g2_dfrbp_1 \shift_storage.storage[889]$_SDFFE_PN0P_  (.CLK(clknet_leaf_216_clk_p2c),
    .RESET_B(net2354),
    .D(_01578_),
    .Q_N(_05389_),
    .Q(\shift_storage.storage[889] ));
 sg13g2_dfrbp_1 \shift_storage.storage[88]$_SDFFE_PN0P_  (.CLK(clknet_leaf_95_clk_p2c),
    .RESET_B(net2355),
    .D(_01579_),
    .Q_N(_05388_),
    .Q(\shift_storage.storage[88] ));
 sg13g2_dfrbp_1 \shift_storage.storage[890]$_SDFFE_PN0P_  (.CLK(clknet_leaf_216_clk_p2c),
    .RESET_B(net2356),
    .D(_01580_),
    .Q_N(_05387_),
    .Q(\shift_storage.storage[890] ));
 sg13g2_dfrbp_1 \shift_storage.storage[891]$_SDFFE_PN0P_  (.CLK(clknet_leaf_216_clk_p2c),
    .RESET_B(net2357),
    .D(_01581_),
    .Q_N(_05386_),
    .Q(\shift_storage.storage[891] ));
 sg13g2_dfrbp_1 \shift_storage.storage[892]$_SDFFE_PN0P_  (.CLK(clknet_leaf_216_clk_p2c),
    .RESET_B(net2358),
    .D(_01582_),
    .Q_N(_05385_),
    .Q(\shift_storage.storage[892] ));
 sg13g2_dfrbp_1 \shift_storage.storage[893]$_SDFFE_PN0P_  (.CLK(clknet_leaf_217_clk_p2c),
    .RESET_B(net2359),
    .D(_01583_),
    .Q_N(_05384_),
    .Q(\shift_storage.storage[893] ));
 sg13g2_dfrbp_1 \shift_storage.storage[894]$_SDFFE_PN0P_  (.CLK(clknet_leaf_211_clk_p2c),
    .RESET_B(net2360),
    .D(_01584_),
    .Q_N(_05383_),
    .Q(\shift_storage.storage[894] ));
 sg13g2_dfrbp_1 \shift_storage.storage[895]$_SDFFE_PN0P_  (.CLK(clknet_leaf_211_clk_p2c),
    .RESET_B(net2361),
    .D(_01585_),
    .Q_N(_05382_),
    .Q(\shift_storage.storage[895] ));
 sg13g2_dfrbp_1 \shift_storage.storage[896]$_SDFFE_PN0P_  (.CLK(clknet_leaf_211_clk_p2c),
    .RESET_B(net2362),
    .D(_01586_),
    .Q_N(_05381_),
    .Q(\shift_storage.storage[896] ));
 sg13g2_dfrbp_1 \shift_storage.storage[897]$_SDFFE_PN0P_  (.CLK(clknet_leaf_211_clk_p2c),
    .RESET_B(net2363),
    .D(_01587_),
    .Q_N(_05380_),
    .Q(\shift_storage.storage[897] ));
 sg13g2_dfrbp_1 \shift_storage.storage[898]$_SDFFE_PN0P_  (.CLK(clknet_leaf_211_clk_p2c),
    .RESET_B(net2364),
    .D(_01588_),
    .Q_N(_05379_),
    .Q(\shift_storage.storage[898] ));
 sg13g2_dfrbp_1 \shift_storage.storage[899]$_SDFFE_PN0P_  (.CLK(clknet_leaf_210_clk_p2c),
    .RESET_B(net2365),
    .D(_01589_),
    .Q_N(_05378_),
    .Q(\shift_storage.storage[899] ));
 sg13g2_dfrbp_1 \shift_storage.storage[89]$_SDFFE_PN0P_  (.CLK(clknet_leaf_48_clk_p2c),
    .RESET_B(net2366),
    .D(_01590_),
    .Q_N(_05377_),
    .Q(\shift_storage.storage[89] ));
 sg13g2_dfrbp_1 \shift_storage.storage[8]$_SDFFE_PN0P_  (.CLK(clknet_leaf_73_clk_p2c),
    .RESET_B(net2367),
    .D(_01591_),
    .Q_N(_05376_),
    .Q(\shift_storage.storage[8] ));
 sg13g2_dfrbp_1 \shift_storage.storage[900]$_SDFFE_PN0P_  (.CLK(clknet_leaf_210_clk_p2c),
    .RESET_B(net2368),
    .D(_01592_),
    .Q_N(_05375_),
    .Q(\shift_storage.storage[900] ));
 sg13g2_dfrbp_1 \shift_storage.storage[901]$_SDFFE_PN0P_  (.CLK(clknet_leaf_210_clk_p2c),
    .RESET_B(net2369),
    .D(_01593_),
    .Q_N(_05374_),
    .Q(\shift_storage.storage[901] ));
 sg13g2_dfrbp_1 \shift_storage.storage[902]$_SDFFE_PN0P_  (.CLK(clknet_leaf_209_clk_p2c),
    .RESET_B(net2370),
    .D(_01594_),
    .Q_N(_05373_),
    .Q(\shift_storage.storage[902] ));
 sg13g2_dfrbp_1 \shift_storage.storage[903]$_SDFFE_PN0P_  (.CLK(clknet_leaf_209_clk_p2c),
    .RESET_B(net2371),
    .D(_01595_),
    .Q_N(_05372_),
    .Q(\shift_storage.storage[903] ));
 sg13g2_dfrbp_1 \shift_storage.storage[904]$_SDFFE_PN0P_  (.CLK(clknet_leaf_209_clk_p2c),
    .RESET_B(net2372),
    .D(_01596_),
    .Q_N(_05371_),
    .Q(\shift_storage.storage[904] ));
 sg13g2_dfrbp_1 \shift_storage.storage[905]$_SDFFE_PN0P_  (.CLK(clknet_leaf_209_clk_p2c),
    .RESET_B(net2373),
    .D(_01597_),
    .Q_N(_05370_),
    .Q(\shift_storage.storage[905] ));
 sg13g2_dfrbp_1 \shift_storage.storage[906]$_SDFFE_PN0P_  (.CLK(clknet_leaf_207_clk_p2c),
    .RESET_B(net2374),
    .D(_01598_),
    .Q_N(_05369_),
    .Q(\shift_storage.storage[906] ));
 sg13g2_dfrbp_1 \shift_storage.storage[907]$_SDFFE_PN0P_  (.CLK(clknet_leaf_207_clk_p2c),
    .RESET_B(net2375),
    .D(_01599_),
    .Q_N(_05368_),
    .Q(\shift_storage.storage[907] ));
 sg13g2_dfrbp_1 \shift_storage.storage[908]$_SDFFE_PN0P_  (.CLK(clknet_leaf_207_clk_p2c),
    .RESET_B(net2376),
    .D(_01600_),
    .Q_N(_05367_),
    .Q(\shift_storage.storage[908] ));
 sg13g2_dfrbp_1 \shift_storage.storage[909]$_SDFFE_PN0P_  (.CLK(clknet_leaf_206_clk_p2c),
    .RESET_B(net2377),
    .D(_01601_),
    .Q_N(_05366_),
    .Q(\shift_storage.storage[909] ));
 sg13g2_dfrbp_1 \shift_storage.storage[90]$_SDFFE_PN0P_  (.CLK(clknet_leaf_48_clk_p2c),
    .RESET_B(net2378),
    .D(_01602_),
    .Q_N(_05365_),
    .Q(\shift_storage.storage[90] ));
 sg13g2_dfrbp_1 \shift_storage.storage[910]$_SDFFE_PN0P_  (.CLK(clknet_leaf_207_clk_p2c),
    .RESET_B(net2379),
    .D(_01603_),
    .Q_N(_05364_),
    .Q(\shift_storage.storage[910] ));
 sg13g2_dfrbp_1 \shift_storage.storage[911]$_SDFFE_PN0P_  (.CLK(clknet_leaf_207_clk_p2c),
    .RESET_B(net2380),
    .D(_01604_),
    .Q_N(_05363_),
    .Q(\shift_storage.storage[911] ));
 sg13g2_dfrbp_1 \shift_storage.storage[912]$_SDFFE_PN0P_  (.CLK(clknet_leaf_207_clk_p2c),
    .RESET_B(net2381),
    .D(_01605_),
    .Q_N(_05362_),
    .Q(\shift_storage.storage[912] ));
 sg13g2_dfrbp_1 \shift_storage.storage[913]$_SDFFE_PN0P_  (.CLK(clknet_leaf_208_clk_p2c),
    .RESET_B(net2382),
    .D(_01606_),
    .Q_N(_05361_),
    .Q(\shift_storage.storage[913] ));
 sg13g2_dfrbp_1 \shift_storage.storage[914]$_SDFFE_PN0P_  (.CLK(clknet_leaf_205_clk_p2c),
    .RESET_B(net2383),
    .D(_01607_),
    .Q_N(_05360_),
    .Q(\shift_storage.storage[914] ));
 sg13g2_dfrbp_1 \shift_storage.storage[915]$_SDFFE_PN0P_  (.CLK(clknet_leaf_205_clk_p2c),
    .RESET_B(net2384),
    .D(_01608_),
    .Q_N(_05359_),
    .Q(\shift_storage.storage[915] ));
 sg13g2_dfrbp_1 \shift_storage.storage[916]$_SDFFE_PN0P_  (.CLK(clknet_leaf_205_clk_p2c),
    .RESET_B(net2385),
    .D(_01609_),
    .Q_N(_05358_),
    .Q(\shift_storage.storage[916] ));
 sg13g2_dfrbp_1 \shift_storage.storage[917]$_SDFFE_PN0P_  (.CLK(clknet_leaf_205_clk_p2c),
    .RESET_B(net2386),
    .D(_01610_),
    .Q_N(_05357_),
    .Q(\shift_storage.storage[917] ));
 sg13g2_dfrbp_1 \shift_storage.storage[918]$_SDFFE_PN0P_  (.CLK(clknet_leaf_206_clk_p2c),
    .RESET_B(net2387),
    .D(_01611_),
    .Q_N(_05356_),
    .Q(\shift_storage.storage[918] ));
 sg13g2_dfrbp_1 \shift_storage.storage[919]$_SDFFE_PN0P_  (.CLK(clknet_leaf_206_clk_p2c),
    .RESET_B(net2388),
    .D(_01612_),
    .Q_N(_05355_),
    .Q(\shift_storage.storage[919] ));
 sg13g2_dfrbp_1 \shift_storage.storage[91]$_SDFFE_PN0P_  (.CLK(clknet_leaf_47_clk_p2c),
    .RESET_B(net2389),
    .D(_01613_),
    .Q_N(_05354_),
    .Q(\shift_storage.storage[91] ));
 sg13g2_dfrbp_1 \shift_storage.storage[920]$_SDFFE_PN0P_  (.CLK(clknet_leaf_201_clk_p2c),
    .RESET_B(net2390),
    .D(_01614_),
    .Q_N(_05353_),
    .Q(\shift_storage.storage[920] ));
 sg13g2_dfrbp_1 \shift_storage.storage[921]$_SDFFE_PN0P_  (.CLK(clknet_leaf_201_clk_p2c),
    .RESET_B(net2391),
    .D(_01615_),
    .Q_N(_05352_),
    .Q(\shift_storage.storage[921] ));
 sg13g2_dfrbp_1 \shift_storage.storage[922]$_SDFFE_PN0P_  (.CLK(clknet_leaf_202_clk_p2c),
    .RESET_B(net2392),
    .D(_01616_),
    .Q_N(_05351_),
    .Q(\shift_storage.storage[922] ));
 sg13g2_dfrbp_1 \shift_storage.storage[923]$_SDFFE_PN0P_  (.CLK(clknet_leaf_202_clk_p2c),
    .RESET_B(net2393),
    .D(_01617_),
    .Q_N(_05350_),
    .Q(\shift_storage.storage[923] ));
 sg13g2_dfrbp_1 \shift_storage.storage[924]$_SDFFE_PN0P_  (.CLK(clknet_leaf_201_clk_p2c),
    .RESET_B(net2394),
    .D(_01618_),
    .Q_N(_05349_),
    .Q(\shift_storage.storage[924] ));
 sg13g2_dfrbp_1 \shift_storage.storage[925]$_SDFFE_PN0P_  (.CLK(clknet_leaf_199_clk_p2c),
    .RESET_B(net2395),
    .D(_01619_),
    .Q_N(_05348_),
    .Q(\shift_storage.storage[925] ));
 sg13g2_dfrbp_1 \shift_storage.storage[926]$_SDFFE_PN0P_  (.CLK(clknet_leaf_199_clk_p2c),
    .RESET_B(net2396),
    .D(_01620_),
    .Q_N(_05347_),
    .Q(\shift_storage.storage[926] ));
 sg13g2_dfrbp_1 \shift_storage.storage[927]$_SDFFE_PN0P_  (.CLK(clknet_leaf_199_clk_p2c),
    .RESET_B(net2397),
    .D(_01621_),
    .Q_N(_05346_),
    .Q(\shift_storage.storage[927] ));
 sg13g2_dfrbp_1 \shift_storage.storage[928]$_SDFFE_PN0P_  (.CLK(clknet_leaf_202_clk_p2c),
    .RESET_B(net2398),
    .D(_01622_),
    .Q_N(_05345_),
    .Q(\shift_storage.storage[928] ));
 sg13g2_dfrbp_1 \shift_storage.storage[929]$_SDFFE_PN0P_  (.CLK(clknet_leaf_202_clk_p2c),
    .RESET_B(net2399),
    .D(_01623_),
    .Q_N(_05344_),
    .Q(\shift_storage.storage[929] ));
 sg13g2_dfrbp_1 \shift_storage.storage[92]$_SDFFE_PN0P_  (.CLK(clknet_leaf_47_clk_p2c),
    .RESET_B(net2400),
    .D(_01624_),
    .Q_N(_05343_),
    .Q(\shift_storage.storage[92] ));
 sg13g2_dfrbp_1 \shift_storage.storage[930]$_SDFFE_PN0P_  (.CLK(clknet_leaf_202_clk_p2c),
    .RESET_B(net2401),
    .D(_01625_),
    .Q_N(_05342_),
    .Q(\shift_storage.storage[930] ));
 sg13g2_dfrbp_1 \shift_storage.storage[931]$_SDFFE_PN0P_  (.CLK(clknet_leaf_202_clk_p2c),
    .RESET_B(net2402),
    .D(_01626_),
    .Q_N(_05341_),
    .Q(\shift_storage.storage[931] ));
 sg13g2_dfrbp_1 \shift_storage.storage[932]$_SDFFE_PN0P_  (.CLK(clknet_leaf_203_clk_p2c),
    .RESET_B(net2403),
    .D(_01627_),
    .Q_N(_05340_),
    .Q(\shift_storage.storage[932] ));
 sg13g2_dfrbp_1 \shift_storage.storage[933]$_SDFFE_PN0P_  (.CLK(clknet_leaf_203_clk_p2c),
    .RESET_B(net2404),
    .D(_01628_),
    .Q_N(_05339_),
    .Q(\shift_storage.storage[933] ));
 sg13g2_dfrbp_1 \shift_storage.storage[934]$_SDFFE_PN0P_  (.CLK(clknet_leaf_203_clk_p2c),
    .RESET_B(net2405),
    .D(_01629_),
    .Q_N(_05338_),
    .Q(\shift_storage.storage[934] ));
 sg13g2_dfrbp_1 \shift_storage.storage[935]$_SDFFE_PN0P_  (.CLK(clknet_leaf_203_clk_p2c),
    .RESET_B(net2406),
    .D(_01630_),
    .Q_N(_05337_),
    .Q(\shift_storage.storage[935] ));
 sg13g2_dfrbp_1 \shift_storage.storage[936]$_SDFFE_PN0P_  (.CLK(clknet_leaf_203_clk_p2c),
    .RESET_B(net2407),
    .D(_01631_),
    .Q_N(_05336_),
    .Q(\shift_storage.storage[936] ));
 sg13g2_dfrbp_1 \shift_storage.storage[937]$_SDFFE_PN0P_  (.CLK(clknet_leaf_204_clk_p2c),
    .RESET_B(net2408),
    .D(_01632_),
    .Q_N(_05335_),
    .Q(\shift_storage.storage[937] ));
 sg13g2_dfrbp_1 \shift_storage.storage[938]$_SDFFE_PN0P_  (.CLK(clknet_leaf_204_clk_p2c),
    .RESET_B(net2409),
    .D(_01633_),
    .Q_N(_05334_),
    .Q(\shift_storage.storage[938] ));
 sg13g2_dfrbp_1 \shift_storage.storage[939]$_SDFFE_PN0P_  (.CLK(clknet_leaf_204_clk_p2c),
    .RESET_B(net2410),
    .D(_01634_),
    .Q_N(_05333_),
    .Q(\shift_storage.storage[939] ));
 sg13g2_dfrbp_1 \shift_storage.storage[93]$_SDFFE_PN0P_  (.CLK(clknet_leaf_46_clk_p2c),
    .RESET_B(net2411),
    .D(_01635_),
    .Q_N(_05332_),
    .Q(\shift_storage.storage[93] ));
 sg13g2_dfrbp_1 \shift_storage.storage[940]$_SDFFE_PN0P_  (.CLK(clknet_leaf_205_clk_p2c),
    .RESET_B(net2412),
    .D(_01636_),
    .Q_N(_05331_),
    .Q(\shift_storage.storage[940] ));
 sg13g2_dfrbp_1 \shift_storage.storage[941]$_SDFFE_PN0P_  (.CLK(clknet_leaf_204_clk_p2c),
    .RESET_B(net2413),
    .D(_01637_),
    .Q_N(_05330_),
    .Q(\shift_storage.storage[941] ));
 sg13g2_dfrbp_1 \shift_storage.storage[942]$_SDFFE_PN0P_  (.CLK(clknet_leaf_204_clk_p2c),
    .RESET_B(net2414),
    .D(_01638_),
    .Q_N(_05329_),
    .Q(\shift_storage.storage[942] ));
 sg13g2_dfrbp_1 \shift_storage.storage[943]$_SDFFE_PN0P_  (.CLK(clknet_leaf_204_clk_p2c),
    .RESET_B(net2415),
    .D(_01639_),
    .Q_N(_05328_),
    .Q(\shift_storage.storage[943] ));
 sg13g2_dfrbp_1 \shift_storage.storage[944]$_SDFFE_PN0P_  (.CLK(clknet_leaf_205_clk_p2c),
    .RESET_B(net2416),
    .D(_01640_),
    .Q_N(_05327_),
    .Q(\shift_storage.storage[944] ));
 sg13g2_dfrbp_1 \shift_storage.storage[945]$_SDFFE_PN0P_  (.CLK(clknet_leaf_206_clk_p2c),
    .RESET_B(net2417),
    .D(_01641_),
    .Q_N(_05326_),
    .Q(\shift_storage.storage[945] ));
 sg13g2_dfrbp_1 \shift_storage.storage[946]$_SDFFE_PN0P_  (.CLK(clknet_leaf_206_clk_p2c),
    .RESET_B(net2418),
    .D(_01642_),
    .Q_N(_05325_),
    .Q(\shift_storage.storage[946] ));
 sg13g2_dfrbp_1 \shift_storage.storage[947]$_SDFFE_PN0P_  (.CLK(clknet_leaf_206_clk_p2c),
    .RESET_B(net2419),
    .D(_01643_),
    .Q_N(_05324_),
    .Q(\shift_storage.storage[947] ));
 sg13g2_dfrbp_1 \shift_storage.storage[948]$_SDFFE_PN0P_  (.CLK(clknet_leaf_201_clk_p2c),
    .RESET_B(net2420),
    .D(_01644_),
    .Q_N(_05323_),
    .Q(\shift_storage.storage[948] ));
 sg13g2_dfrbp_1 \shift_storage.storage[949]$_SDFFE_PN0P_  (.CLK(clknet_leaf_201_clk_p2c),
    .RESET_B(net2421),
    .D(_01645_),
    .Q_N(_05322_),
    .Q(\shift_storage.storage[949] ));
 sg13g2_dfrbp_1 \shift_storage.storage[94]$_SDFFE_PN0P_  (.CLK(clknet_leaf_46_clk_p2c),
    .RESET_B(net2422),
    .D(_01646_),
    .Q_N(_05321_),
    .Q(\shift_storage.storage[94] ));
 sg13g2_dfrbp_1 \shift_storage.storage[950]$_SDFFE_PN0P_  (.CLK(clknet_leaf_201_clk_p2c),
    .RESET_B(net2423),
    .D(_01647_),
    .Q_N(_05320_),
    .Q(\shift_storage.storage[950] ));
 sg13g2_dfrbp_1 \shift_storage.storage[951]$_SDFFE_PN0P_  (.CLK(clknet_leaf_200_clk_p2c),
    .RESET_B(net2424),
    .D(_01648_),
    .Q_N(_05319_),
    .Q(\shift_storage.storage[951] ));
 sg13g2_dfrbp_1 \shift_storage.storage[952]$_SDFFE_PN0P_  (.CLK(clknet_leaf_200_clk_p2c),
    .RESET_B(net2425),
    .D(_01649_),
    .Q_N(_05318_),
    .Q(\shift_storage.storage[952] ));
 sg13g2_dfrbp_1 \shift_storage.storage[953]$_SDFFE_PN0P_  (.CLK(clknet_leaf_196_clk_p2c),
    .RESET_B(net2426),
    .D(_01650_),
    .Q_N(_05317_),
    .Q(\shift_storage.storage[953] ));
 sg13g2_dfrbp_1 \shift_storage.storage[954]$_SDFFE_PN0P_  (.CLK(clknet_leaf_210_clk_p2c),
    .RESET_B(net2427),
    .D(_01651_),
    .Q_N(_05316_),
    .Q(\shift_storage.storage[954] ));
 sg13g2_dfrbp_1 \shift_storage.storage[955]$_SDFFE_PN0P_  (.CLK(clknet_leaf_210_clk_p2c),
    .RESET_B(net2428),
    .D(_01652_),
    .Q_N(_05315_),
    .Q(\shift_storage.storage[955] ));
 sg13g2_dfrbp_1 \shift_storage.storage[956]$_SDFFE_PN0P_  (.CLK(clknet_leaf_195_clk_p2c),
    .RESET_B(net2429),
    .D(_01653_),
    .Q_N(_05314_),
    .Q(\shift_storage.storage[956] ));
 sg13g2_dfrbp_1 \shift_storage.storage[957]$_SDFFE_PN0P_  (.CLK(clknet_leaf_195_clk_p2c),
    .RESET_B(net2430),
    .D(_01654_),
    .Q_N(_05313_),
    .Q(\shift_storage.storage[957] ));
 sg13g2_dfrbp_1 \shift_storage.storage[958]$_SDFFE_PN0P_  (.CLK(clknet_leaf_195_clk_p2c),
    .RESET_B(net2431),
    .D(_01655_),
    .Q_N(_05312_),
    .Q(\shift_storage.storage[958] ));
 sg13g2_dfrbp_1 \shift_storage.storage[959]$_SDFFE_PN0P_  (.CLK(clknet_leaf_195_clk_p2c),
    .RESET_B(net2432),
    .D(_01656_),
    .Q_N(_05311_),
    .Q(\shift_storage.storage[959] ));
 sg13g2_dfrbp_1 \shift_storage.storage[95]$_SDFFE_PN0P_  (.CLK(clknet_leaf_47_clk_p2c),
    .RESET_B(net2433),
    .D(_01657_),
    .Q_N(_05310_),
    .Q(\shift_storage.storage[95] ));
 sg13g2_dfrbp_1 \shift_storage.storage[960]$_SDFFE_PN0P_  (.CLK(clknet_leaf_194_clk_p2c),
    .RESET_B(net2434),
    .D(_01658_),
    .Q_N(_05309_),
    .Q(\shift_storage.storage[960] ));
 sg13g2_dfrbp_1 \shift_storage.storage[961]$_SDFFE_PN0P_  (.CLK(clknet_leaf_194_clk_p2c),
    .RESET_B(net2435),
    .D(_01659_),
    .Q_N(_05308_),
    .Q(\shift_storage.storage[961] ));
 sg13g2_dfrbp_1 \shift_storage.storage[962]$_SDFFE_PN0P_  (.CLK(clknet_leaf_194_clk_p2c),
    .RESET_B(net2436),
    .D(_01660_),
    .Q_N(_05307_),
    .Q(\shift_storage.storage[962] ));
 sg13g2_dfrbp_1 \shift_storage.storage[963]$_SDFFE_PN0P_  (.CLK(clknet_leaf_192_clk_p2c),
    .RESET_B(net2437),
    .D(_01661_),
    .Q_N(_05306_),
    .Q(\shift_storage.storage[963] ));
 sg13g2_dfrbp_1 \shift_storage.storage[964]$_SDFFE_PN0P_  (.CLK(clknet_leaf_192_clk_p2c),
    .RESET_B(net2438),
    .D(_01662_),
    .Q_N(_05305_),
    .Q(\shift_storage.storage[964] ));
 sg13g2_dfrbp_1 \shift_storage.storage[965]$_SDFFE_PN0P_  (.CLK(clknet_leaf_190_clk_p2c),
    .RESET_B(net2439),
    .D(_01663_),
    .Q_N(_05304_),
    .Q(\shift_storage.storage[965] ));
 sg13g2_dfrbp_1 \shift_storage.storage[966]$_SDFFE_PN0P_  (.CLK(clknet_leaf_190_clk_p2c),
    .RESET_B(net2440),
    .D(_01664_),
    .Q_N(_05303_),
    .Q(\shift_storage.storage[966] ));
 sg13g2_dfrbp_1 \shift_storage.storage[967]$_SDFFE_PN0P_  (.CLK(clknet_leaf_197_clk_p2c),
    .RESET_B(net2441),
    .D(_01665_),
    .Q_N(_05302_),
    .Q(\shift_storage.storage[967] ));
 sg13g2_dfrbp_1 \shift_storage.storage[968]$_SDFFE_PN0P_  (.CLK(clknet_leaf_197_clk_p2c),
    .RESET_B(net2442),
    .D(_01666_),
    .Q_N(_05301_),
    .Q(\shift_storage.storage[968] ));
 sg13g2_dfrbp_1 \shift_storage.storage[969]$_SDFFE_PN0P_  (.CLK(clknet_leaf_197_clk_p2c),
    .RESET_B(net2443),
    .D(_01667_),
    .Q_N(_05300_),
    .Q(\shift_storage.storage[969] ));
 sg13g2_dfrbp_1 \shift_storage.storage[96]$_SDFFE_PN0P_  (.CLK(clknet_leaf_44_clk_p2c),
    .RESET_B(net2444),
    .D(_01668_),
    .Q_N(_05299_),
    .Q(\shift_storage.storage[96] ));
 sg13g2_dfrbp_1 \shift_storage.storage[970]$_SDFFE_PN0P_  (.CLK(clknet_leaf_197_clk_p2c),
    .RESET_B(net2445),
    .D(_01669_),
    .Q_N(_05298_),
    .Q(\shift_storage.storage[970] ));
 sg13g2_dfrbp_1 \shift_storage.storage[971]$_SDFFE_PN0P_  (.CLK(clknet_leaf_198_clk_p2c),
    .RESET_B(net2446),
    .D(_01670_),
    .Q_N(_05297_),
    .Q(\shift_storage.storage[971] ));
 sg13g2_dfrbp_1 \shift_storage.storage[972]$_SDFFE_PN0P_  (.CLK(clknet_leaf_197_clk_p2c),
    .RESET_B(net2447),
    .D(_01671_),
    .Q_N(_05296_),
    .Q(\shift_storage.storage[972] ));
 sg13g2_dfrbp_1 \shift_storage.storage[973]$_SDFFE_PN0P_  (.CLK(clknet_leaf_196_clk_p2c),
    .RESET_B(net2448),
    .D(_01672_),
    .Q_N(_05295_),
    .Q(\shift_storage.storage[973] ));
 sg13g2_dfrbp_1 \shift_storage.storage[974]$_SDFFE_PN0P_  (.CLK(clknet_leaf_196_clk_p2c),
    .RESET_B(net2449),
    .D(_01673_),
    .Q_N(_05294_),
    .Q(\shift_storage.storage[974] ));
 sg13g2_dfrbp_1 \shift_storage.storage[975]$_SDFFE_PN0P_  (.CLK(clknet_leaf_196_clk_p2c),
    .RESET_B(net2450),
    .D(_01674_),
    .Q_N(_05293_),
    .Q(\shift_storage.storage[975] ));
 sg13g2_dfrbp_1 \shift_storage.storage[976]$_SDFFE_PN0P_  (.CLK(clknet_leaf_196_clk_p2c),
    .RESET_B(net2451),
    .D(_01675_),
    .Q_N(_05292_),
    .Q(\shift_storage.storage[976] ));
 sg13g2_dfrbp_1 \shift_storage.storage[977]$_SDFFE_PN0P_  (.CLK(clknet_leaf_196_clk_p2c),
    .RESET_B(net2452),
    .D(_01676_),
    .Q_N(_05291_),
    .Q(\shift_storage.storage[977] ));
 sg13g2_dfrbp_1 \shift_storage.storage[978]$_SDFFE_PN0P_  (.CLK(clknet_leaf_200_clk_p2c),
    .RESET_B(net2453),
    .D(_01677_),
    .Q_N(_05290_),
    .Q(\shift_storage.storage[978] ));
 sg13g2_dfrbp_1 \shift_storage.storage[979]$_SDFFE_PN0P_  (.CLK(clknet_leaf_200_clk_p2c),
    .RESET_B(net2454),
    .D(_01678_),
    .Q_N(_05289_),
    .Q(\shift_storage.storage[979] ));
 sg13g2_dfrbp_1 \shift_storage.storage[97]$_SDFFE_PN0P_  (.CLK(clknet_leaf_44_clk_p2c),
    .RESET_B(net2455),
    .D(_01679_),
    .Q_N(_05288_),
    .Q(\shift_storage.storage[97] ));
 sg13g2_dfrbp_1 \shift_storage.storage[980]$_SDFFE_PN0P_  (.CLK(clknet_leaf_200_clk_p2c),
    .RESET_B(net2456),
    .D(_01680_),
    .Q_N(_05287_),
    .Q(\shift_storage.storage[980] ));
 sg13g2_dfrbp_1 \shift_storage.storage[981]$_SDFFE_PN0P_  (.CLK(clknet_leaf_199_clk_p2c),
    .RESET_B(net2457),
    .D(_01681_),
    .Q_N(_05286_),
    .Q(\shift_storage.storage[981] ));
 sg13g2_dfrbp_1 \shift_storage.storage[982]$_SDFFE_PN0P_  (.CLK(clknet_leaf_199_clk_p2c),
    .RESET_B(net2458),
    .D(_01682_),
    .Q_N(_05285_),
    .Q(\shift_storage.storage[982] ));
 sg13g2_dfrbp_1 \shift_storage.storage[983]$_SDFFE_PN0P_  (.CLK(clknet_leaf_199_clk_p2c),
    .RESET_B(net2459),
    .D(_01683_),
    .Q_N(_05284_),
    .Q(\shift_storage.storage[983] ));
 sg13g2_dfrbp_1 \shift_storage.storage[984]$_SDFFE_PN0P_  (.CLK(clknet_leaf_198_clk_p2c),
    .RESET_B(net2460),
    .D(_01684_),
    .Q_N(_05283_),
    .Q(\shift_storage.storage[984] ));
 sg13g2_dfrbp_1 \shift_storage.storage[985]$_SDFFE_PN0P_  (.CLK(clknet_leaf_198_clk_p2c),
    .RESET_B(net2461),
    .D(_01685_),
    .Q_N(_05282_),
    .Q(\shift_storage.storage[985] ));
 sg13g2_dfrbp_1 \shift_storage.storage[986]$_SDFFE_PN0P_  (.CLK(clknet_leaf_198_clk_p2c),
    .RESET_B(net2462),
    .D(_01686_),
    .Q_N(_05281_),
    .Q(\shift_storage.storage[986] ));
 sg13g2_dfrbp_1 \shift_storage.storage[987]$_SDFFE_PN0P_  (.CLK(clknet_leaf_198_clk_p2c),
    .RESET_B(net2463),
    .D(_01687_),
    .Q_N(_05280_),
    .Q(\shift_storage.storage[987] ));
 sg13g2_dfrbp_1 \shift_storage.storage[988]$_SDFFE_PN0P_  (.CLK(clknet_leaf_198_clk_p2c),
    .RESET_B(net2464),
    .D(_01688_),
    .Q_N(_05279_),
    .Q(\shift_storage.storage[988] ));
 sg13g2_dfrbp_1 \shift_storage.storage[989]$_SDFFE_PN0P_  (.CLK(clknet_leaf_189_clk_p2c),
    .RESET_B(net2465),
    .D(_01689_),
    .Q_N(_05278_),
    .Q(\shift_storage.storage[989] ));
 sg13g2_dfrbp_1 \shift_storage.storage[98]$_SDFFE_PN0P_  (.CLK(clknet_leaf_43_clk_p2c),
    .RESET_B(net2466),
    .D(_01690_),
    .Q_N(_05277_),
    .Q(\shift_storage.storage[98] ));
 sg13g2_dfrbp_1 \shift_storage.storage[990]$_SDFFE_PN0P_  (.CLK(clknet_leaf_189_clk_p2c),
    .RESET_B(net2467),
    .D(_01691_),
    .Q_N(_05276_),
    .Q(\shift_storage.storage[990] ));
 sg13g2_dfrbp_1 \shift_storage.storage[991]$_SDFFE_PN0P_  (.CLK(clknet_leaf_189_clk_p2c),
    .RESET_B(net2468),
    .D(_01692_),
    .Q_N(_05275_),
    .Q(\shift_storage.storage[991] ));
 sg13g2_dfrbp_1 \shift_storage.storage[992]$_SDFFE_PN0P_  (.CLK(clknet_leaf_188_clk_p2c),
    .RESET_B(net2469),
    .D(_01693_),
    .Q_N(_05274_),
    .Q(\shift_storage.storage[992] ));
 sg13g2_dfrbp_1 \shift_storage.storage[993]$_SDFFE_PN0P_  (.CLK(clknet_leaf_188_clk_p2c),
    .RESET_B(net2470),
    .D(_01694_),
    .Q_N(_05273_),
    .Q(\shift_storage.storage[993] ));
 sg13g2_dfrbp_1 \shift_storage.storage[994]$_SDFFE_PN0P_  (.CLK(clknet_leaf_188_clk_p2c),
    .RESET_B(net2471),
    .D(_01695_),
    .Q_N(_05272_),
    .Q(\shift_storage.storage[994] ));
 sg13g2_dfrbp_1 \shift_storage.storage[995]$_SDFFE_PN0P_  (.CLK(clknet_leaf_189_clk_p2c),
    .RESET_B(net2472),
    .D(_01696_),
    .Q_N(_05271_),
    .Q(\shift_storage.storage[995] ));
 sg13g2_dfrbp_1 \shift_storage.storage[996]$_SDFFE_PN0P_  (.CLK(clknet_leaf_189_clk_p2c),
    .RESET_B(net2473),
    .D(_01697_),
    .Q_N(_05270_),
    .Q(\shift_storage.storage[996] ));
 sg13g2_dfrbp_1 \shift_storage.storage[997]$_SDFFE_PN0P_  (.CLK(clknet_leaf_189_clk_p2c),
    .RESET_B(net2474),
    .D(_01698_),
    .Q_N(_05269_),
    .Q(\shift_storage.storage[997] ));
 sg13g2_dfrbp_1 \shift_storage.storage[998]$_SDFFE_PN0P_  (.CLK(clknet_leaf_189_clk_p2c),
    .RESET_B(net2475),
    .D(_01699_),
    .Q_N(_05268_),
    .Q(\shift_storage.storage[998] ));
 sg13g2_dfrbp_1 \shift_storage.storage[999]$_SDFFE_PN0P_  (.CLK(clknet_leaf_198_clk_p2c),
    .RESET_B(net2476),
    .D(_01700_),
    .Q_N(_05267_),
    .Q(\shift_storage.storage[999] ));
 sg13g2_dfrbp_1 \shift_storage.storage[99]$_SDFFE_PN0P_  (.CLK(clknet_leaf_43_clk_p2c),
    .RESET_B(net2477),
    .D(_01701_),
    .Q_N(_05266_),
    .Q(\shift_storage.storage[99] ));
 sg13g2_dfrbp_1 \shift_storage.storage[9]$_SDFFE_PN0P_  (.CLK(clknet_leaf_74_clk_p2c),
    .RESET_B(net2478),
    .D(_01702_),
    .Q_N(_05265_),
    .Q(\shift_storage.storage[9] ));
 sg13g2_IOPadVdd VDD ();
 sg13g2_IOPadIOVdd IOVDD ();
 sg13g2_IOPadVss VSS ();
 sg13g2_IOPadIOVss IOVSS ();
 sg13g2_Corner IO_CORNER_NORTH_WEST_INST ();
 sg13g2_Corner IO_CORNER_NORTH_EAST_INST ();
 sg13g2_Corner IO_CORNER_SOUTH_WEST_INST ();
 sg13g2_Corner IO_CORNER_SOUTH_EAST_INST ();
 sg13g2_Filler200 IO_FILL_IO_NORTH_0_0 ();
 sg13g2_Filler200 IO_FILL_IO_NORTH_0_1 ();
 sg13g2_Filler200 IO_FILL_IO_NORTH_0_2 ();
 sg13g2_Filler200 IO_FILL_IO_NORTH_0_3 ();
 sg13g2_Filler200 IO_FILL_IO_NORTH_0_4 ();
 sg13g2_Filler200 IO_FILL_IO_NORTH_0_5 ();
 sg13g2_Filler200 IO_FILL_IO_NORTH_0_6 ();
 sg13g2_Filler200 IO_FILL_IO_NORTH_0_7 ();
 sg13g2_Filler200 IO_FILL_IO_NORTH_0_8 ();
 sg13g2_Filler200 IO_FILL_IO_NORTH_0_9 ();
 sg13g2_Filler200 IO_FILL_IO_NORTH_1_0 ();
 sg13g2_Filler200 IO_FILL_IO_NORTH_1_1 ();
 sg13g2_Filler200 IO_FILL_IO_NORTH_1_2 ();
 sg13g2_Filler200 IO_FILL_IO_NORTH_1_3 ();
 sg13g2_Filler200 IO_FILL_IO_NORTH_1_4 ();
 sg13g2_Filler200 IO_FILL_IO_NORTH_1_5 ();
 sg13g2_Filler200 IO_FILL_IO_NORTH_1_6 ();
 sg13g2_Filler200 IO_FILL_IO_NORTH_1_7 ();
 sg13g2_Filler200 IO_FILL_IO_NORTH_1_8 ();
 sg13g2_Filler200 IO_FILL_IO_NORTH_1_9 ();
 sg13g2_Filler200 IO_FILL_IO_NORTH_2_0 ();
 sg13g2_Filler200 IO_FILL_IO_NORTH_2_1 ();
 sg13g2_Filler200 IO_FILL_IO_NORTH_2_2 ();
 sg13g2_Filler200 IO_FILL_IO_NORTH_2_3 ();
 sg13g2_Filler200 IO_FILL_IO_NORTH_2_4 ();
 sg13g2_Filler200 IO_FILL_IO_NORTH_2_5 ();
 sg13g2_Filler200 IO_FILL_IO_NORTH_2_6 ();
 sg13g2_Filler200 IO_FILL_IO_NORTH_2_7 ();
 sg13g2_Filler200 IO_FILL_IO_NORTH_2_8 ();
 sg13g2_Filler200 IO_FILL_IO_NORTH_2_9 ();
 sg13g2_Filler200 IO_FILL_IO_NORTH_3_0 ();
 sg13g2_Filler200 IO_FILL_IO_NORTH_3_1 ();
 sg13g2_Filler200 IO_FILL_IO_NORTH_3_2 ();
 sg13g2_Filler200 IO_FILL_IO_NORTH_3_3 ();
 sg13g2_Filler200 IO_FILL_IO_NORTH_3_4 ();
 sg13g2_Filler200 IO_FILL_IO_NORTH_3_5 ();
 sg13g2_Filler200 IO_FILL_IO_NORTH_3_6 ();
 sg13g2_Filler200 IO_FILL_IO_NORTH_3_7 ();
 sg13g2_Filler200 IO_FILL_IO_NORTH_3_8 ();
 sg13g2_Filler200 IO_FILL_IO_NORTH_3_9 ();
 sg13g2_Filler200 IO_FILL_IO_NORTH_4_0 ();
 sg13g2_Filler200 IO_FILL_IO_NORTH_4_1 ();
 sg13g2_Filler200 IO_FILL_IO_NORTH_4_2 ();
 sg13g2_Filler200 IO_FILL_IO_NORTH_4_3 ();
 sg13g2_Filler200 IO_FILL_IO_NORTH_4_4 ();
 sg13g2_Filler200 IO_FILL_IO_NORTH_4_5 ();
 sg13g2_Filler200 IO_FILL_IO_NORTH_4_6 ();
 sg13g2_Filler200 IO_FILL_IO_NORTH_4_7 ();
 sg13g2_Filler200 IO_FILL_IO_NORTH_4_8 ();
 sg13g2_Filler200 IO_FILL_IO_NORTH_4_9 ();
 sg13g2_Filler200 IO_FILL_IO_NORTH_5_0 ();
 sg13g2_Filler200 IO_FILL_IO_NORTH_5_1 ();
 sg13g2_Filler200 IO_FILL_IO_NORTH_5_2 ();
 sg13g2_Filler200 IO_FILL_IO_NORTH_5_3 ();
 sg13g2_Filler200 IO_FILL_IO_NORTH_5_4 ();
 sg13g2_Filler200 IO_FILL_IO_NORTH_5_5 ();
 sg13g2_Filler200 IO_FILL_IO_NORTH_5_6 ();
 sg13g2_Filler200 IO_FILL_IO_NORTH_5_7 ();
 sg13g2_Filler200 IO_FILL_IO_NORTH_5_8 ();
 sg13g2_Filler200 IO_FILL_IO_NORTH_5_9 ();
 sg13g2_Filler200 IO_FILL_IO_NORTH_6_0 ();
 sg13g2_Filler200 IO_FILL_IO_NORTH_6_1 ();
 sg13g2_Filler200 IO_FILL_IO_NORTH_6_2 ();
 sg13g2_Filler200 IO_FILL_IO_NORTH_6_3 ();
 sg13g2_Filler200 IO_FILL_IO_NORTH_6_4 ();
 sg13g2_Filler200 IO_FILL_IO_NORTH_6_5 ();
 sg13g2_Filler200 IO_FILL_IO_NORTH_6_6 ();
 sg13g2_Filler200 IO_FILL_IO_NORTH_6_7 ();
 sg13g2_Filler200 IO_FILL_IO_NORTH_6_8 ();
 sg13g2_Filler200 IO_FILL_IO_NORTH_6_9 ();
 sg13g2_Filler200 IO_FILL_IO_NORTH_7_0 ();
 sg13g2_Filler200 IO_FILL_IO_NORTH_7_1 ();
 sg13g2_Filler200 IO_FILL_IO_NORTH_7_2 ();
 sg13g2_Filler200 IO_FILL_IO_NORTH_7_3 ();
 sg13g2_Filler200 IO_FILL_IO_NORTH_7_4 ();
 sg13g2_Filler200 IO_FILL_IO_NORTH_7_5 ();
 sg13g2_Filler200 IO_FILL_IO_NORTH_7_6 ();
 sg13g2_Filler200 IO_FILL_IO_NORTH_7_7 ();
 sg13g2_Filler200 IO_FILL_IO_NORTH_7_8 ();
 sg13g2_Filler200 IO_FILL_IO_NORTH_7_9 ();
 sg13g2_Filler200 IO_FILL_IO_NORTH_8_0 ();
 sg13g2_Filler200 IO_FILL_IO_NORTH_8_1 ();
 sg13g2_Filler200 IO_FILL_IO_NORTH_8_2 ();
 sg13g2_Filler200 IO_FILL_IO_NORTH_8_3 ();
 sg13g2_Filler200 IO_FILL_IO_NORTH_8_4 ();
 sg13g2_Filler200 IO_FILL_IO_NORTH_8_5 ();
 sg13g2_Filler200 IO_FILL_IO_NORTH_8_6 ();
 sg13g2_Filler200 IO_FILL_IO_NORTH_8_7 ();
 sg13g2_Filler200 IO_FILL_IO_NORTH_8_8 ();
 sg13g2_Filler200 IO_FILL_IO_NORTH_8_9 ();
 sg13g2_Filler200 IO_FILL_IO_SOUTH_0_0 ();
 sg13g2_Filler200 IO_FILL_IO_SOUTH_0_1 ();
 sg13g2_Filler200 IO_FILL_IO_SOUTH_0_2 ();
 sg13g2_Filler200 IO_FILL_IO_SOUTH_0_3 ();
 sg13g2_Filler200 IO_FILL_IO_SOUTH_0_4 ();
 sg13g2_Filler200 IO_FILL_IO_SOUTH_0_5 ();
 sg13g2_Filler200 IO_FILL_IO_SOUTH_0_6 ();
 sg13g2_Filler200 IO_FILL_IO_SOUTH_0_7 ();
 sg13g2_Filler200 IO_FILL_IO_SOUTH_0_8 ();
 sg13g2_Filler200 IO_FILL_IO_SOUTH_0_9 ();
 sg13g2_Filler200 IO_FILL_IO_SOUTH_1_0 ();
 sg13g2_Filler200 IO_FILL_IO_SOUTH_1_1 ();
 sg13g2_Filler200 IO_FILL_IO_SOUTH_1_2 ();
 sg13g2_Filler200 IO_FILL_IO_SOUTH_1_3 ();
 sg13g2_Filler200 IO_FILL_IO_SOUTH_1_4 ();
 sg13g2_Filler200 IO_FILL_IO_SOUTH_1_5 ();
 sg13g2_Filler200 IO_FILL_IO_SOUTH_1_6 ();
 sg13g2_Filler200 IO_FILL_IO_SOUTH_1_7 ();
 sg13g2_Filler200 IO_FILL_IO_SOUTH_1_8 ();
 sg13g2_Filler200 IO_FILL_IO_SOUTH_1_9 ();
 sg13g2_Filler200 IO_FILL_IO_SOUTH_2_0 ();
 sg13g2_Filler200 IO_FILL_IO_SOUTH_2_1 ();
 sg13g2_Filler200 IO_FILL_IO_SOUTH_2_2 ();
 sg13g2_Filler200 IO_FILL_IO_SOUTH_2_3 ();
 sg13g2_Filler200 IO_FILL_IO_SOUTH_2_4 ();
 sg13g2_Filler200 IO_FILL_IO_SOUTH_2_5 ();
 sg13g2_Filler200 IO_FILL_IO_SOUTH_2_6 ();
 sg13g2_Filler200 IO_FILL_IO_SOUTH_2_7 ();
 sg13g2_Filler200 IO_FILL_IO_SOUTH_2_8 ();
 sg13g2_Filler200 IO_FILL_IO_SOUTH_2_9 ();
 sg13g2_Filler200 IO_FILL_IO_SOUTH_3_0 ();
 sg13g2_Filler200 IO_FILL_IO_SOUTH_3_1 ();
 sg13g2_Filler200 IO_FILL_IO_SOUTH_3_2 ();
 sg13g2_Filler200 IO_FILL_IO_SOUTH_3_3 ();
 sg13g2_Filler200 IO_FILL_IO_SOUTH_3_4 ();
 sg13g2_Filler200 IO_FILL_IO_SOUTH_3_5 ();
 sg13g2_Filler200 IO_FILL_IO_SOUTH_3_6 ();
 sg13g2_Filler200 IO_FILL_IO_SOUTH_3_7 ();
 sg13g2_Filler200 IO_FILL_IO_SOUTH_3_8 ();
 sg13g2_Filler200 IO_FILL_IO_SOUTH_3_9 ();
 sg13g2_Filler200 IO_FILL_IO_SOUTH_4_0 ();
 sg13g2_Filler200 IO_FILL_IO_SOUTH_4_1 ();
 sg13g2_Filler200 IO_FILL_IO_SOUTH_4_2 ();
 sg13g2_Filler200 IO_FILL_IO_SOUTH_4_3 ();
 sg13g2_Filler200 IO_FILL_IO_SOUTH_4_4 ();
 sg13g2_Filler200 IO_FILL_IO_SOUTH_4_5 ();
 sg13g2_Filler200 IO_FILL_IO_SOUTH_4_6 ();
 sg13g2_Filler200 IO_FILL_IO_SOUTH_4_7 ();
 sg13g2_Filler200 IO_FILL_IO_SOUTH_4_8 ();
 sg13g2_Filler200 IO_FILL_IO_SOUTH_4_9 ();
 sg13g2_Filler200 IO_FILL_IO_SOUTH_5_0 ();
 sg13g2_Filler200 IO_FILL_IO_SOUTH_5_1 ();
 sg13g2_Filler200 IO_FILL_IO_SOUTH_5_2 ();
 sg13g2_Filler200 IO_FILL_IO_SOUTH_5_3 ();
 sg13g2_Filler200 IO_FILL_IO_SOUTH_5_4 ();
 sg13g2_Filler200 IO_FILL_IO_SOUTH_5_5 ();
 sg13g2_Filler200 IO_FILL_IO_SOUTH_5_6 ();
 sg13g2_Filler200 IO_FILL_IO_SOUTH_5_7 ();
 sg13g2_Filler200 IO_FILL_IO_SOUTH_5_8 ();
 sg13g2_Filler200 IO_FILL_IO_SOUTH_5_9 ();
 sg13g2_Filler200 IO_FILL_IO_SOUTH_6_0 ();
 sg13g2_Filler200 IO_FILL_IO_SOUTH_6_1 ();
 sg13g2_Filler200 IO_FILL_IO_SOUTH_6_2 ();
 sg13g2_Filler200 IO_FILL_IO_SOUTH_6_3 ();
 sg13g2_Filler200 IO_FILL_IO_SOUTH_6_4 ();
 sg13g2_Filler200 IO_FILL_IO_SOUTH_6_5 ();
 sg13g2_Filler200 IO_FILL_IO_SOUTH_6_6 ();
 sg13g2_Filler200 IO_FILL_IO_SOUTH_6_7 ();
 sg13g2_Filler200 IO_FILL_IO_SOUTH_6_8 ();
 sg13g2_Filler200 IO_FILL_IO_SOUTH_6_9 ();
 sg13g2_Filler200 IO_FILL_IO_SOUTH_7_0 ();
 sg13g2_Filler200 IO_FILL_IO_SOUTH_7_1 ();
 sg13g2_Filler200 IO_FILL_IO_SOUTH_7_2 ();
 sg13g2_Filler200 IO_FILL_IO_SOUTH_7_3 ();
 sg13g2_Filler200 IO_FILL_IO_SOUTH_7_4 ();
 sg13g2_Filler200 IO_FILL_IO_SOUTH_7_5 ();
 sg13g2_Filler200 IO_FILL_IO_SOUTH_7_6 ();
 sg13g2_Filler200 IO_FILL_IO_SOUTH_7_7 ();
 sg13g2_Filler200 IO_FILL_IO_SOUTH_7_8 ();
 sg13g2_Filler200 IO_FILL_IO_SOUTH_7_9 ();
 sg13g2_Filler200 IO_FILL_IO_SOUTH_8_0 ();
 sg13g2_Filler200 IO_FILL_IO_SOUTH_8_1 ();
 sg13g2_Filler200 IO_FILL_IO_SOUTH_8_2 ();
 sg13g2_Filler200 IO_FILL_IO_SOUTH_8_3 ();
 sg13g2_Filler200 IO_FILL_IO_SOUTH_8_4 ();
 sg13g2_Filler200 IO_FILL_IO_SOUTH_8_5 ();
 sg13g2_Filler200 IO_FILL_IO_SOUTH_8_6 ();
 sg13g2_Filler200 IO_FILL_IO_SOUTH_8_7 ();
 sg13g2_Filler200 IO_FILL_IO_SOUTH_8_8 ();
 sg13g2_Filler200 IO_FILL_IO_SOUTH_8_9 ();
 sg13g2_Filler200 IO_FILL_IO_WEST_0_0 ();
 sg13g2_Filler200 IO_FILL_IO_WEST_0_1 ();
 sg13g2_Filler200 IO_FILL_IO_WEST_0_2 ();
 sg13g2_Filler200 IO_FILL_IO_WEST_0_3 ();
 sg13g2_Filler200 IO_FILL_IO_WEST_0_4 ();
 sg13g2_Filler200 IO_FILL_IO_WEST_0_5 ();
 sg13g2_Filler200 IO_FILL_IO_WEST_0_6 ();
 sg13g2_Filler200 IO_FILL_IO_WEST_0_7 ();
 sg13g2_Filler200 IO_FILL_IO_WEST_0_8 ();
 sg13g2_Filler200 IO_FILL_IO_WEST_0_9 ();
 sg13g2_Filler200 IO_FILL_IO_WEST_1_0 ();
 sg13g2_Filler200 IO_FILL_IO_WEST_1_1 ();
 sg13g2_Filler200 IO_FILL_IO_WEST_1_2 ();
 sg13g2_Filler200 IO_FILL_IO_WEST_1_3 ();
 sg13g2_Filler200 IO_FILL_IO_WEST_1_4 ();
 sg13g2_Filler200 IO_FILL_IO_WEST_1_5 ();
 sg13g2_Filler200 IO_FILL_IO_WEST_1_6 ();
 sg13g2_Filler200 IO_FILL_IO_WEST_1_7 ();
 sg13g2_Filler200 IO_FILL_IO_WEST_1_8 ();
 sg13g2_Filler200 IO_FILL_IO_WEST_1_9 ();
 sg13g2_Filler200 IO_FILL_IO_WEST_2_0 ();
 sg13g2_Filler200 IO_FILL_IO_WEST_2_1 ();
 sg13g2_Filler200 IO_FILL_IO_WEST_2_2 ();
 sg13g2_Filler200 IO_FILL_IO_WEST_2_3 ();
 sg13g2_Filler200 IO_FILL_IO_WEST_2_4 ();
 sg13g2_Filler200 IO_FILL_IO_WEST_2_5 ();
 sg13g2_Filler200 IO_FILL_IO_WEST_2_6 ();
 sg13g2_Filler200 IO_FILL_IO_WEST_2_7 ();
 sg13g2_Filler200 IO_FILL_IO_WEST_2_8 ();
 sg13g2_Filler200 IO_FILL_IO_WEST_2_9 ();
 sg13g2_Filler200 IO_FILL_IO_WEST_3_0 ();
 sg13g2_Filler200 IO_FILL_IO_WEST_3_1 ();
 sg13g2_Filler200 IO_FILL_IO_WEST_3_2 ();
 sg13g2_Filler200 IO_FILL_IO_WEST_3_3 ();
 sg13g2_Filler200 IO_FILL_IO_WEST_3_4 ();
 sg13g2_Filler200 IO_FILL_IO_WEST_3_5 ();
 sg13g2_Filler200 IO_FILL_IO_WEST_3_6 ();
 sg13g2_Filler200 IO_FILL_IO_WEST_3_7 ();
 sg13g2_Filler200 IO_FILL_IO_WEST_3_8 ();
 sg13g2_Filler200 IO_FILL_IO_WEST_3_9 ();
 sg13g2_Filler200 IO_FILL_IO_WEST_4_0 ();
 sg13g2_Filler200 IO_FILL_IO_WEST_4_1 ();
 sg13g2_Filler200 IO_FILL_IO_WEST_4_2 ();
 sg13g2_Filler200 IO_FILL_IO_WEST_4_3 ();
 sg13g2_Filler200 IO_FILL_IO_WEST_4_4 ();
 sg13g2_Filler200 IO_FILL_IO_WEST_4_5 ();
 sg13g2_Filler200 IO_FILL_IO_WEST_4_6 ();
 sg13g2_Filler200 IO_FILL_IO_WEST_4_7 ();
 sg13g2_Filler200 IO_FILL_IO_WEST_4_8 ();
 sg13g2_Filler200 IO_FILL_IO_WEST_4_9 ();
 sg13g2_Filler200 IO_FILL_IO_WEST_5_0 ();
 sg13g2_Filler200 IO_FILL_IO_WEST_5_1 ();
 sg13g2_Filler200 IO_FILL_IO_WEST_5_2 ();
 sg13g2_Filler200 IO_FILL_IO_WEST_5_3 ();
 sg13g2_Filler200 IO_FILL_IO_WEST_5_4 ();
 sg13g2_Filler200 IO_FILL_IO_WEST_5_5 ();
 sg13g2_Filler200 IO_FILL_IO_WEST_5_6 ();
 sg13g2_Filler200 IO_FILL_IO_WEST_5_7 ();
 sg13g2_Filler200 IO_FILL_IO_WEST_5_8 ();
 sg13g2_Filler200 IO_FILL_IO_WEST_5_9 ();
 sg13g2_Filler200 IO_FILL_IO_WEST_6_0 ();
 sg13g2_Filler200 IO_FILL_IO_WEST_6_1 ();
 sg13g2_Filler200 IO_FILL_IO_WEST_6_2 ();
 sg13g2_Filler200 IO_FILL_IO_WEST_6_3 ();
 sg13g2_Filler200 IO_FILL_IO_WEST_6_4 ();
 sg13g2_Filler200 IO_FILL_IO_WEST_6_5 ();
 sg13g2_Filler200 IO_FILL_IO_WEST_6_6 ();
 sg13g2_Filler200 IO_FILL_IO_WEST_6_7 ();
 sg13g2_Filler200 IO_FILL_IO_WEST_6_8 ();
 sg13g2_Filler200 IO_FILL_IO_WEST_6_9 ();
 sg13g2_Filler200 IO_FILL_IO_WEST_7_0 ();
 sg13g2_Filler200 IO_FILL_IO_WEST_7_1 ();
 sg13g2_Filler200 IO_FILL_IO_WEST_7_2 ();
 sg13g2_Filler200 IO_FILL_IO_WEST_7_3 ();
 sg13g2_Filler200 IO_FILL_IO_WEST_7_4 ();
 sg13g2_Filler200 IO_FILL_IO_WEST_7_5 ();
 sg13g2_Filler200 IO_FILL_IO_WEST_7_6 ();
 sg13g2_Filler200 IO_FILL_IO_WEST_7_7 ();
 sg13g2_Filler200 IO_FILL_IO_WEST_7_8 ();
 sg13g2_Filler200 IO_FILL_IO_WEST_7_9 ();
 sg13g2_Filler200 IO_FILL_IO_WEST_8_0 ();
 sg13g2_Filler200 IO_FILL_IO_WEST_8_1 ();
 sg13g2_Filler200 IO_FILL_IO_WEST_8_2 ();
 sg13g2_Filler200 IO_FILL_IO_WEST_8_3 ();
 sg13g2_Filler200 IO_FILL_IO_WEST_8_4 ();
 sg13g2_Filler200 IO_FILL_IO_WEST_8_5 ();
 sg13g2_Filler200 IO_FILL_IO_WEST_8_6 ();
 sg13g2_Filler200 IO_FILL_IO_WEST_8_7 ();
 sg13g2_Filler200 IO_FILL_IO_WEST_8_8 ();
 sg13g2_Filler200 IO_FILL_IO_WEST_8_9 ();
 sg13g2_Filler200 IO_FILL_IO_EAST_0_0 ();
 sg13g2_Filler200 IO_FILL_IO_EAST_0_1 ();
 sg13g2_Filler200 IO_FILL_IO_EAST_0_2 ();
 sg13g2_Filler200 IO_FILL_IO_EAST_0_3 ();
 sg13g2_Filler200 IO_FILL_IO_EAST_0_4 ();
 sg13g2_Filler200 IO_FILL_IO_EAST_0_5 ();
 sg13g2_Filler200 IO_FILL_IO_EAST_0_6 ();
 sg13g2_Filler200 IO_FILL_IO_EAST_0_7 ();
 sg13g2_Filler200 IO_FILL_IO_EAST_0_8 ();
 sg13g2_Filler200 IO_FILL_IO_EAST_0_9 ();
 sg13g2_Filler200 IO_FILL_IO_EAST_1_0 ();
 sg13g2_Filler200 IO_FILL_IO_EAST_1_1 ();
 sg13g2_Filler200 IO_FILL_IO_EAST_1_2 ();
 sg13g2_Filler200 IO_FILL_IO_EAST_1_3 ();
 sg13g2_Filler200 IO_FILL_IO_EAST_1_4 ();
 sg13g2_Filler200 IO_FILL_IO_EAST_1_5 ();
 sg13g2_Filler200 IO_FILL_IO_EAST_1_6 ();
 sg13g2_Filler200 IO_FILL_IO_EAST_1_7 ();
 sg13g2_Filler200 IO_FILL_IO_EAST_1_8 ();
 sg13g2_Filler200 IO_FILL_IO_EAST_1_9 ();
 sg13g2_Filler200 IO_FILL_IO_EAST_2_0 ();
 sg13g2_Filler200 IO_FILL_IO_EAST_2_1 ();
 sg13g2_Filler200 IO_FILL_IO_EAST_2_2 ();
 sg13g2_Filler200 IO_FILL_IO_EAST_2_3 ();
 sg13g2_Filler200 IO_FILL_IO_EAST_2_4 ();
 sg13g2_Filler200 IO_FILL_IO_EAST_2_5 ();
 sg13g2_Filler200 IO_FILL_IO_EAST_2_6 ();
 sg13g2_Filler200 IO_FILL_IO_EAST_2_7 ();
 sg13g2_Filler200 IO_FILL_IO_EAST_2_8 ();
 sg13g2_Filler200 IO_FILL_IO_EAST_2_9 ();
 sg13g2_Filler200 IO_FILL_IO_EAST_3_0 ();
 sg13g2_Filler200 IO_FILL_IO_EAST_3_1 ();
 sg13g2_Filler200 IO_FILL_IO_EAST_3_2 ();
 sg13g2_Filler200 IO_FILL_IO_EAST_3_3 ();
 sg13g2_Filler200 IO_FILL_IO_EAST_3_4 ();
 sg13g2_Filler200 IO_FILL_IO_EAST_3_5 ();
 sg13g2_Filler200 IO_FILL_IO_EAST_3_6 ();
 sg13g2_Filler200 IO_FILL_IO_EAST_3_7 ();
 sg13g2_Filler200 IO_FILL_IO_EAST_3_8 ();
 sg13g2_Filler200 IO_FILL_IO_EAST_3_9 ();
 sg13g2_Filler200 IO_FILL_IO_EAST_4_0 ();
 sg13g2_Filler200 IO_FILL_IO_EAST_4_1 ();
 sg13g2_Filler200 IO_FILL_IO_EAST_4_2 ();
 sg13g2_Filler200 IO_FILL_IO_EAST_4_3 ();
 sg13g2_Filler200 IO_FILL_IO_EAST_4_4 ();
 sg13g2_Filler200 IO_FILL_IO_EAST_4_5 ();
 sg13g2_Filler200 IO_FILL_IO_EAST_4_6 ();
 sg13g2_Filler200 IO_FILL_IO_EAST_4_7 ();
 sg13g2_Filler200 IO_FILL_IO_EAST_4_8 ();
 sg13g2_Filler200 IO_FILL_IO_EAST_4_9 ();
 sg13g2_Filler200 IO_FILL_IO_EAST_5_0 ();
 sg13g2_Filler200 IO_FILL_IO_EAST_5_1 ();
 sg13g2_Filler200 IO_FILL_IO_EAST_5_2 ();
 sg13g2_Filler200 IO_FILL_IO_EAST_5_3 ();
 sg13g2_Filler200 IO_FILL_IO_EAST_5_4 ();
 sg13g2_Filler200 IO_FILL_IO_EAST_5_5 ();
 sg13g2_Filler200 IO_FILL_IO_EAST_5_6 ();
 sg13g2_Filler200 IO_FILL_IO_EAST_5_7 ();
 sg13g2_Filler200 IO_FILL_IO_EAST_5_8 ();
 sg13g2_Filler200 IO_FILL_IO_EAST_5_9 ();
 sg13g2_Filler200 IO_FILL_IO_EAST_6_0 ();
 sg13g2_Filler200 IO_FILL_IO_EAST_6_1 ();
 sg13g2_Filler200 IO_FILL_IO_EAST_6_2 ();
 sg13g2_Filler200 IO_FILL_IO_EAST_6_3 ();
 sg13g2_Filler200 IO_FILL_IO_EAST_6_4 ();
 sg13g2_Filler200 IO_FILL_IO_EAST_6_5 ();
 sg13g2_Filler200 IO_FILL_IO_EAST_6_6 ();
 sg13g2_Filler200 IO_FILL_IO_EAST_6_7 ();
 sg13g2_Filler200 IO_FILL_IO_EAST_6_8 ();
 sg13g2_Filler200 IO_FILL_IO_EAST_6_9 ();
 sg13g2_Filler200 IO_FILL_IO_EAST_7_0 ();
 sg13g2_Filler200 IO_FILL_IO_EAST_7_1 ();
 sg13g2_Filler200 IO_FILL_IO_EAST_7_2 ();
 sg13g2_Filler200 IO_FILL_IO_EAST_7_3 ();
 sg13g2_Filler200 IO_FILL_IO_EAST_7_4 ();
 sg13g2_Filler200 IO_FILL_IO_EAST_7_5 ();
 sg13g2_Filler200 IO_FILL_IO_EAST_7_6 ();
 sg13g2_Filler200 IO_FILL_IO_EAST_7_7 ();
 sg13g2_Filler200 IO_FILL_IO_EAST_7_8 ();
 sg13g2_Filler200 IO_FILL_IO_EAST_7_9 ();
 sg13g2_Filler200 IO_FILL_IO_EAST_8_0 ();
 sg13g2_Filler200 IO_FILL_IO_EAST_8_1 ();
 sg13g2_Filler200 IO_FILL_IO_EAST_8_2 ();
 sg13g2_Filler200 IO_FILL_IO_EAST_8_3 ();
 sg13g2_Filler200 IO_FILL_IO_EAST_8_4 ();
 sg13g2_Filler200 IO_FILL_IO_EAST_8_5 ();
 sg13g2_Filler200 IO_FILL_IO_EAST_8_6 ();
 sg13g2_Filler200 IO_FILL_IO_EAST_8_7 ();
 sg13g2_Filler200 IO_FILL_IO_EAST_8_8 ();
 sg13g2_Filler200 IO_FILL_IO_EAST_8_9 ();
 bondpad_70x70 IO_BOND_port_aux_enable_cell (.pad(aux_enable_pad));
 bondpad_70x70 IO_BOND_port_clk_cell (.pad(clk_pad));
 bondpad_70x70 IO_BOND_port_data_in1_cell (.pad(data_in_pad[0]));
 bondpad_70x70 IO_BOND_port_data_in2_cell (.pad(data_in_pad[1]));
 bondpad_70x70 IO_BOND_port_data_in3_cell (.pad(data_in_pad[2]));
 bondpad_70x70 IO_BOND_port_data_in4_cell (.pad(data_in_pad[3]));
 bondpad_70x70 IO_BOND_port_data_in5_cell (.pad(data_in_pad[4]));
 bondpad_70x70 IO_BOND_port_data_in6_cell (.pad(data_in_pad[5]));
 bondpad_70x70 IO_BOND_port_data_in7_cell (.pad(data_in_pad[6]));
 bondpad_70x70 IO_BOND_port_data_in8_cell (.pad(data_in_pad[7]));
 bondpad_70x70 IO_BOND_port_data_out1_cell (.pad(data_out_pad[0]));
 bondpad_70x70 IO_BOND_port_data_out2_cell (.pad(data_out_pad[1]));
 bondpad_70x70 IO_BOND_port_data_out3_cell (.pad(data_out_pad[2]));
 bondpad_70x70 IO_BOND_port_data_out4_cell (.pad(data_out_pad[3]));
 bondpad_70x70 IO_BOND_port_data_out5_cell (.pad(data_out_pad[4]));
 bondpad_70x70 IO_BOND_port_data_out6_cell (.pad(data_out_pad[5]));
 bondpad_70x70 IO_BOND_port_data_out7_cell (.pad(data_out_pad[6]));
 bondpad_70x70 IO_BOND_port_data_out8_cell (.pad(data_out_pad[7]));
 bondpad_70x70 IO_BOND_port_lfsr_out_cell (.pad(lfsr_out_pad));
 bondpad_70x70 IO_BOND_port_out_select1_cell (.pad(out_select_pad[0]));
 bondpad_70x70 IO_BOND_port_out_select2_cell (.pad(out_select_pad[1]));
 bondpad_70x70 IO_BOND_port_reg_addr1_cell (.pad(reg_addr_pad[0]));
 bondpad_70x70 IO_BOND_port_reg_addr2_cell (.pad(reg_addr_pad[1]));
 bondpad_70x70 IO_BOND_port_reg_addr3_cell (.pad(reg_addr_pad[2]));
 bondpad_70x70 IO_BOND_port_rst_cell (.pad(rst_pad));
 bondpad_70x70 IO_BOND_port_shreg_in_cell (.pad(shreg_in_pad));
 bondpad_70x70 IO_BOND_port_shreg_out_cell (.pad(shreg_out_pad));
 bondpad_70x70 IO_BOND_port_wr_enable_cell (.pad(wr_enable_pad));
 bondpad_70x70 IO_BOND_VSS (.pad(\IO_CORNER_NORTH_WEST_INST.vss_RING ));
 bondpad_70x70 IO_BOND_VDD (.pad(\IO_CORNER_NORTH_WEST_INST.vdd_RING ));
 bondpad_70x70 IO_BOND_IOVDD (.pad(\IO_CORNER_NORTH_WEST_INST.iovdd_RING ));
 bondpad_70x70 IO_BOND_IOVSS (.pad(\IO_CORNER_NORTH_WEST_INST.iovss_RING ));
 sg13g2_buf_4 fanout609 (.X(net609),
    .A(net611));
 sg13g2_buf_1 fanout610 (.A(net611),
    .X(net610));
 sg13g2_buf_1 fanout611 (.A(net618),
    .X(net611));
 sg13g2_buf_4 fanout612 (.X(net612),
    .A(net613));
 sg13g2_buf_2 fanout613 (.A(net618),
    .X(net613));
 sg13g2_buf_4 fanout614 (.X(net614),
    .A(net615));
 sg13g2_buf_4 fanout615 (.X(net615),
    .A(net616));
 sg13g2_buf_2 fanout616 (.A(net617),
    .X(net616));
 sg13g2_buf_2 fanout617 (.A(net618),
    .X(net617));
 sg13g2_buf_1 fanout618 (.A(net653),
    .X(net618));
 sg13g2_buf_4 fanout619 (.X(net619),
    .A(net624));
 sg13g2_buf_4 fanout620 (.X(net620),
    .A(net624));
 sg13g2_buf_4 fanout621 (.X(net621),
    .A(net623));
 sg13g2_buf_4 fanout622 (.X(net622),
    .A(net624));
 sg13g2_buf_1 fanout623 (.A(net624),
    .X(net623));
 sg13g2_buf_1 fanout624 (.A(net640),
    .X(net624));
 sg13g2_buf_4 fanout625 (.X(net625),
    .A(net626));
 sg13g2_buf_4 fanout626 (.X(net626),
    .A(net629));
 sg13g2_buf_4 fanout627 (.X(net627),
    .A(net629));
 sg13g2_buf_2 fanout628 (.A(net629),
    .X(net628));
 sg13g2_buf_1 fanout629 (.A(net640),
    .X(net629));
 sg13g2_buf_4 fanout630 (.X(net630),
    .A(net634));
 sg13g2_buf_2 fanout631 (.A(net634),
    .X(net631));
 sg13g2_buf_4 fanout632 (.X(net632),
    .A(net634));
 sg13g2_buf_4 fanout633 (.X(net633),
    .A(net634));
 sg13g2_buf_2 fanout634 (.A(net640),
    .X(net634));
 sg13g2_buf_4 fanout635 (.X(net635),
    .A(net636));
 sg13g2_buf_4 fanout636 (.X(net636),
    .A(net639));
 sg13g2_buf_4 fanout637 (.X(net637),
    .A(net639));
 sg13g2_buf_2 fanout638 (.A(net639),
    .X(net638));
 sg13g2_buf_2 fanout639 (.A(net640),
    .X(net639));
 sg13g2_buf_1 fanout640 (.A(net653),
    .X(net640));
 sg13g2_buf_4 fanout641 (.X(net641),
    .A(net644));
 sg13g2_buf_4 fanout642 (.X(net642),
    .A(net643));
 sg13g2_buf_4 fanout643 (.X(net643),
    .A(net644));
 sg13g2_buf_1 fanout644 (.A(net646),
    .X(net644));
 sg13g2_buf_4 fanout645 (.X(net645),
    .A(net646));
 sg13g2_buf_1 fanout646 (.A(net653),
    .X(net646));
 sg13g2_buf_4 fanout647 (.X(net647),
    .A(net648));
 sg13g2_buf_4 fanout648 (.X(net648),
    .A(net652));
 sg13g2_buf_4 fanout649 (.X(net649),
    .A(net651));
 sg13g2_buf_4 fanout650 (.X(net650),
    .A(net651));
 sg13g2_buf_1 fanout651 (.A(net652),
    .X(net651));
 sg13g2_buf_2 fanout652 (.A(net653),
    .X(net652));
 sg13g2_buf_1 fanout653 (.A(net775),
    .X(net653));
 sg13g2_buf_4 fanout654 (.X(net654),
    .A(net655));
 sg13g2_buf_2 fanout655 (.A(net662),
    .X(net655));
 sg13g2_buf_4 fanout656 (.X(net656),
    .A(net662));
 sg13g2_buf_4 fanout657 (.X(net657),
    .A(net661));
 sg13g2_buf_4 fanout658 (.X(net658),
    .A(net661));
 sg13g2_buf_4 fanout659 (.X(net659),
    .A(net661));
 sg13g2_buf_4 fanout660 (.X(net660),
    .A(net661));
 sg13g2_buf_1 fanout661 (.A(net662),
    .X(net661));
 sg13g2_buf_1 fanout662 (.A(net693),
    .X(net662));
 sg13g2_buf_4 fanout663 (.X(net663),
    .A(net666));
 sg13g2_buf_4 fanout664 (.X(net664),
    .A(net665));
 sg13g2_buf_2 fanout665 (.A(net666),
    .X(net665));
 sg13g2_buf_2 fanout666 (.A(net693),
    .X(net666));
 sg13g2_buf_4 fanout667 (.X(net667),
    .A(net668));
 sg13g2_buf_4 fanout668 (.X(net668),
    .A(net671));
 sg13g2_buf_4 fanout669 (.X(net669),
    .A(net671));
 sg13g2_buf_2 fanout670 (.A(net671),
    .X(net670));
 sg13g2_buf_2 fanout671 (.A(net693),
    .X(net671));
 sg13g2_buf_4 fanout672 (.X(net672),
    .A(net673));
 sg13g2_buf_2 fanout673 (.A(net681),
    .X(net673));
 sg13g2_buf_4 fanout674 (.X(net674),
    .A(net675));
 sg13g2_buf_2 fanout675 (.A(net681),
    .X(net675));
 sg13g2_buf_4 fanout676 (.X(net676),
    .A(net677));
 sg13g2_buf_4 fanout677 (.X(net677),
    .A(net680));
 sg13g2_buf_4 fanout678 (.X(net678),
    .A(net679));
 sg13g2_buf_4 fanout679 (.X(net679),
    .A(net680));
 sg13g2_buf_2 fanout680 (.A(net681),
    .X(net680));
 sg13g2_buf_1 fanout681 (.A(net693),
    .X(net681));
 sg13g2_buf_4 fanout682 (.X(net682),
    .A(net686));
 sg13g2_buf_2 fanout683 (.A(net686),
    .X(net683));
 sg13g2_buf_4 fanout684 (.X(net684),
    .A(net686));
 sg13g2_buf_2 fanout685 (.A(net686),
    .X(net685));
 sg13g2_buf_1 fanout686 (.A(net692),
    .X(net686));
 sg13g2_buf_4 fanout687 (.X(net687),
    .A(net688));
 sg13g2_buf_4 fanout688 (.X(net688),
    .A(net692));
 sg13g2_buf_4 fanout689 (.X(net689),
    .A(net691));
 sg13g2_buf_4 fanout690 (.X(net690),
    .A(net691));
 sg13g2_buf_2 fanout691 (.A(net692),
    .X(net691));
 sg13g2_buf_1 fanout692 (.A(net693),
    .X(net692));
 sg13g2_buf_1 fanout693 (.A(net728),
    .X(net693));
 sg13g2_buf_4 fanout694 (.X(net694),
    .A(net695));
 sg13g2_buf_4 fanout695 (.X(net695),
    .A(net712));
 sg13g2_buf_4 fanout696 (.X(net696),
    .A(net697));
 sg13g2_buf_4 fanout697 (.X(net697),
    .A(net700));
 sg13g2_buf_4 fanout698 (.X(net698),
    .A(net699));
 sg13g2_buf_2 fanout699 (.A(net700),
    .X(net699));
 sg13g2_buf_2 fanout700 (.A(net712),
    .X(net700));
 sg13g2_buf_4 fanout701 (.X(net701),
    .A(net702));
 sg13g2_buf_2 fanout702 (.A(net711),
    .X(net702));
 sg13g2_buf_4 fanout703 (.X(net703),
    .A(net705));
 sg13g2_buf_4 fanout704 (.X(net704),
    .A(net705));
 sg13g2_buf_2 fanout705 (.A(net711),
    .X(net705));
 sg13g2_buf_4 fanout706 (.X(net706),
    .A(net710));
 sg13g2_buf_2 fanout707 (.A(net710),
    .X(net707));
 sg13g2_buf_4 fanout708 (.X(net708),
    .A(net709));
 sg13g2_buf_4 fanout709 (.X(net709),
    .A(net710));
 sg13g2_buf_1 fanout710 (.A(net711),
    .X(net710));
 sg13g2_buf_1 fanout711 (.A(net712),
    .X(net711));
 sg13g2_buf_1 fanout712 (.A(net728),
    .X(net712));
 sg13g2_buf_4 fanout713 (.X(net713),
    .A(net715));
 sg13g2_buf_4 fanout714 (.X(net714),
    .A(net715));
 sg13g2_buf_2 fanout715 (.A(net722),
    .X(net715));
 sg13g2_buf_4 fanout716 (.X(net716),
    .A(net722));
 sg13g2_buf_2 fanout717 (.A(net722),
    .X(net717));
 sg13g2_buf_4 fanout718 (.X(net718),
    .A(net721));
 sg13g2_buf_2 fanout719 (.A(net721),
    .X(net719));
 sg13g2_buf_4 fanout720 (.X(net720),
    .A(net721));
 sg13g2_buf_2 fanout721 (.A(net722),
    .X(net721));
 sg13g2_buf_1 fanout722 (.A(net728),
    .X(net722));
 sg13g2_buf_4 fanout723 (.X(net723),
    .A(net724));
 sg13g2_buf_2 fanout724 (.A(net726),
    .X(net724));
 sg13g2_buf_4 fanout725 (.X(net725),
    .A(net726));
 sg13g2_buf_1 fanout726 (.A(net727),
    .X(net726));
 sg13g2_buf_2 fanout727 (.A(net728),
    .X(net727));
 sg13g2_buf_1 fanout728 (.A(net775),
    .X(net728));
 sg13g2_buf_4 fanout729 (.X(net729),
    .A(net730));
 sg13g2_buf_2 fanout730 (.A(net733),
    .X(net730));
 sg13g2_buf_4 fanout731 (.X(net731),
    .A(net733));
 sg13g2_buf_2 fanout732 (.A(net733),
    .X(net732));
 sg13g2_buf_1 fanout733 (.A(net739),
    .X(net733));
 sg13g2_buf_4 fanout734 (.X(net734),
    .A(net736));
 sg13g2_buf_4 fanout735 (.X(net735),
    .A(net736));
 sg13g2_buf_2 fanout736 (.A(net739),
    .X(net736));
 sg13g2_buf_4 fanout737 (.X(net737),
    .A(net739));
 sg13g2_buf_4 fanout738 (.X(net738),
    .A(net739));
 sg13g2_buf_1 fanout739 (.A(net774),
    .X(net739));
 sg13g2_buf_4 fanout740 (.X(net740),
    .A(net744));
 sg13g2_buf_4 fanout741 (.X(net741),
    .A(net744));
 sg13g2_buf_4 fanout742 (.X(net742),
    .A(net743));
 sg13g2_buf_4 fanout743 (.X(net743),
    .A(net744));
 sg13g2_buf_2 fanout744 (.A(net745),
    .X(net744));
 sg13g2_buf_2 fanout745 (.A(net774),
    .X(net745));
 sg13g2_buf_4 fanout746 (.X(net746),
    .A(net749));
 sg13g2_buf_4 fanout747 (.X(net747),
    .A(net748));
 sg13g2_buf_2 fanout748 (.A(net749),
    .X(net748));
 sg13g2_buf_2 fanout749 (.A(net757),
    .X(net749));
 sg13g2_buf_4 fanout750 (.X(net750),
    .A(net751));
 sg13g2_buf_1 fanout751 (.A(net757),
    .X(net751));
 sg13g2_buf_4 fanout752 (.X(net752),
    .A(net754));
 sg13g2_buf_4 fanout753 (.X(net753),
    .A(net754));
 sg13g2_buf_1 fanout754 (.A(net757),
    .X(net754));
 sg13g2_buf_4 fanout755 (.X(net755),
    .A(net756));
 sg13g2_buf_1 fanout756 (.A(net757),
    .X(net756));
 sg13g2_buf_1 fanout757 (.A(net774),
    .X(net757));
 sg13g2_buf_4 fanout758 (.X(net758),
    .A(net759));
 sg13g2_buf_4 fanout759 (.X(net759),
    .A(net762));
 sg13g2_buf_4 fanout760 (.X(net760),
    .A(net761));
 sg13g2_buf_2 fanout761 (.A(net762),
    .X(net761));
 sg13g2_buf_1 fanout762 (.A(net764),
    .X(net762));
 sg13g2_buf_4 fanout763 (.X(net763),
    .A(net764));
 sg13g2_buf_1 fanout764 (.A(net774),
    .X(net764));
 sg13g2_buf_4 fanout765 (.X(net765),
    .A(net767));
 sg13g2_buf_4 fanout766 (.X(net766),
    .A(net767));
 sg13g2_buf_2 fanout767 (.A(net774),
    .X(net767));
 sg13g2_buf_4 fanout768 (.X(net768),
    .A(net773));
 sg13g2_buf_4 fanout769 (.X(net769),
    .A(net770));
 sg13g2_buf_2 fanout770 (.A(net773),
    .X(net770));
 sg13g2_buf_4 fanout771 (.X(net771),
    .A(net773));
 sg13g2_buf_4 fanout772 (.X(net772),
    .A(net773));
 sg13g2_buf_2 fanout773 (.A(net774),
    .X(net773));
 sg13g2_buf_2 fanout774 (.A(net775),
    .X(net774));
 sg13g2_buf_1 fanout775 (.A(aux_enable_p2c),
    .X(net775));
 sg13g2_tiehi \median_processor.input_storage[0]$_SDFFE_PN0P__776  (.L_HI(net776));
 sg13g2_tiehi \median_processor.input_storage[10]$_SDFFE_PN0P__777  (.L_HI(net777));
 sg13g2_tiehi \median_processor.input_storage[11]$_SDFFE_PN0P__778  (.L_HI(net778));
 sg13g2_tiehi \median_processor.input_storage[12]$_SDFFE_PN0P__779  (.L_HI(net779));
 sg13g2_tiehi \median_processor.input_storage[13]$_SDFFE_PN0P__780  (.L_HI(net780));
 sg13g2_tiehi \median_processor.input_storage[14]$_SDFFE_PN0P__781  (.L_HI(net781));
 sg13g2_tiehi \median_processor.input_storage[15]$_SDFFE_PN0P__782  (.L_HI(net782));
 sg13g2_tiehi \median_processor.input_storage[16]$_SDFFE_PN0P__783  (.L_HI(net783));
 sg13g2_tiehi \median_processor.input_storage[17]$_SDFFE_PN0P__784  (.L_HI(net784));
 sg13g2_tiehi \median_processor.input_storage[18]$_SDFFE_PN0P__785  (.L_HI(net785));
 sg13g2_tiehi \median_processor.input_storage[19]$_SDFFE_PN0P__786  (.L_HI(net786));
 sg13g2_tiehi \median_processor.input_storage[1]$_SDFFE_PN0P__787  (.L_HI(net787));
 sg13g2_tiehi \median_processor.input_storage[20]$_SDFFE_PN0P__788  (.L_HI(net788));
 sg13g2_tiehi \median_processor.input_storage[21]$_SDFFE_PN0P__789  (.L_HI(net789));
 sg13g2_tiehi \median_processor.input_storage[22]$_SDFFE_PN0P__790  (.L_HI(net790));
 sg13g2_tiehi \median_processor.input_storage[23]$_SDFFE_PN0P__791  (.L_HI(net791));
 sg13g2_tiehi \median_processor.input_storage[24]$_SDFFE_PN0P__792  (.L_HI(net792));
 sg13g2_tiehi \median_processor.input_storage[25]$_SDFFE_PN0P__793  (.L_HI(net793));
 sg13g2_tiehi \median_processor.input_storage[26]$_SDFFE_PN0P__794  (.L_HI(net794));
 sg13g2_tiehi \median_processor.input_storage[27]$_SDFFE_PN0P__795  (.L_HI(net795));
 sg13g2_tiehi \median_processor.input_storage[28]$_SDFFE_PN0P__796  (.L_HI(net796));
 sg13g2_tiehi \median_processor.input_storage[29]$_SDFFE_PN0P__797  (.L_HI(net797));
 sg13g2_tiehi \median_processor.input_storage[2]$_SDFFE_PN0P__798  (.L_HI(net798));
 sg13g2_tiehi \median_processor.input_storage[30]$_SDFFE_PN0P__799  (.L_HI(net799));
 sg13g2_tiehi \median_processor.input_storage[31]$_SDFFE_PN0P__800  (.L_HI(net800));
 sg13g2_tiehi \median_processor.input_storage[32]$_SDFFE_PN0P__801  (.L_HI(net801));
 sg13g2_tiehi \median_processor.input_storage[33]$_SDFFE_PN0P__802  (.L_HI(net802));
 sg13g2_tiehi \median_processor.input_storage[34]$_SDFFE_PN0P__803  (.L_HI(net803));
 sg13g2_tiehi \median_processor.input_storage[35]$_SDFFE_PN0P__804  (.L_HI(net804));
 sg13g2_tiehi \median_processor.input_storage[36]$_SDFFE_PN0P__805  (.L_HI(net805));
 sg13g2_tiehi \median_processor.input_storage[37]$_SDFFE_PN0P__806  (.L_HI(net806));
 sg13g2_tiehi \median_processor.input_storage[38]$_SDFFE_PN0P__807  (.L_HI(net807));
 sg13g2_tiehi \median_processor.input_storage[39]$_SDFFE_PN0P__808  (.L_HI(net808));
 sg13g2_tiehi \median_processor.input_storage[3]$_SDFFE_PN0P__809  (.L_HI(net809));
 sg13g2_tiehi \median_processor.input_storage[40]$_SDFFE_PN0P__810  (.L_HI(net810));
 sg13g2_tiehi \median_processor.input_storage[41]$_SDFFE_PN0P__811  (.L_HI(net811));
 sg13g2_tiehi \median_processor.input_storage[42]$_SDFFE_PN0P__812  (.L_HI(net812));
 sg13g2_tiehi \median_processor.input_storage[43]$_SDFFE_PN0P__813  (.L_HI(net813));
 sg13g2_tiehi \median_processor.input_storage[44]$_SDFFE_PN0P__814  (.L_HI(net814));
 sg13g2_tiehi \median_processor.input_storage[45]$_SDFFE_PN0P__815  (.L_HI(net815));
 sg13g2_tiehi \median_processor.input_storage[46]$_SDFFE_PN0P__816  (.L_HI(net816));
 sg13g2_tiehi \median_processor.input_storage[47]$_SDFFE_PN0P__817  (.L_HI(net817));
 sg13g2_tiehi \median_processor.input_storage[48]$_SDFFE_PN0P__818  (.L_HI(net818));
 sg13g2_tiehi \median_processor.input_storage[49]$_SDFFE_PN0P__819  (.L_HI(net819));
 sg13g2_tiehi \median_processor.input_storage[4]$_SDFFE_PN0P__820  (.L_HI(net820));
 sg13g2_tiehi \median_processor.input_storage[50]$_SDFFE_PN0P__821  (.L_HI(net821));
 sg13g2_tiehi \median_processor.input_storage[51]$_SDFFE_PN0P__822  (.L_HI(net822));
 sg13g2_tiehi \median_processor.input_storage[52]$_SDFFE_PN0P__823  (.L_HI(net823));
 sg13g2_tiehi \median_processor.input_storage[53]$_SDFFE_PN0P__824  (.L_HI(net824));
 sg13g2_tiehi \median_processor.input_storage[54]$_SDFFE_PN0P__825  (.L_HI(net825));
 sg13g2_tiehi \median_processor.input_storage[55]$_SDFFE_PN0P__826  (.L_HI(net826));
 sg13g2_tiehi \median_processor.input_storage[56]$_SDFFE_PN0P__827  (.L_HI(net827));
 sg13g2_tiehi \median_processor.input_storage[57]$_SDFFE_PN0P__828  (.L_HI(net828));
 sg13g2_tiehi \median_processor.input_storage[58]$_SDFFE_PN0P__829  (.L_HI(net829));
 sg13g2_tiehi \median_processor.input_storage[59]$_SDFFE_PN0P__830  (.L_HI(net830));
 sg13g2_tiehi \median_processor.input_storage[5]$_SDFFE_PN0P__831  (.L_HI(net831));
 sg13g2_tiehi \median_processor.input_storage[60]$_SDFFE_PN0P__832  (.L_HI(net832));
 sg13g2_tiehi \median_processor.input_storage[61]$_SDFFE_PN0P__833  (.L_HI(net833));
 sg13g2_tiehi \median_processor.input_storage[62]$_SDFFE_PN0P__834  (.L_HI(net834));
 sg13g2_tiehi \median_processor.input_storage[63]$_SDFFE_PN0P__835  (.L_HI(net835));
 sg13g2_tiehi \median_processor.input_storage[6]$_SDFFE_PN0P__836  (.L_HI(net836));
 sg13g2_tiehi \median_processor.input_storage[7]$_SDFFE_PN0P__837  (.L_HI(net837));
 sg13g2_tiehi \median_processor.input_storage[8]$_SDFFE_PN0P__838  (.L_HI(net838));
 sg13g2_tiehi \median_processor.input_storage[9]$_SDFFE_PN0P__839  (.L_HI(net839));
 sg13g2_tiehi \median_processor.median_processor.median_out[0]$_DFFE_PP__840  (.L_HI(net840));
 sg13g2_tiehi \median_processor.median_processor.median_out[1]$_DFFE_PP__841  (.L_HI(net841));
 sg13g2_tiehi \median_processor.median_processor.median_out[2]$_DFFE_PP__842  (.L_HI(net842));
 sg13g2_tiehi \median_processor.median_processor.median_out[3]$_DFFE_PP__843  (.L_HI(net843));
 sg13g2_tiehi \median_processor.median_processor.median_out[4]$_DFFE_PP__844  (.L_HI(net844));
 sg13g2_tiehi \median_processor.median_processor.median_out[5]$_DFFE_PP__845  (.L_HI(net845));
 sg13g2_tiehi \median_processor.median_processor.median_out[6]$_DFFE_PP__846  (.L_HI(net846));
 sg13g2_tiehi \median_processor.median_processor.median_out[7]$_DFFE_PP__847  (.L_HI(net847));
 sg13g2_tiehi \rando_generator.lfsr_reg[0]$_SDFF_PN0__848  (.L_HI(net848));
 sg13g2_tiehi \rando_generator.lfsr_reg[10]$_SDFF_PN0__849  (.L_HI(net849));
 sg13g2_tiehi \rando_generator.lfsr_reg[11]$_SDFF_PN0__850  (.L_HI(net850));
 sg13g2_tiehi \rando_generator.lfsr_reg[12]$_SDFF_PN0__851  (.L_HI(net851));
 sg13g2_tiehi \rando_generator.lfsr_reg[13]$_SDFF_PN0__852  (.L_HI(net852));
 sg13g2_tiehi \rando_generator.lfsr_reg[14]$_SDFF_PN0__853  (.L_HI(net853));
 sg13g2_tiehi \rando_generator.lfsr_reg[15]$_SDFF_PN0__854  (.L_HI(net854));
 sg13g2_tiehi \rando_generator.lfsr_reg[16]$_SDFF_PN0__855  (.L_HI(net855));
 sg13g2_tiehi \rando_generator.lfsr_reg[17]$_SDFF_PN0__856  (.L_HI(net856));
 sg13g2_tiehi \rando_generator.lfsr_reg[18]$_SDFF_PN0__857  (.L_HI(net857));
 sg13g2_tiehi \rando_generator.lfsr_reg[19]$_SDFF_PN0__858  (.L_HI(net858));
 sg13g2_tiehi \rando_generator.lfsr_reg[1]$_SDFF_PN0__859  (.L_HI(net859));
 sg13g2_tiehi \rando_generator.lfsr_reg[20]$_SDFF_PN0__860  (.L_HI(net860));
 sg13g2_tiehi \rando_generator.lfsr_reg[21]$_SDFF_PN0__861  (.L_HI(net861));
 sg13g2_tiehi \rando_generator.lfsr_reg[22]$_SDFF_PN0__862  (.L_HI(net862));
 sg13g2_tiehi \rando_generator.lfsr_reg[23]$_SDFF_PN0__863  (.L_HI(net863));
 sg13g2_tiehi \rando_generator.lfsr_reg[24]$_SDFF_PN0__864  (.L_HI(net864));
 sg13g2_tiehi \rando_generator.lfsr_reg[25]$_SDFF_PN0__865  (.L_HI(net865));
 sg13g2_tiehi \rando_generator.lfsr_reg[26]$_SDFF_PN0__866  (.L_HI(net866));
 sg13g2_tiehi \rando_generator.lfsr_reg[27]$_SDFF_PN0__867  (.L_HI(net867));
 sg13g2_tiehi \rando_generator.lfsr_reg[28]$_SDFF_PN0__868  (.L_HI(net868));
 sg13g2_tiehi \rando_generator.lfsr_reg[29]$_SDFF_PN0__869  (.L_HI(net869));
 sg13g2_tiehi \rando_generator.lfsr_reg[2]$_SDFF_PN0__870  (.L_HI(net870));
 sg13g2_tiehi \rando_generator.lfsr_reg[30]$_SDFF_PN0__871  (.L_HI(net871));
 sg13g2_tiehi \rando_generator.lfsr_reg[3]$_SDFF_PN0__872  (.L_HI(net872));
 sg13g2_tiehi \rando_generator.lfsr_reg[4]$_SDFF_PN0__873  (.L_HI(net873));
 sg13g2_tiehi \rando_generator.lfsr_reg[5]$_SDFF_PN0__874  (.L_HI(net874));
 sg13g2_tiehi \rando_generator.lfsr_reg[6]$_SDFF_PN0__875  (.L_HI(net875));
 sg13g2_tiehi \rando_generator.lfsr_reg[7]$_SDFF_PN0__876  (.L_HI(net876));
 sg13g2_tiehi \rando_generator.lfsr_reg[8]$_SDFF_PN0__877  (.L_HI(net877));
 sg13g2_tiehi \rando_generator.lfsr_reg[9]$_SDFF_PN0__878  (.L_HI(net878));
 sg13g2_tiehi \shift_storage.storage[0]$_SDFFE_PN0P__879  (.L_HI(net879));
 sg13g2_tiehi \shift_storage.storage[1000]$_SDFFE_PN0P__880  (.L_HI(net880));
 sg13g2_tiehi \shift_storage.storage[1001]$_SDFFE_PN0P__881  (.L_HI(net881));
 sg13g2_tiehi \shift_storage.storage[1002]$_SDFFE_PN0P__882  (.L_HI(net882));
 sg13g2_tiehi \shift_storage.storage[1003]$_SDFFE_PN0P__883  (.L_HI(net883));
 sg13g2_tiehi \shift_storage.storage[1004]$_SDFFE_PN0P__884  (.L_HI(net884));
 sg13g2_tiehi \shift_storage.storage[1005]$_SDFFE_PN0P__885  (.L_HI(net885));
 sg13g2_tiehi \shift_storage.storage[1006]$_SDFFE_PN0P__886  (.L_HI(net886));
 sg13g2_tiehi \shift_storage.storage[1007]$_SDFFE_PN0P__887  (.L_HI(net887));
 sg13g2_tiehi \shift_storage.storage[1008]$_SDFFE_PN0P__888  (.L_HI(net888));
 sg13g2_tiehi \shift_storage.storage[1009]$_SDFFE_PN0P__889  (.L_HI(net889));
 sg13g2_tiehi \shift_storage.storage[100]$_SDFFE_PN0P__890  (.L_HI(net890));
 sg13g2_tiehi \shift_storage.storage[1010]$_SDFFE_PN0P__891  (.L_HI(net891));
 sg13g2_tiehi \shift_storage.storage[1011]$_SDFFE_PN0P__892  (.L_HI(net892));
 sg13g2_tiehi \shift_storage.storage[1012]$_SDFFE_PN0P__893  (.L_HI(net893));
 sg13g2_tiehi \shift_storage.storage[1013]$_SDFFE_PN0P__894  (.L_HI(net894));
 sg13g2_tiehi \shift_storage.storage[1014]$_SDFFE_PN0P__895  (.L_HI(net895));
 sg13g2_tiehi \shift_storage.storage[1015]$_SDFFE_PN0P__896  (.L_HI(net896));
 sg13g2_tiehi \shift_storage.storage[1016]$_SDFFE_PN0P__897  (.L_HI(net897));
 sg13g2_tiehi \shift_storage.storage[1017]$_SDFFE_PN0P__898  (.L_HI(net898));
 sg13g2_tiehi \shift_storage.storage[1018]$_SDFFE_PN0P__899  (.L_HI(net899));
 sg13g2_tiehi \shift_storage.storage[1019]$_SDFFE_PN0P__900  (.L_HI(net900));
 sg13g2_tiehi \shift_storage.storage[101]$_SDFFE_PN0P__901  (.L_HI(net901));
 sg13g2_tiehi \shift_storage.storage[1020]$_SDFFE_PN0P__902  (.L_HI(net902));
 sg13g2_tiehi \shift_storage.storage[1021]$_SDFFE_PN0P__903  (.L_HI(net903));
 sg13g2_tiehi \shift_storage.storage[1022]$_SDFFE_PN0P__904  (.L_HI(net904));
 sg13g2_tiehi \shift_storage.storage[1023]$_SDFFE_PN0P__905  (.L_HI(net905));
 sg13g2_tiehi \shift_storage.storage[1024]$_SDFFE_PN0P__906  (.L_HI(net906));
 sg13g2_tiehi \shift_storage.storage[1025]$_SDFFE_PN0P__907  (.L_HI(net907));
 sg13g2_tiehi \shift_storage.storage[1026]$_SDFFE_PN0P__908  (.L_HI(net908));
 sg13g2_tiehi \shift_storage.storage[1027]$_SDFFE_PN0P__909  (.L_HI(net909));
 sg13g2_tiehi \shift_storage.storage[1028]$_SDFFE_PN0P__910  (.L_HI(net910));
 sg13g2_tiehi \shift_storage.storage[1029]$_SDFFE_PN0P__911  (.L_HI(net911));
 sg13g2_tiehi \shift_storage.storage[102]$_SDFFE_PN0P__912  (.L_HI(net912));
 sg13g2_tiehi \shift_storage.storage[1030]$_SDFFE_PN0P__913  (.L_HI(net913));
 sg13g2_tiehi \shift_storage.storage[1031]$_SDFFE_PN0P__914  (.L_HI(net914));
 sg13g2_tiehi \shift_storage.storage[1032]$_SDFFE_PN0P__915  (.L_HI(net915));
 sg13g2_tiehi \shift_storage.storage[1033]$_SDFFE_PN0P__916  (.L_HI(net916));
 sg13g2_tiehi \shift_storage.storage[1034]$_SDFFE_PN0P__917  (.L_HI(net917));
 sg13g2_tiehi \shift_storage.storage[1035]$_SDFFE_PN0P__918  (.L_HI(net918));
 sg13g2_tiehi \shift_storage.storage[1036]$_SDFFE_PN0P__919  (.L_HI(net919));
 sg13g2_tiehi \shift_storage.storage[1037]$_SDFFE_PN0P__920  (.L_HI(net920));
 sg13g2_tiehi \shift_storage.storage[1038]$_SDFFE_PN0P__921  (.L_HI(net921));
 sg13g2_tiehi \shift_storage.storage[1039]$_SDFFE_PN0P__922  (.L_HI(net922));
 sg13g2_tiehi \shift_storage.storage[103]$_SDFFE_PN0P__923  (.L_HI(net923));
 sg13g2_tiehi \shift_storage.storage[1040]$_SDFFE_PN0P__924  (.L_HI(net924));
 sg13g2_tiehi \shift_storage.storage[1041]$_SDFFE_PN0P__925  (.L_HI(net925));
 sg13g2_tiehi \shift_storage.storage[1042]$_SDFFE_PN0P__926  (.L_HI(net926));
 sg13g2_tiehi \shift_storage.storage[1043]$_SDFFE_PN0P__927  (.L_HI(net927));
 sg13g2_tiehi \shift_storage.storage[1044]$_SDFFE_PN0P__928  (.L_HI(net928));
 sg13g2_tiehi \shift_storage.storage[1045]$_SDFFE_PN0P__929  (.L_HI(net929));
 sg13g2_tiehi \shift_storage.storage[1046]$_SDFFE_PN0P__930  (.L_HI(net930));
 sg13g2_tiehi \shift_storage.storage[1047]$_SDFFE_PN0P__931  (.L_HI(net931));
 sg13g2_tiehi \shift_storage.storage[1048]$_SDFFE_PN0P__932  (.L_HI(net932));
 sg13g2_tiehi \shift_storage.storage[1049]$_SDFFE_PN0P__933  (.L_HI(net933));
 sg13g2_tiehi \shift_storage.storage[104]$_SDFFE_PN0P__934  (.L_HI(net934));
 sg13g2_tiehi \shift_storage.storage[1050]$_SDFFE_PN0P__935  (.L_HI(net935));
 sg13g2_tiehi \shift_storage.storage[1051]$_SDFFE_PN0P__936  (.L_HI(net936));
 sg13g2_tiehi \shift_storage.storage[1052]$_SDFFE_PN0P__937  (.L_HI(net937));
 sg13g2_tiehi \shift_storage.storage[1053]$_SDFFE_PN0P__938  (.L_HI(net938));
 sg13g2_tiehi \shift_storage.storage[1054]$_SDFFE_PN0P__939  (.L_HI(net939));
 sg13g2_tiehi \shift_storage.storage[1055]$_SDFFE_PN0P__940  (.L_HI(net940));
 sg13g2_tiehi \shift_storage.storage[1056]$_SDFFE_PN0P__941  (.L_HI(net941));
 sg13g2_tiehi \shift_storage.storage[1057]$_SDFFE_PN0P__942  (.L_HI(net942));
 sg13g2_tiehi \shift_storage.storage[1058]$_SDFFE_PN0P__943  (.L_HI(net943));
 sg13g2_tiehi \shift_storage.storage[1059]$_SDFFE_PN0P__944  (.L_HI(net944));
 sg13g2_tiehi \shift_storage.storage[105]$_SDFFE_PN0P__945  (.L_HI(net945));
 sg13g2_tiehi \shift_storage.storage[1060]$_SDFFE_PN0P__946  (.L_HI(net946));
 sg13g2_tiehi \shift_storage.storage[1061]$_SDFFE_PN0P__947  (.L_HI(net947));
 sg13g2_tiehi \shift_storage.storage[1062]$_SDFFE_PN0P__948  (.L_HI(net948));
 sg13g2_tiehi \shift_storage.storage[1063]$_SDFFE_PN0P__949  (.L_HI(net949));
 sg13g2_tiehi \shift_storage.storage[1064]$_SDFFE_PN0P__950  (.L_HI(net950));
 sg13g2_tiehi \shift_storage.storage[1065]$_SDFFE_PN0P__951  (.L_HI(net951));
 sg13g2_tiehi \shift_storage.storage[1066]$_SDFFE_PN0P__952  (.L_HI(net952));
 sg13g2_tiehi \shift_storage.storage[1067]$_SDFFE_PN0P__953  (.L_HI(net953));
 sg13g2_tiehi \shift_storage.storage[1068]$_SDFFE_PN0P__954  (.L_HI(net954));
 sg13g2_tiehi \shift_storage.storage[1069]$_SDFFE_PN0P__955  (.L_HI(net955));
 sg13g2_tiehi \shift_storage.storage[106]$_SDFFE_PN0P__956  (.L_HI(net956));
 sg13g2_tiehi \shift_storage.storage[1070]$_SDFFE_PN0P__957  (.L_HI(net957));
 sg13g2_tiehi \shift_storage.storage[1071]$_SDFFE_PN0P__958  (.L_HI(net958));
 sg13g2_tiehi \shift_storage.storage[1072]$_SDFFE_PN0P__959  (.L_HI(net959));
 sg13g2_tiehi \shift_storage.storage[1073]$_SDFFE_PN0P__960  (.L_HI(net960));
 sg13g2_tiehi \shift_storage.storage[1074]$_SDFFE_PN0P__961  (.L_HI(net961));
 sg13g2_tiehi \shift_storage.storage[1075]$_SDFFE_PN0P__962  (.L_HI(net962));
 sg13g2_tiehi \shift_storage.storage[1076]$_SDFFE_PN0P__963  (.L_HI(net963));
 sg13g2_tiehi \shift_storage.storage[1077]$_SDFFE_PN0P__964  (.L_HI(net964));
 sg13g2_tiehi \shift_storage.storage[1078]$_SDFFE_PN0P__965  (.L_HI(net965));
 sg13g2_tiehi \shift_storage.storage[1079]$_SDFFE_PN0P__966  (.L_HI(net966));
 sg13g2_tiehi \shift_storage.storage[107]$_SDFFE_PN0P__967  (.L_HI(net967));
 sg13g2_tiehi \shift_storage.storage[1080]$_SDFFE_PN0P__968  (.L_HI(net968));
 sg13g2_tiehi \shift_storage.storage[1081]$_SDFFE_PN0P__969  (.L_HI(net969));
 sg13g2_tiehi \shift_storage.storage[1082]$_SDFFE_PN0P__970  (.L_HI(net970));
 sg13g2_tiehi \shift_storage.storage[1083]$_SDFFE_PN0P__971  (.L_HI(net971));
 sg13g2_tiehi \shift_storage.storage[1084]$_SDFFE_PN0P__972  (.L_HI(net972));
 sg13g2_tiehi \shift_storage.storage[1085]$_SDFFE_PN0P__973  (.L_HI(net973));
 sg13g2_tiehi \shift_storage.storage[1086]$_SDFFE_PN0P__974  (.L_HI(net974));
 sg13g2_tiehi \shift_storage.storage[1087]$_SDFFE_PN0P__975  (.L_HI(net975));
 sg13g2_tiehi \shift_storage.storage[1088]$_SDFFE_PN0P__976  (.L_HI(net976));
 sg13g2_tiehi \shift_storage.storage[1089]$_SDFFE_PN0P__977  (.L_HI(net977));
 sg13g2_tiehi \shift_storage.storage[108]$_SDFFE_PN0P__978  (.L_HI(net978));
 sg13g2_tiehi \shift_storage.storage[1090]$_SDFFE_PN0P__979  (.L_HI(net979));
 sg13g2_tiehi \shift_storage.storage[1091]$_SDFFE_PN0P__980  (.L_HI(net980));
 sg13g2_tiehi \shift_storage.storage[1092]$_SDFFE_PN0P__981  (.L_HI(net981));
 sg13g2_tiehi \shift_storage.storage[1093]$_SDFFE_PN0P__982  (.L_HI(net982));
 sg13g2_tiehi \shift_storage.storage[1094]$_SDFFE_PN0P__983  (.L_HI(net983));
 sg13g2_tiehi \shift_storage.storage[1095]$_SDFFE_PN0P__984  (.L_HI(net984));
 sg13g2_tiehi \shift_storage.storage[1096]$_SDFFE_PN0P__985  (.L_HI(net985));
 sg13g2_tiehi \shift_storage.storage[1097]$_SDFFE_PN0P__986  (.L_HI(net986));
 sg13g2_tiehi \shift_storage.storage[1098]$_SDFFE_PN0P__987  (.L_HI(net987));
 sg13g2_tiehi \shift_storage.storage[1099]$_SDFFE_PN0P__988  (.L_HI(net988));
 sg13g2_tiehi \shift_storage.storage[109]$_SDFFE_PN0P__989  (.L_HI(net989));
 sg13g2_tiehi \shift_storage.storage[10]$_SDFFE_PN0P__990  (.L_HI(net990));
 sg13g2_tiehi \shift_storage.storage[1100]$_SDFFE_PN0P__991  (.L_HI(net991));
 sg13g2_tiehi \shift_storage.storage[1101]$_SDFFE_PN0P__992  (.L_HI(net992));
 sg13g2_tiehi \shift_storage.storage[1102]$_SDFFE_PN0P__993  (.L_HI(net993));
 sg13g2_tiehi \shift_storage.storage[1103]$_SDFFE_PN0P__994  (.L_HI(net994));
 sg13g2_tiehi \shift_storage.storage[1104]$_SDFFE_PN0P__995  (.L_HI(net995));
 sg13g2_tiehi \shift_storage.storage[1105]$_SDFFE_PN0P__996  (.L_HI(net996));
 sg13g2_tiehi \shift_storage.storage[1106]$_SDFFE_PN0P__997  (.L_HI(net997));
 sg13g2_tiehi \shift_storage.storage[1107]$_SDFFE_PN0P__998  (.L_HI(net998));
 sg13g2_tiehi \shift_storage.storage[1108]$_SDFFE_PN0P__999  (.L_HI(net999));
 sg13g2_tiehi \shift_storage.storage[1109]$_SDFFE_PN0P__1000  (.L_HI(net1000));
 sg13g2_tiehi \shift_storage.storage[110]$_SDFFE_PN0P__1001  (.L_HI(net1001));
 sg13g2_tiehi \shift_storage.storage[1110]$_SDFFE_PN0P__1002  (.L_HI(net1002));
 sg13g2_tiehi \shift_storage.storage[1111]$_SDFFE_PN0P__1003  (.L_HI(net1003));
 sg13g2_tiehi \shift_storage.storage[1112]$_SDFFE_PN0P__1004  (.L_HI(net1004));
 sg13g2_tiehi \shift_storage.storage[1113]$_SDFFE_PN0P__1005  (.L_HI(net1005));
 sg13g2_tiehi \shift_storage.storage[1114]$_SDFFE_PN0P__1006  (.L_HI(net1006));
 sg13g2_tiehi \shift_storage.storage[1115]$_SDFFE_PN0P__1007  (.L_HI(net1007));
 sg13g2_tiehi \shift_storage.storage[1116]$_SDFFE_PN0P__1008  (.L_HI(net1008));
 sg13g2_tiehi \shift_storage.storage[1117]$_SDFFE_PN0P__1009  (.L_HI(net1009));
 sg13g2_tiehi \shift_storage.storage[1118]$_SDFFE_PN0P__1010  (.L_HI(net1010));
 sg13g2_tiehi \shift_storage.storage[1119]$_SDFFE_PN0P__1011  (.L_HI(net1011));
 sg13g2_tiehi \shift_storage.storage[111]$_SDFFE_PN0P__1012  (.L_HI(net1012));
 sg13g2_tiehi \shift_storage.storage[1120]$_SDFFE_PN0P__1013  (.L_HI(net1013));
 sg13g2_tiehi \shift_storage.storage[1121]$_SDFFE_PN0P__1014  (.L_HI(net1014));
 sg13g2_tiehi \shift_storage.storage[1122]$_SDFFE_PN0P__1015  (.L_HI(net1015));
 sg13g2_tiehi \shift_storage.storage[1123]$_SDFFE_PN0P__1016  (.L_HI(net1016));
 sg13g2_tiehi \shift_storage.storage[1124]$_SDFFE_PN0P__1017  (.L_HI(net1017));
 sg13g2_tiehi \shift_storage.storage[1125]$_SDFFE_PN0P__1018  (.L_HI(net1018));
 sg13g2_tiehi \shift_storage.storage[1126]$_SDFFE_PN0P__1019  (.L_HI(net1019));
 sg13g2_tiehi \shift_storage.storage[1127]$_SDFFE_PN0P__1020  (.L_HI(net1020));
 sg13g2_tiehi \shift_storage.storage[1128]$_SDFFE_PN0P__1021  (.L_HI(net1021));
 sg13g2_tiehi \shift_storage.storage[1129]$_SDFFE_PN0P__1022  (.L_HI(net1022));
 sg13g2_tiehi \shift_storage.storage[112]$_SDFFE_PN0P__1023  (.L_HI(net1023));
 sg13g2_tiehi \shift_storage.storage[1130]$_SDFFE_PN0P__1024  (.L_HI(net1024));
 sg13g2_tiehi \shift_storage.storage[1131]$_SDFFE_PN0P__1025  (.L_HI(net1025));
 sg13g2_tiehi \shift_storage.storage[1132]$_SDFFE_PN0P__1026  (.L_HI(net1026));
 sg13g2_tiehi \shift_storage.storage[1133]$_SDFFE_PN0P__1027  (.L_HI(net1027));
 sg13g2_tiehi \shift_storage.storage[1134]$_SDFFE_PN0P__1028  (.L_HI(net1028));
 sg13g2_tiehi \shift_storage.storage[1135]$_SDFFE_PN0P__1029  (.L_HI(net1029));
 sg13g2_tiehi \shift_storage.storage[1136]$_SDFFE_PN0P__1030  (.L_HI(net1030));
 sg13g2_tiehi \shift_storage.storage[1137]$_SDFFE_PN0P__1031  (.L_HI(net1031));
 sg13g2_tiehi \shift_storage.storage[1138]$_SDFFE_PN0P__1032  (.L_HI(net1032));
 sg13g2_tiehi \shift_storage.storage[1139]$_SDFFE_PN0P__1033  (.L_HI(net1033));
 sg13g2_tiehi \shift_storage.storage[113]$_SDFFE_PN0P__1034  (.L_HI(net1034));
 sg13g2_tiehi \shift_storage.storage[1140]$_SDFFE_PN0P__1035  (.L_HI(net1035));
 sg13g2_tiehi \shift_storage.storage[1141]$_SDFFE_PN0P__1036  (.L_HI(net1036));
 sg13g2_tiehi \shift_storage.storage[1142]$_SDFFE_PN0P__1037  (.L_HI(net1037));
 sg13g2_tiehi \shift_storage.storage[1143]$_SDFFE_PN0P__1038  (.L_HI(net1038));
 sg13g2_tiehi \shift_storage.storage[1144]$_SDFFE_PN0P__1039  (.L_HI(net1039));
 sg13g2_tiehi \shift_storage.storage[1145]$_SDFFE_PN0P__1040  (.L_HI(net1040));
 sg13g2_tiehi \shift_storage.storage[1146]$_SDFFE_PN0P__1041  (.L_HI(net1041));
 sg13g2_tiehi \shift_storage.storage[1147]$_SDFFE_PN0P__1042  (.L_HI(net1042));
 sg13g2_tiehi \shift_storage.storage[1148]$_SDFFE_PN0P__1043  (.L_HI(net1043));
 sg13g2_tiehi \shift_storage.storage[1149]$_SDFFE_PN0P__1044  (.L_HI(net1044));
 sg13g2_tiehi \shift_storage.storage[114]$_SDFFE_PN0P__1045  (.L_HI(net1045));
 sg13g2_tiehi \shift_storage.storage[1150]$_SDFFE_PN0P__1046  (.L_HI(net1046));
 sg13g2_tiehi \shift_storage.storage[1151]$_SDFFE_PN0P__1047  (.L_HI(net1047));
 sg13g2_tiehi \shift_storage.storage[1152]$_SDFFE_PN0P__1048  (.L_HI(net1048));
 sg13g2_tiehi \shift_storage.storage[1153]$_SDFFE_PN0P__1049  (.L_HI(net1049));
 sg13g2_tiehi \shift_storage.storage[1154]$_SDFFE_PN0P__1050  (.L_HI(net1050));
 sg13g2_tiehi \shift_storage.storage[1155]$_SDFFE_PN0P__1051  (.L_HI(net1051));
 sg13g2_tiehi \shift_storage.storage[1156]$_SDFFE_PN0P__1052  (.L_HI(net1052));
 sg13g2_tiehi \shift_storage.storage[1157]$_SDFFE_PN0P__1053  (.L_HI(net1053));
 sg13g2_tiehi \shift_storage.storage[1158]$_SDFFE_PN0P__1054  (.L_HI(net1054));
 sg13g2_tiehi \shift_storage.storage[1159]$_SDFFE_PN0P__1055  (.L_HI(net1055));
 sg13g2_tiehi \shift_storage.storage[115]$_SDFFE_PN0P__1056  (.L_HI(net1056));
 sg13g2_tiehi \shift_storage.storage[1160]$_SDFFE_PN0P__1057  (.L_HI(net1057));
 sg13g2_tiehi \shift_storage.storage[1161]$_SDFFE_PN0P__1058  (.L_HI(net1058));
 sg13g2_tiehi \shift_storage.storage[1162]$_SDFFE_PN0P__1059  (.L_HI(net1059));
 sg13g2_tiehi \shift_storage.storage[1163]$_SDFFE_PN0P__1060  (.L_HI(net1060));
 sg13g2_tiehi \shift_storage.storage[1164]$_SDFFE_PN0P__1061  (.L_HI(net1061));
 sg13g2_tiehi \shift_storage.storage[1165]$_SDFFE_PN0P__1062  (.L_HI(net1062));
 sg13g2_tiehi \shift_storage.storage[1166]$_SDFFE_PN0P__1063  (.L_HI(net1063));
 sg13g2_tiehi \shift_storage.storage[1167]$_SDFFE_PN0P__1064  (.L_HI(net1064));
 sg13g2_tiehi \shift_storage.storage[1168]$_SDFFE_PN0P__1065  (.L_HI(net1065));
 sg13g2_tiehi \shift_storage.storage[1169]$_SDFFE_PN0P__1066  (.L_HI(net1066));
 sg13g2_tiehi \shift_storage.storage[116]$_SDFFE_PN0P__1067  (.L_HI(net1067));
 sg13g2_tiehi \shift_storage.storage[1170]$_SDFFE_PN0P__1068  (.L_HI(net1068));
 sg13g2_tiehi \shift_storage.storage[1171]$_SDFFE_PN0P__1069  (.L_HI(net1069));
 sg13g2_tiehi \shift_storage.storage[1172]$_SDFFE_PN0P__1070  (.L_HI(net1070));
 sg13g2_tiehi \shift_storage.storage[1173]$_SDFFE_PN0P__1071  (.L_HI(net1071));
 sg13g2_tiehi \shift_storage.storage[1174]$_SDFFE_PN0P__1072  (.L_HI(net1072));
 sg13g2_tiehi \shift_storage.storage[1175]$_SDFFE_PN0P__1073  (.L_HI(net1073));
 sg13g2_tiehi \shift_storage.storage[1176]$_SDFFE_PN0P__1074  (.L_HI(net1074));
 sg13g2_tiehi \shift_storage.storage[1177]$_SDFFE_PN0P__1075  (.L_HI(net1075));
 sg13g2_tiehi \shift_storage.storage[1178]$_SDFFE_PN0P__1076  (.L_HI(net1076));
 sg13g2_tiehi \shift_storage.storage[1179]$_SDFFE_PN0P__1077  (.L_HI(net1077));
 sg13g2_tiehi \shift_storage.storage[117]$_SDFFE_PN0P__1078  (.L_HI(net1078));
 sg13g2_tiehi \shift_storage.storage[1180]$_SDFFE_PN0P__1079  (.L_HI(net1079));
 sg13g2_tiehi \shift_storage.storage[1181]$_SDFFE_PN0P__1080  (.L_HI(net1080));
 sg13g2_tiehi \shift_storage.storage[1182]$_SDFFE_PN0P__1081  (.L_HI(net1081));
 sg13g2_tiehi \shift_storage.storage[1183]$_SDFFE_PN0P__1082  (.L_HI(net1082));
 sg13g2_tiehi \shift_storage.storage[1184]$_SDFFE_PN0P__1083  (.L_HI(net1083));
 sg13g2_tiehi \shift_storage.storage[1185]$_SDFFE_PN0P__1084  (.L_HI(net1084));
 sg13g2_tiehi \shift_storage.storage[1186]$_SDFFE_PN0P__1085  (.L_HI(net1085));
 sg13g2_tiehi \shift_storage.storage[1187]$_SDFFE_PN0P__1086  (.L_HI(net1086));
 sg13g2_tiehi \shift_storage.storage[1188]$_SDFFE_PN0P__1087  (.L_HI(net1087));
 sg13g2_tiehi \shift_storage.storage[1189]$_SDFFE_PN0P__1088  (.L_HI(net1088));
 sg13g2_tiehi \shift_storage.storage[118]$_SDFFE_PN0P__1089  (.L_HI(net1089));
 sg13g2_tiehi \shift_storage.storage[1190]$_SDFFE_PN0P__1090  (.L_HI(net1090));
 sg13g2_tiehi \shift_storage.storage[1191]$_SDFFE_PN0P__1091  (.L_HI(net1091));
 sg13g2_tiehi \shift_storage.storage[1192]$_SDFFE_PN0P__1092  (.L_HI(net1092));
 sg13g2_tiehi \shift_storage.storage[1193]$_SDFFE_PN0P__1093  (.L_HI(net1093));
 sg13g2_tiehi \shift_storage.storage[1194]$_SDFFE_PN0P__1094  (.L_HI(net1094));
 sg13g2_tiehi \shift_storage.storage[1195]$_SDFFE_PN0P__1095  (.L_HI(net1095));
 sg13g2_tiehi \shift_storage.storage[1196]$_SDFFE_PN0P__1096  (.L_HI(net1096));
 sg13g2_tiehi \shift_storage.storage[1197]$_SDFFE_PN0P__1097  (.L_HI(net1097));
 sg13g2_tiehi \shift_storage.storage[1198]$_SDFFE_PN0P__1098  (.L_HI(net1098));
 sg13g2_tiehi \shift_storage.storage[1199]$_SDFFE_PN0P__1099  (.L_HI(net1099));
 sg13g2_tiehi \shift_storage.storage[119]$_SDFFE_PN0P__1100  (.L_HI(net1100));
 sg13g2_tiehi \shift_storage.storage[11]$_SDFFE_PN0P__1101  (.L_HI(net1101));
 sg13g2_tiehi \shift_storage.storage[1200]$_SDFFE_PN0P__1102  (.L_HI(net1102));
 sg13g2_tiehi \shift_storage.storage[1201]$_SDFFE_PN0P__1103  (.L_HI(net1103));
 sg13g2_tiehi \shift_storage.storage[1202]$_SDFFE_PN0P__1104  (.L_HI(net1104));
 sg13g2_tiehi \shift_storage.storage[1203]$_SDFFE_PN0P__1105  (.L_HI(net1105));
 sg13g2_tiehi \shift_storage.storage[1204]$_SDFFE_PN0P__1106  (.L_HI(net1106));
 sg13g2_tiehi \shift_storage.storage[1205]$_SDFFE_PN0P__1107  (.L_HI(net1107));
 sg13g2_tiehi \shift_storage.storage[1206]$_SDFFE_PN0P__1108  (.L_HI(net1108));
 sg13g2_tiehi \shift_storage.storage[1207]$_SDFFE_PN0P__1109  (.L_HI(net1109));
 sg13g2_tiehi \shift_storage.storage[1208]$_SDFFE_PN0P__1110  (.L_HI(net1110));
 sg13g2_tiehi \shift_storage.storage[1209]$_SDFFE_PN0P__1111  (.L_HI(net1111));
 sg13g2_tiehi \shift_storage.storage[120]$_SDFFE_PN0P__1112  (.L_HI(net1112));
 sg13g2_tiehi \shift_storage.storage[1210]$_SDFFE_PN0P__1113  (.L_HI(net1113));
 sg13g2_tiehi \shift_storage.storage[1211]$_SDFFE_PN0P__1114  (.L_HI(net1114));
 sg13g2_tiehi \shift_storage.storage[1212]$_SDFFE_PN0P__1115  (.L_HI(net1115));
 sg13g2_tiehi \shift_storage.storage[1213]$_SDFFE_PN0P__1116  (.L_HI(net1116));
 sg13g2_tiehi \shift_storage.storage[1214]$_SDFFE_PN0P__1117  (.L_HI(net1117));
 sg13g2_tiehi \shift_storage.storage[1215]$_SDFFE_PN0P__1118  (.L_HI(net1118));
 sg13g2_tiehi \shift_storage.storage[1216]$_SDFFE_PN0P__1119  (.L_HI(net1119));
 sg13g2_tiehi \shift_storage.storage[1217]$_SDFFE_PN0P__1120  (.L_HI(net1120));
 sg13g2_tiehi \shift_storage.storage[1218]$_SDFFE_PN0P__1121  (.L_HI(net1121));
 sg13g2_tiehi \shift_storage.storage[1219]$_SDFFE_PN0P__1122  (.L_HI(net1122));
 sg13g2_tiehi \shift_storage.storage[121]$_SDFFE_PN0P__1123  (.L_HI(net1123));
 sg13g2_tiehi \shift_storage.storage[1220]$_SDFFE_PN0P__1124  (.L_HI(net1124));
 sg13g2_tiehi \shift_storage.storage[1221]$_SDFFE_PN0P__1125  (.L_HI(net1125));
 sg13g2_tiehi \shift_storage.storage[1222]$_SDFFE_PN0P__1126  (.L_HI(net1126));
 sg13g2_tiehi \shift_storage.storage[1223]$_SDFFE_PN0P__1127  (.L_HI(net1127));
 sg13g2_tiehi \shift_storage.storage[1224]$_SDFFE_PN0P__1128  (.L_HI(net1128));
 sg13g2_tiehi \shift_storage.storage[1225]$_SDFFE_PN0P__1129  (.L_HI(net1129));
 sg13g2_tiehi \shift_storage.storage[1226]$_SDFFE_PN0P__1130  (.L_HI(net1130));
 sg13g2_tiehi \shift_storage.storage[1227]$_SDFFE_PN0P__1131  (.L_HI(net1131));
 sg13g2_tiehi \shift_storage.storage[1228]$_SDFFE_PN0P__1132  (.L_HI(net1132));
 sg13g2_tiehi \shift_storage.storage[1229]$_SDFFE_PN0P__1133  (.L_HI(net1133));
 sg13g2_tiehi \shift_storage.storage[122]$_SDFFE_PN0P__1134  (.L_HI(net1134));
 sg13g2_tiehi \shift_storage.storage[1230]$_SDFFE_PN0P__1135  (.L_HI(net1135));
 sg13g2_tiehi \shift_storage.storage[1231]$_SDFFE_PN0P__1136  (.L_HI(net1136));
 sg13g2_tiehi \shift_storage.storage[1232]$_SDFFE_PN0P__1137  (.L_HI(net1137));
 sg13g2_tiehi \shift_storage.storage[1233]$_SDFFE_PN0P__1138  (.L_HI(net1138));
 sg13g2_tiehi \shift_storage.storage[1234]$_SDFFE_PN0P__1139  (.L_HI(net1139));
 sg13g2_tiehi \shift_storage.storage[1235]$_SDFFE_PN0P__1140  (.L_HI(net1140));
 sg13g2_tiehi \shift_storage.storage[1236]$_SDFFE_PN0P__1141  (.L_HI(net1141));
 sg13g2_tiehi \shift_storage.storage[1237]$_SDFFE_PN0P__1142  (.L_HI(net1142));
 sg13g2_tiehi \shift_storage.storage[1238]$_SDFFE_PN0P__1143  (.L_HI(net1143));
 sg13g2_tiehi \shift_storage.storage[1239]$_SDFFE_PN0P__1144  (.L_HI(net1144));
 sg13g2_tiehi \shift_storage.storage[123]$_SDFFE_PN0P__1145  (.L_HI(net1145));
 sg13g2_tiehi \shift_storage.storage[1240]$_SDFFE_PN0P__1146  (.L_HI(net1146));
 sg13g2_tiehi \shift_storage.storage[1241]$_SDFFE_PN0P__1147  (.L_HI(net1147));
 sg13g2_tiehi \shift_storage.storage[1242]$_SDFFE_PN0P__1148  (.L_HI(net1148));
 sg13g2_tiehi \shift_storage.storage[1243]$_SDFFE_PN0P__1149  (.L_HI(net1149));
 sg13g2_tiehi \shift_storage.storage[1244]$_SDFFE_PN0P__1150  (.L_HI(net1150));
 sg13g2_tiehi \shift_storage.storage[1245]$_SDFFE_PN0P__1151  (.L_HI(net1151));
 sg13g2_tiehi \shift_storage.storage[1246]$_SDFFE_PN0P__1152  (.L_HI(net1152));
 sg13g2_tiehi \shift_storage.storage[1247]$_SDFFE_PN0P__1153  (.L_HI(net1153));
 sg13g2_tiehi \shift_storage.storage[1248]$_SDFFE_PN0P__1154  (.L_HI(net1154));
 sg13g2_tiehi \shift_storage.storage[1249]$_SDFFE_PN0P__1155  (.L_HI(net1155));
 sg13g2_tiehi \shift_storage.storage[124]$_SDFFE_PN0P__1156  (.L_HI(net1156));
 sg13g2_tiehi \shift_storage.storage[1250]$_SDFFE_PN0P__1157  (.L_HI(net1157));
 sg13g2_tiehi \shift_storage.storage[1251]$_SDFFE_PN0P__1158  (.L_HI(net1158));
 sg13g2_tiehi \shift_storage.storage[1252]$_SDFFE_PN0P__1159  (.L_HI(net1159));
 sg13g2_tiehi \shift_storage.storage[1253]$_SDFFE_PN0P__1160  (.L_HI(net1160));
 sg13g2_tiehi \shift_storage.storage[1254]$_SDFFE_PN0P__1161  (.L_HI(net1161));
 sg13g2_tiehi \shift_storage.storage[1255]$_SDFFE_PN0P__1162  (.L_HI(net1162));
 sg13g2_tiehi \shift_storage.storage[1256]$_SDFFE_PN0P__1163  (.L_HI(net1163));
 sg13g2_tiehi \shift_storage.storage[1257]$_SDFFE_PN0P__1164  (.L_HI(net1164));
 sg13g2_tiehi \shift_storage.storage[1258]$_SDFFE_PN0P__1165  (.L_HI(net1165));
 sg13g2_tiehi \shift_storage.storage[1259]$_SDFFE_PN0P__1166  (.L_HI(net1166));
 sg13g2_tiehi \shift_storage.storage[125]$_SDFFE_PN0P__1167  (.L_HI(net1167));
 sg13g2_tiehi \shift_storage.storage[1260]$_SDFFE_PN0P__1168  (.L_HI(net1168));
 sg13g2_tiehi \shift_storage.storage[1261]$_SDFFE_PN0P__1169  (.L_HI(net1169));
 sg13g2_tiehi \shift_storage.storage[1262]$_SDFFE_PN0P__1170  (.L_HI(net1170));
 sg13g2_tiehi \shift_storage.storage[1263]$_SDFFE_PN0P__1171  (.L_HI(net1171));
 sg13g2_tiehi \shift_storage.storage[1264]$_SDFFE_PN0P__1172  (.L_HI(net1172));
 sg13g2_tiehi \shift_storage.storage[1265]$_SDFFE_PN0P__1173  (.L_HI(net1173));
 sg13g2_tiehi \shift_storage.storage[1266]$_SDFFE_PN0P__1174  (.L_HI(net1174));
 sg13g2_tiehi \shift_storage.storage[1267]$_SDFFE_PN0P__1175  (.L_HI(net1175));
 sg13g2_tiehi \shift_storage.storage[1268]$_SDFFE_PN0P__1176  (.L_HI(net1176));
 sg13g2_tiehi \shift_storage.storage[1269]$_SDFFE_PN0P__1177  (.L_HI(net1177));
 sg13g2_tiehi \shift_storage.storage[126]$_SDFFE_PN0P__1178  (.L_HI(net1178));
 sg13g2_tiehi \shift_storage.storage[1270]$_SDFFE_PN0P__1179  (.L_HI(net1179));
 sg13g2_tiehi \shift_storage.storage[1271]$_SDFFE_PN0P__1180  (.L_HI(net1180));
 sg13g2_tiehi \shift_storage.storage[1272]$_SDFFE_PN0P__1181  (.L_HI(net1181));
 sg13g2_tiehi \shift_storage.storage[1273]$_SDFFE_PN0P__1182  (.L_HI(net1182));
 sg13g2_tiehi \shift_storage.storage[1274]$_SDFFE_PN0P__1183  (.L_HI(net1183));
 sg13g2_tiehi \shift_storage.storage[1275]$_SDFFE_PN0P__1184  (.L_HI(net1184));
 sg13g2_tiehi \shift_storage.storage[1276]$_SDFFE_PN0P__1185  (.L_HI(net1185));
 sg13g2_tiehi \shift_storage.storage[1277]$_SDFFE_PN0P__1186  (.L_HI(net1186));
 sg13g2_tiehi \shift_storage.storage[1278]$_SDFFE_PN0P__1187  (.L_HI(net1187));
 sg13g2_tiehi \shift_storage.storage[1279]$_SDFFE_PN0P__1188  (.L_HI(net1188));
 sg13g2_tiehi \shift_storage.storage[127]$_SDFFE_PN0P__1189  (.L_HI(net1189));
 sg13g2_tiehi \shift_storage.storage[1280]$_SDFFE_PN0P__1190  (.L_HI(net1190));
 sg13g2_tiehi \shift_storage.storage[1281]$_SDFFE_PN0P__1191  (.L_HI(net1191));
 sg13g2_tiehi \shift_storage.storage[1282]$_SDFFE_PN0P__1192  (.L_HI(net1192));
 sg13g2_tiehi \shift_storage.storage[1283]$_SDFFE_PN0P__1193  (.L_HI(net1193));
 sg13g2_tiehi \shift_storage.storage[1284]$_SDFFE_PN0P__1194  (.L_HI(net1194));
 sg13g2_tiehi \shift_storage.storage[1285]$_SDFFE_PN0P__1195  (.L_HI(net1195));
 sg13g2_tiehi \shift_storage.storage[1286]$_SDFFE_PN0P__1196  (.L_HI(net1196));
 sg13g2_tiehi \shift_storage.storage[1287]$_SDFFE_PN0P__1197  (.L_HI(net1197));
 sg13g2_tiehi \shift_storage.storage[1288]$_SDFFE_PN0P__1198  (.L_HI(net1198));
 sg13g2_tiehi \shift_storage.storage[1289]$_SDFFE_PN0P__1199  (.L_HI(net1199));
 sg13g2_tiehi \shift_storage.storage[128]$_SDFFE_PN0P__1200  (.L_HI(net1200));
 sg13g2_tiehi \shift_storage.storage[1290]$_SDFFE_PN0P__1201  (.L_HI(net1201));
 sg13g2_tiehi \shift_storage.storage[1291]$_SDFFE_PN0P__1202  (.L_HI(net1202));
 sg13g2_tiehi \shift_storage.storage[1292]$_SDFFE_PN0P__1203  (.L_HI(net1203));
 sg13g2_tiehi \shift_storage.storage[1293]$_SDFFE_PN0P__1204  (.L_HI(net1204));
 sg13g2_tiehi \shift_storage.storage[1294]$_SDFFE_PN0P__1205  (.L_HI(net1205));
 sg13g2_tiehi \shift_storage.storage[1295]$_SDFFE_PN0P__1206  (.L_HI(net1206));
 sg13g2_tiehi \shift_storage.storage[1296]$_SDFFE_PN0P__1207  (.L_HI(net1207));
 sg13g2_tiehi \shift_storage.storage[1297]$_SDFFE_PN0P__1208  (.L_HI(net1208));
 sg13g2_tiehi \shift_storage.storage[1298]$_SDFFE_PN0P__1209  (.L_HI(net1209));
 sg13g2_tiehi \shift_storage.storage[1299]$_SDFFE_PN0P__1210  (.L_HI(net1210));
 sg13g2_tiehi \shift_storage.storage[129]$_SDFFE_PN0P__1211  (.L_HI(net1211));
 sg13g2_tiehi \shift_storage.storage[12]$_SDFFE_PN0P__1212  (.L_HI(net1212));
 sg13g2_tiehi \shift_storage.storage[1300]$_SDFFE_PN0P__1213  (.L_HI(net1213));
 sg13g2_tiehi \shift_storage.storage[1301]$_SDFFE_PN0P__1214  (.L_HI(net1214));
 sg13g2_tiehi \shift_storage.storage[1302]$_SDFFE_PN0P__1215  (.L_HI(net1215));
 sg13g2_tiehi \shift_storage.storage[1303]$_SDFFE_PN0P__1216  (.L_HI(net1216));
 sg13g2_tiehi \shift_storage.storage[1304]$_SDFFE_PN0P__1217  (.L_HI(net1217));
 sg13g2_tiehi \shift_storage.storage[1305]$_SDFFE_PN0P__1218  (.L_HI(net1218));
 sg13g2_tiehi \shift_storage.storage[1306]$_SDFFE_PN0P__1219  (.L_HI(net1219));
 sg13g2_tiehi \shift_storage.storage[1307]$_SDFFE_PN0P__1220  (.L_HI(net1220));
 sg13g2_tiehi \shift_storage.storage[1308]$_SDFFE_PN0P__1221  (.L_HI(net1221));
 sg13g2_tiehi \shift_storage.storage[1309]$_SDFFE_PN0P__1222  (.L_HI(net1222));
 sg13g2_tiehi \shift_storage.storage[130]$_SDFFE_PN0P__1223  (.L_HI(net1223));
 sg13g2_tiehi \shift_storage.storage[1310]$_SDFFE_PN0P__1224  (.L_HI(net1224));
 sg13g2_tiehi \shift_storage.storage[1311]$_SDFFE_PN0P__1225  (.L_HI(net1225));
 sg13g2_tiehi \shift_storage.storage[1312]$_SDFFE_PN0P__1226  (.L_HI(net1226));
 sg13g2_tiehi \shift_storage.storage[1313]$_SDFFE_PN0P__1227  (.L_HI(net1227));
 sg13g2_tiehi \shift_storage.storage[1314]$_SDFFE_PN0P__1228  (.L_HI(net1228));
 sg13g2_tiehi \shift_storage.storage[1315]$_SDFFE_PN0P__1229  (.L_HI(net1229));
 sg13g2_tiehi \shift_storage.storage[1316]$_SDFFE_PN0P__1230  (.L_HI(net1230));
 sg13g2_tiehi \shift_storage.storage[1317]$_SDFFE_PN0P__1231  (.L_HI(net1231));
 sg13g2_tiehi \shift_storage.storage[1318]$_SDFFE_PN0P__1232  (.L_HI(net1232));
 sg13g2_tiehi \shift_storage.storage[1319]$_SDFFE_PN0P__1233  (.L_HI(net1233));
 sg13g2_tiehi \shift_storage.storage[131]$_SDFFE_PN0P__1234  (.L_HI(net1234));
 sg13g2_tiehi \shift_storage.storage[1320]$_SDFFE_PN0P__1235  (.L_HI(net1235));
 sg13g2_tiehi \shift_storage.storage[1321]$_SDFFE_PN0P__1236  (.L_HI(net1236));
 sg13g2_tiehi \shift_storage.storage[1322]$_SDFFE_PN0P__1237  (.L_HI(net1237));
 sg13g2_tiehi \shift_storage.storage[1323]$_SDFFE_PN0P__1238  (.L_HI(net1238));
 sg13g2_tiehi \shift_storage.storage[1324]$_SDFFE_PN0P__1239  (.L_HI(net1239));
 sg13g2_tiehi \shift_storage.storage[1325]$_SDFFE_PN0P__1240  (.L_HI(net1240));
 sg13g2_tiehi \shift_storage.storage[1326]$_SDFFE_PN0P__1241  (.L_HI(net1241));
 sg13g2_tiehi \shift_storage.storage[1327]$_SDFFE_PN0P__1242  (.L_HI(net1242));
 sg13g2_tiehi \shift_storage.storage[1328]$_SDFFE_PN0P__1243  (.L_HI(net1243));
 sg13g2_tiehi \shift_storage.storage[1329]$_SDFFE_PN0P__1244  (.L_HI(net1244));
 sg13g2_tiehi \shift_storage.storage[132]$_SDFFE_PN0P__1245  (.L_HI(net1245));
 sg13g2_tiehi \shift_storage.storage[1330]$_SDFFE_PN0P__1246  (.L_HI(net1246));
 sg13g2_tiehi \shift_storage.storage[1331]$_SDFFE_PN0P__1247  (.L_HI(net1247));
 sg13g2_tiehi \shift_storage.storage[1332]$_SDFFE_PN0P__1248  (.L_HI(net1248));
 sg13g2_tiehi \shift_storage.storage[1333]$_SDFFE_PN0P__1249  (.L_HI(net1249));
 sg13g2_tiehi \shift_storage.storage[1334]$_SDFFE_PN0P__1250  (.L_HI(net1250));
 sg13g2_tiehi \shift_storage.storage[1335]$_SDFFE_PN0P__1251  (.L_HI(net1251));
 sg13g2_tiehi \shift_storage.storage[1336]$_SDFFE_PN0P__1252  (.L_HI(net1252));
 sg13g2_tiehi \shift_storage.storage[1337]$_SDFFE_PN0P__1253  (.L_HI(net1253));
 sg13g2_tiehi \shift_storage.storage[1338]$_SDFFE_PN0P__1254  (.L_HI(net1254));
 sg13g2_tiehi \shift_storage.storage[1339]$_SDFFE_PN0P__1255  (.L_HI(net1255));
 sg13g2_tiehi \shift_storage.storage[133]$_SDFFE_PN0P__1256  (.L_HI(net1256));
 sg13g2_tiehi \shift_storage.storage[1340]$_SDFFE_PN0P__1257  (.L_HI(net1257));
 sg13g2_tiehi \shift_storage.storage[1341]$_SDFFE_PN0P__1258  (.L_HI(net1258));
 sg13g2_tiehi \shift_storage.storage[1342]$_SDFFE_PN0P__1259  (.L_HI(net1259));
 sg13g2_tiehi \shift_storage.storage[1343]$_SDFFE_PN0P__1260  (.L_HI(net1260));
 sg13g2_tiehi \shift_storage.storage[1344]$_SDFFE_PN0P__1261  (.L_HI(net1261));
 sg13g2_tiehi \shift_storage.storage[1345]$_SDFFE_PN0P__1262  (.L_HI(net1262));
 sg13g2_tiehi \shift_storage.storage[1346]$_SDFFE_PN0P__1263  (.L_HI(net1263));
 sg13g2_tiehi \shift_storage.storage[1347]$_SDFFE_PN0P__1264  (.L_HI(net1264));
 sg13g2_tiehi \shift_storage.storage[1348]$_SDFFE_PN0P__1265  (.L_HI(net1265));
 sg13g2_tiehi \shift_storage.storage[1349]$_SDFFE_PN0P__1266  (.L_HI(net1266));
 sg13g2_tiehi \shift_storage.storage[134]$_SDFFE_PN0P__1267  (.L_HI(net1267));
 sg13g2_tiehi \shift_storage.storage[1350]$_SDFFE_PN0P__1268  (.L_HI(net1268));
 sg13g2_tiehi \shift_storage.storage[1351]$_SDFFE_PN0P__1269  (.L_HI(net1269));
 sg13g2_tiehi \shift_storage.storage[1352]$_SDFFE_PN0P__1270  (.L_HI(net1270));
 sg13g2_tiehi \shift_storage.storage[1353]$_SDFFE_PN0P__1271  (.L_HI(net1271));
 sg13g2_tiehi \shift_storage.storage[1354]$_SDFFE_PN0P__1272  (.L_HI(net1272));
 sg13g2_tiehi \shift_storage.storage[1355]$_SDFFE_PN0P__1273  (.L_HI(net1273));
 sg13g2_tiehi \shift_storage.storage[1356]$_SDFFE_PN0P__1274  (.L_HI(net1274));
 sg13g2_tiehi \shift_storage.storage[1357]$_SDFFE_PN0P__1275  (.L_HI(net1275));
 sg13g2_tiehi \shift_storage.storage[1358]$_SDFFE_PN0P__1276  (.L_HI(net1276));
 sg13g2_tiehi \shift_storage.storage[1359]$_SDFFE_PN0P__1277  (.L_HI(net1277));
 sg13g2_tiehi \shift_storage.storage[135]$_SDFFE_PN0P__1278  (.L_HI(net1278));
 sg13g2_tiehi \shift_storage.storage[1360]$_SDFFE_PN0P__1279  (.L_HI(net1279));
 sg13g2_tiehi \shift_storage.storage[1361]$_SDFFE_PN0P__1280  (.L_HI(net1280));
 sg13g2_tiehi \shift_storage.storage[1362]$_SDFFE_PN0P__1281  (.L_HI(net1281));
 sg13g2_tiehi \shift_storage.storage[1363]$_SDFFE_PN0P__1282  (.L_HI(net1282));
 sg13g2_tiehi \shift_storage.storage[1364]$_SDFFE_PN0P__1283  (.L_HI(net1283));
 sg13g2_tiehi \shift_storage.storage[1365]$_SDFFE_PN0P__1284  (.L_HI(net1284));
 sg13g2_tiehi \shift_storage.storage[1366]$_SDFFE_PN0P__1285  (.L_HI(net1285));
 sg13g2_tiehi \shift_storage.storage[1367]$_SDFFE_PN0P__1286  (.L_HI(net1286));
 sg13g2_tiehi \shift_storage.storage[1368]$_SDFFE_PN0P__1287  (.L_HI(net1287));
 sg13g2_tiehi \shift_storage.storage[1369]$_SDFFE_PN0P__1288  (.L_HI(net1288));
 sg13g2_tiehi \shift_storage.storage[136]$_SDFFE_PN0P__1289  (.L_HI(net1289));
 sg13g2_tiehi \shift_storage.storage[1370]$_SDFFE_PN0P__1290  (.L_HI(net1290));
 sg13g2_tiehi \shift_storage.storage[1371]$_SDFFE_PN0P__1291  (.L_HI(net1291));
 sg13g2_tiehi \shift_storage.storage[1372]$_SDFFE_PN0P__1292  (.L_HI(net1292));
 sg13g2_tiehi \shift_storage.storage[1373]$_SDFFE_PN0P__1293  (.L_HI(net1293));
 sg13g2_tiehi \shift_storage.storage[1374]$_SDFFE_PN0P__1294  (.L_HI(net1294));
 sg13g2_tiehi \shift_storage.storage[1375]$_SDFFE_PN0P__1295  (.L_HI(net1295));
 sg13g2_tiehi \shift_storage.storage[1376]$_SDFFE_PN0P__1296  (.L_HI(net1296));
 sg13g2_tiehi \shift_storage.storage[1377]$_SDFFE_PN0P__1297  (.L_HI(net1297));
 sg13g2_tiehi \shift_storage.storage[1378]$_SDFFE_PN0P__1298  (.L_HI(net1298));
 sg13g2_tiehi \shift_storage.storage[1379]$_SDFFE_PN0P__1299  (.L_HI(net1299));
 sg13g2_tiehi \shift_storage.storage[137]$_SDFFE_PN0P__1300  (.L_HI(net1300));
 sg13g2_tiehi \shift_storage.storage[1380]$_SDFFE_PN0P__1301  (.L_HI(net1301));
 sg13g2_tiehi \shift_storage.storage[1381]$_SDFFE_PN0P__1302  (.L_HI(net1302));
 sg13g2_tiehi \shift_storage.storage[1382]$_SDFFE_PN0P__1303  (.L_HI(net1303));
 sg13g2_tiehi \shift_storage.storage[1383]$_SDFFE_PN0P__1304  (.L_HI(net1304));
 sg13g2_tiehi \shift_storage.storage[1384]$_SDFFE_PN0P__1305  (.L_HI(net1305));
 sg13g2_tiehi \shift_storage.storage[1385]$_SDFFE_PN0P__1306  (.L_HI(net1306));
 sg13g2_tiehi \shift_storage.storage[1386]$_SDFFE_PN0P__1307  (.L_HI(net1307));
 sg13g2_tiehi \shift_storage.storage[1387]$_SDFFE_PN0P__1308  (.L_HI(net1308));
 sg13g2_tiehi \shift_storage.storage[1388]$_SDFFE_PN0P__1309  (.L_HI(net1309));
 sg13g2_tiehi \shift_storage.storage[1389]$_SDFFE_PN0P__1310  (.L_HI(net1310));
 sg13g2_tiehi \shift_storage.storage[138]$_SDFFE_PN0P__1311  (.L_HI(net1311));
 sg13g2_tiehi \shift_storage.storage[1390]$_SDFFE_PN0P__1312  (.L_HI(net1312));
 sg13g2_tiehi \shift_storage.storage[1391]$_SDFFE_PN0P__1313  (.L_HI(net1313));
 sg13g2_tiehi \shift_storage.storage[1392]$_SDFFE_PN0P__1314  (.L_HI(net1314));
 sg13g2_tiehi \shift_storage.storage[1393]$_SDFFE_PN0P__1315  (.L_HI(net1315));
 sg13g2_tiehi \shift_storage.storage[1394]$_SDFFE_PN0P__1316  (.L_HI(net1316));
 sg13g2_tiehi \shift_storage.storage[1395]$_SDFFE_PN0P__1317  (.L_HI(net1317));
 sg13g2_tiehi \shift_storage.storage[1396]$_SDFFE_PN0P__1318  (.L_HI(net1318));
 sg13g2_tiehi \shift_storage.storage[1397]$_SDFFE_PN0P__1319  (.L_HI(net1319));
 sg13g2_tiehi \shift_storage.storage[1398]$_SDFFE_PN0P__1320  (.L_HI(net1320));
 sg13g2_tiehi \shift_storage.storage[1399]$_SDFFE_PN0P__1321  (.L_HI(net1321));
 sg13g2_tiehi \shift_storage.storage[139]$_SDFFE_PN0P__1322  (.L_HI(net1322));
 sg13g2_tiehi \shift_storage.storage[13]$_SDFFE_PN0P__1323  (.L_HI(net1323));
 sg13g2_tiehi \shift_storage.storage[1400]$_SDFFE_PN0P__1324  (.L_HI(net1324));
 sg13g2_tiehi \shift_storage.storage[1401]$_SDFFE_PN0P__1325  (.L_HI(net1325));
 sg13g2_tiehi \shift_storage.storage[1402]$_SDFFE_PN0P__1326  (.L_HI(net1326));
 sg13g2_tiehi \shift_storage.storage[1403]$_SDFFE_PN0P__1327  (.L_HI(net1327));
 sg13g2_tiehi \shift_storage.storage[1404]$_SDFFE_PN0P__1328  (.L_HI(net1328));
 sg13g2_tiehi \shift_storage.storage[1405]$_SDFFE_PN0P__1329  (.L_HI(net1329));
 sg13g2_tiehi \shift_storage.storage[1406]$_SDFFE_PN0P__1330  (.L_HI(net1330));
 sg13g2_tiehi \shift_storage.storage[1407]$_SDFFE_PN0P__1331  (.L_HI(net1331));
 sg13g2_tiehi \shift_storage.storage[1408]$_SDFFE_PN0P__1332  (.L_HI(net1332));
 sg13g2_tiehi \shift_storage.storage[1409]$_SDFFE_PN0P__1333  (.L_HI(net1333));
 sg13g2_tiehi \shift_storage.storage[140]$_SDFFE_PN0P__1334  (.L_HI(net1334));
 sg13g2_tiehi \shift_storage.storage[1410]$_SDFFE_PN0P__1335  (.L_HI(net1335));
 sg13g2_tiehi \shift_storage.storage[1411]$_SDFFE_PN0P__1336  (.L_HI(net1336));
 sg13g2_tiehi \shift_storage.storage[1412]$_SDFFE_PN0P__1337  (.L_HI(net1337));
 sg13g2_tiehi \shift_storage.storage[1413]$_SDFFE_PN0P__1338  (.L_HI(net1338));
 sg13g2_tiehi \shift_storage.storage[1414]$_SDFFE_PN0P__1339  (.L_HI(net1339));
 sg13g2_tiehi \shift_storage.storage[1415]$_SDFFE_PN0P__1340  (.L_HI(net1340));
 sg13g2_tiehi \shift_storage.storage[1416]$_SDFFE_PN0P__1341  (.L_HI(net1341));
 sg13g2_tiehi \shift_storage.storage[1417]$_SDFFE_PN0P__1342  (.L_HI(net1342));
 sg13g2_tiehi \shift_storage.storage[1418]$_SDFFE_PN0P__1343  (.L_HI(net1343));
 sg13g2_tiehi \shift_storage.storage[1419]$_SDFFE_PN0P__1344  (.L_HI(net1344));
 sg13g2_tiehi \shift_storage.storage[141]$_SDFFE_PN0P__1345  (.L_HI(net1345));
 sg13g2_tiehi \shift_storage.storage[1420]$_SDFFE_PN0P__1346  (.L_HI(net1346));
 sg13g2_tiehi \shift_storage.storage[1421]$_SDFFE_PN0P__1347  (.L_HI(net1347));
 sg13g2_tiehi \shift_storage.storage[1422]$_SDFFE_PN0P__1348  (.L_HI(net1348));
 sg13g2_tiehi \shift_storage.storage[1423]$_SDFFE_PN0P__1349  (.L_HI(net1349));
 sg13g2_tiehi \shift_storage.storage[1424]$_SDFFE_PN0P__1350  (.L_HI(net1350));
 sg13g2_tiehi \shift_storage.storage[1425]$_SDFFE_PN0P__1351  (.L_HI(net1351));
 sg13g2_tiehi \shift_storage.storage[1426]$_SDFFE_PN0P__1352  (.L_HI(net1352));
 sg13g2_tiehi \shift_storage.storage[1427]$_SDFFE_PN0P__1353  (.L_HI(net1353));
 sg13g2_tiehi \shift_storage.storage[1428]$_SDFFE_PN0P__1354  (.L_HI(net1354));
 sg13g2_tiehi \shift_storage.storage[1429]$_SDFFE_PN0P__1355  (.L_HI(net1355));
 sg13g2_tiehi \shift_storage.storage[142]$_SDFFE_PN0P__1356  (.L_HI(net1356));
 sg13g2_tiehi \shift_storage.storage[1430]$_SDFFE_PN0P__1357  (.L_HI(net1357));
 sg13g2_tiehi \shift_storage.storage[1431]$_SDFFE_PN0P__1358  (.L_HI(net1358));
 sg13g2_tiehi \shift_storage.storage[1432]$_SDFFE_PN0P__1359  (.L_HI(net1359));
 sg13g2_tiehi \shift_storage.storage[1433]$_SDFFE_PN0P__1360  (.L_HI(net1360));
 sg13g2_tiehi \shift_storage.storage[1434]$_SDFFE_PN0P__1361  (.L_HI(net1361));
 sg13g2_tiehi \shift_storage.storage[1435]$_SDFFE_PN0P__1362  (.L_HI(net1362));
 sg13g2_tiehi \shift_storage.storage[1436]$_SDFFE_PN0P__1363  (.L_HI(net1363));
 sg13g2_tiehi \shift_storage.storage[1437]$_SDFFE_PN0P__1364  (.L_HI(net1364));
 sg13g2_tiehi \shift_storage.storage[1438]$_SDFFE_PN0P__1365  (.L_HI(net1365));
 sg13g2_tiehi \shift_storage.storage[1439]$_SDFFE_PN0P__1366  (.L_HI(net1366));
 sg13g2_tiehi \shift_storage.storage[143]$_SDFFE_PN0P__1367  (.L_HI(net1367));
 sg13g2_tiehi \shift_storage.storage[1440]$_SDFFE_PN0P__1368  (.L_HI(net1368));
 sg13g2_tiehi \shift_storage.storage[1441]$_SDFFE_PN0P__1369  (.L_HI(net1369));
 sg13g2_tiehi \shift_storage.storage[1442]$_SDFFE_PN0P__1370  (.L_HI(net1370));
 sg13g2_tiehi \shift_storage.storage[1443]$_SDFFE_PN0P__1371  (.L_HI(net1371));
 sg13g2_tiehi \shift_storage.storage[1444]$_SDFFE_PN0P__1372  (.L_HI(net1372));
 sg13g2_tiehi \shift_storage.storage[1445]$_SDFFE_PN0P__1373  (.L_HI(net1373));
 sg13g2_tiehi \shift_storage.storage[1446]$_SDFFE_PN0P__1374  (.L_HI(net1374));
 sg13g2_tiehi \shift_storage.storage[1447]$_SDFFE_PN0P__1375  (.L_HI(net1375));
 sg13g2_tiehi \shift_storage.storage[1448]$_SDFFE_PN0P__1376  (.L_HI(net1376));
 sg13g2_tiehi \shift_storage.storage[1449]$_SDFFE_PN0P__1377  (.L_HI(net1377));
 sg13g2_tiehi \shift_storage.storage[144]$_SDFFE_PN0P__1378  (.L_HI(net1378));
 sg13g2_tiehi \shift_storage.storage[1450]$_SDFFE_PN0P__1379  (.L_HI(net1379));
 sg13g2_tiehi \shift_storage.storage[1451]$_SDFFE_PN0P__1380  (.L_HI(net1380));
 sg13g2_tiehi \shift_storage.storage[1452]$_SDFFE_PN0P__1381  (.L_HI(net1381));
 sg13g2_tiehi \shift_storage.storage[1453]$_SDFFE_PN0P__1382  (.L_HI(net1382));
 sg13g2_tiehi \shift_storage.storage[1454]$_SDFFE_PN0P__1383  (.L_HI(net1383));
 sg13g2_tiehi \shift_storage.storage[1455]$_SDFFE_PN0P__1384  (.L_HI(net1384));
 sg13g2_tiehi \shift_storage.storage[1456]$_SDFFE_PN0P__1385  (.L_HI(net1385));
 sg13g2_tiehi \shift_storage.storage[1457]$_SDFFE_PN0P__1386  (.L_HI(net1386));
 sg13g2_tiehi \shift_storage.storage[1458]$_SDFFE_PN0P__1387  (.L_HI(net1387));
 sg13g2_tiehi \shift_storage.storage[1459]$_SDFFE_PN0P__1388  (.L_HI(net1388));
 sg13g2_tiehi \shift_storage.storage[145]$_SDFFE_PN0P__1389  (.L_HI(net1389));
 sg13g2_tiehi \shift_storage.storage[1460]$_SDFFE_PN0P__1390  (.L_HI(net1390));
 sg13g2_tiehi \shift_storage.storage[1461]$_SDFFE_PN0P__1391  (.L_HI(net1391));
 sg13g2_tiehi \shift_storage.storage[1462]$_SDFFE_PN0P__1392  (.L_HI(net1392));
 sg13g2_tiehi \shift_storage.storage[1463]$_SDFFE_PN0P__1393  (.L_HI(net1393));
 sg13g2_tiehi \shift_storage.storage[1464]$_SDFFE_PN0P__1394  (.L_HI(net1394));
 sg13g2_tiehi \shift_storage.storage[1465]$_SDFFE_PN0P__1395  (.L_HI(net1395));
 sg13g2_tiehi \shift_storage.storage[1466]$_SDFFE_PN0P__1396  (.L_HI(net1396));
 sg13g2_tiehi \shift_storage.storage[1467]$_SDFFE_PN0P__1397  (.L_HI(net1397));
 sg13g2_tiehi \shift_storage.storage[1468]$_SDFFE_PN0P__1398  (.L_HI(net1398));
 sg13g2_tiehi \shift_storage.storage[1469]$_SDFFE_PN0P__1399  (.L_HI(net1399));
 sg13g2_tiehi \shift_storage.storage[146]$_SDFFE_PN0P__1400  (.L_HI(net1400));
 sg13g2_tiehi \shift_storage.storage[1470]$_SDFFE_PN0P__1401  (.L_HI(net1401));
 sg13g2_tiehi \shift_storage.storage[1471]$_SDFFE_PN0P__1402  (.L_HI(net1402));
 sg13g2_tiehi \shift_storage.storage[1472]$_SDFFE_PN0P__1403  (.L_HI(net1403));
 sg13g2_tiehi \shift_storage.storage[1473]$_SDFFE_PN0P__1404  (.L_HI(net1404));
 sg13g2_tiehi \shift_storage.storage[1474]$_SDFFE_PN0P__1405  (.L_HI(net1405));
 sg13g2_tiehi \shift_storage.storage[1475]$_SDFFE_PN0P__1406  (.L_HI(net1406));
 sg13g2_tiehi \shift_storage.storage[1476]$_SDFFE_PN0P__1407  (.L_HI(net1407));
 sg13g2_tiehi \shift_storage.storage[1477]$_SDFFE_PN0P__1408  (.L_HI(net1408));
 sg13g2_tiehi \shift_storage.storage[1478]$_SDFFE_PN0P__1409  (.L_HI(net1409));
 sg13g2_tiehi \shift_storage.storage[1479]$_SDFFE_PN0P__1410  (.L_HI(net1410));
 sg13g2_tiehi \shift_storage.storage[147]$_SDFFE_PN0P__1411  (.L_HI(net1411));
 sg13g2_tiehi \shift_storage.storage[1480]$_SDFFE_PN0P__1412  (.L_HI(net1412));
 sg13g2_tiehi \shift_storage.storage[1481]$_SDFFE_PN0P__1413  (.L_HI(net1413));
 sg13g2_tiehi \shift_storage.storage[1482]$_SDFFE_PN0P__1414  (.L_HI(net1414));
 sg13g2_tiehi \shift_storage.storage[1483]$_SDFFE_PN0P__1415  (.L_HI(net1415));
 sg13g2_tiehi \shift_storage.storage[1484]$_SDFFE_PN0P__1416  (.L_HI(net1416));
 sg13g2_tiehi \shift_storage.storage[1485]$_SDFFE_PN0P__1417  (.L_HI(net1417));
 sg13g2_tiehi \shift_storage.storage[1486]$_SDFFE_PN0P__1418  (.L_HI(net1418));
 sg13g2_tiehi \shift_storage.storage[1487]$_SDFFE_PN0P__1419  (.L_HI(net1419));
 sg13g2_tiehi \shift_storage.storage[1488]$_SDFFE_PN0P__1420  (.L_HI(net1420));
 sg13g2_tiehi \shift_storage.storage[1489]$_SDFFE_PN0P__1421  (.L_HI(net1421));
 sg13g2_tiehi \shift_storage.storage[148]$_SDFFE_PN0P__1422  (.L_HI(net1422));
 sg13g2_tiehi \shift_storage.storage[1490]$_SDFFE_PN0P__1423  (.L_HI(net1423));
 sg13g2_tiehi \shift_storage.storage[1491]$_SDFFE_PN0P__1424  (.L_HI(net1424));
 sg13g2_tiehi \shift_storage.storage[1492]$_SDFFE_PN0P__1425  (.L_HI(net1425));
 sg13g2_tiehi \shift_storage.storage[1493]$_SDFFE_PN0P__1426  (.L_HI(net1426));
 sg13g2_tiehi \shift_storage.storage[1494]$_SDFFE_PN0P__1427  (.L_HI(net1427));
 sg13g2_tiehi \shift_storage.storage[1495]$_SDFFE_PN0P__1428  (.L_HI(net1428));
 sg13g2_tiehi \shift_storage.storage[1496]$_SDFFE_PN0P__1429  (.L_HI(net1429));
 sg13g2_tiehi \shift_storage.storage[1497]$_SDFFE_PN0P__1430  (.L_HI(net1430));
 sg13g2_tiehi \shift_storage.storage[1498]$_SDFFE_PN0P__1431  (.L_HI(net1431));
 sg13g2_tiehi \shift_storage.storage[1499]$_SDFFE_PN0P__1432  (.L_HI(net1432));
 sg13g2_tiehi \shift_storage.storage[149]$_SDFFE_PN0P__1433  (.L_HI(net1433));
 sg13g2_tiehi \shift_storage.storage[14]$_SDFFE_PN0P__1434  (.L_HI(net1434));
 sg13g2_tiehi \shift_storage.storage[1500]$_SDFFE_PN0P__1435  (.L_HI(net1435));
 sg13g2_tiehi \shift_storage.storage[1501]$_SDFFE_PN0P__1436  (.L_HI(net1436));
 sg13g2_tiehi \shift_storage.storage[1502]$_SDFFE_PN0P__1437  (.L_HI(net1437));
 sg13g2_tiehi \shift_storage.storage[1503]$_SDFFE_PN0P__1438  (.L_HI(net1438));
 sg13g2_tiehi \shift_storage.storage[1504]$_SDFFE_PN0P__1439  (.L_HI(net1439));
 sg13g2_tiehi \shift_storage.storage[1505]$_SDFFE_PN0P__1440  (.L_HI(net1440));
 sg13g2_tiehi \shift_storage.storage[1506]$_SDFFE_PN0P__1441  (.L_HI(net1441));
 sg13g2_tiehi \shift_storage.storage[1507]$_SDFFE_PN0P__1442  (.L_HI(net1442));
 sg13g2_tiehi \shift_storage.storage[1508]$_SDFFE_PN0P__1443  (.L_HI(net1443));
 sg13g2_tiehi \shift_storage.storage[1509]$_SDFFE_PN0P__1444  (.L_HI(net1444));
 sg13g2_tiehi \shift_storage.storage[150]$_SDFFE_PN0P__1445  (.L_HI(net1445));
 sg13g2_tiehi \shift_storage.storage[1510]$_SDFFE_PN0P__1446  (.L_HI(net1446));
 sg13g2_tiehi \shift_storage.storage[1511]$_SDFFE_PN0P__1447  (.L_HI(net1447));
 sg13g2_tiehi \shift_storage.storage[1512]$_SDFFE_PN0P__1448  (.L_HI(net1448));
 sg13g2_tiehi \shift_storage.storage[1513]$_SDFFE_PN0P__1449  (.L_HI(net1449));
 sg13g2_tiehi \shift_storage.storage[1514]$_SDFFE_PN0P__1450  (.L_HI(net1450));
 sg13g2_tiehi \shift_storage.storage[1515]$_SDFFE_PN0P__1451  (.L_HI(net1451));
 sg13g2_tiehi \shift_storage.storage[1516]$_SDFFE_PN0P__1452  (.L_HI(net1452));
 sg13g2_tiehi \shift_storage.storage[1517]$_SDFFE_PN0P__1453  (.L_HI(net1453));
 sg13g2_tiehi \shift_storage.storage[1518]$_SDFFE_PN0P__1454  (.L_HI(net1454));
 sg13g2_tiehi \shift_storage.storage[1519]$_SDFFE_PN0P__1455  (.L_HI(net1455));
 sg13g2_tiehi \shift_storage.storage[151]$_SDFFE_PN0P__1456  (.L_HI(net1456));
 sg13g2_tiehi \shift_storage.storage[1520]$_SDFFE_PN0P__1457  (.L_HI(net1457));
 sg13g2_tiehi \shift_storage.storage[1521]$_SDFFE_PN0P__1458  (.L_HI(net1458));
 sg13g2_tiehi \shift_storage.storage[1522]$_SDFFE_PN0P__1459  (.L_HI(net1459));
 sg13g2_tiehi \shift_storage.storage[1523]$_SDFFE_PN0P__1460  (.L_HI(net1460));
 sg13g2_tiehi \shift_storage.storage[1524]$_SDFFE_PN0P__1461  (.L_HI(net1461));
 sg13g2_tiehi \shift_storage.storage[1525]$_SDFFE_PN0P__1462  (.L_HI(net1462));
 sg13g2_tiehi \shift_storage.storage[1526]$_SDFFE_PN0P__1463  (.L_HI(net1463));
 sg13g2_tiehi \shift_storage.storage[1527]$_SDFFE_PN0P__1464  (.L_HI(net1464));
 sg13g2_tiehi \shift_storage.storage[1528]$_SDFFE_PN0P__1465  (.L_HI(net1465));
 sg13g2_tiehi \shift_storage.storage[1529]$_SDFFE_PN0P__1466  (.L_HI(net1466));
 sg13g2_tiehi \shift_storage.storage[152]$_SDFFE_PN0P__1467  (.L_HI(net1467));
 sg13g2_tiehi \shift_storage.storage[1530]$_SDFFE_PN0P__1468  (.L_HI(net1468));
 sg13g2_tiehi \shift_storage.storage[1531]$_SDFFE_PN0P__1469  (.L_HI(net1469));
 sg13g2_tiehi \shift_storage.storage[1532]$_SDFFE_PN0P__1470  (.L_HI(net1470));
 sg13g2_tiehi \shift_storage.storage[1533]$_SDFFE_PN0P__1471  (.L_HI(net1471));
 sg13g2_tiehi \shift_storage.storage[1534]$_SDFFE_PN0P__1472  (.L_HI(net1472));
 sg13g2_tiehi \shift_storage.storage[1535]$_SDFFE_PN0P__1473  (.L_HI(net1473));
 sg13g2_tiehi \shift_storage.storage[1536]$_SDFFE_PN0P__1474  (.L_HI(net1474));
 sg13g2_tiehi \shift_storage.storage[1537]$_SDFFE_PN0P__1475  (.L_HI(net1475));
 sg13g2_tiehi \shift_storage.storage[1538]$_SDFFE_PN0P__1476  (.L_HI(net1476));
 sg13g2_tiehi \shift_storage.storage[1539]$_SDFFE_PN0P__1477  (.L_HI(net1477));
 sg13g2_tiehi \shift_storage.storage[153]$_SDFFE_PN0P__1478  (.L_HI(net1478));
 sg13g2_tiehi \shift_storage.storage[1540]$_SDFFE_PN0P__1479  (.L_HI(net1479));
 sg13g2_tiehi \shift_storage.storage[1541]$_SDFFE_PN0P__1480  (.L_HI(net1480));
 sg13g2_tiehi \shift_storage.storage[1542]$_SDFFE_PN0P__1481  (.L_HI(net1481));
 sg13g2_tiehi \shift_storage.storage[1543]$_SDFFE_PN0P__1482  (.L_HI(net1482));
 sg13g2_tiehi \shift_storage.storage[1544]$_SDFFE_PN0P__1483  (.L_HI(net1483));
 sg13g2_tiehi \shift_storage.storage[1545]$_SDFFE_PN0P__1484  (.L_HI(net1484));
 sg13g2_tiehi \shift_storage.storage[1546]$_SDFFE_PN0P__1485  (.L_HI(net1485));
 sg13g2_tiehi \shift_storage.storage[1547]$_SDFFE_PN0P__1486  (.L_HI(net1486));
 sg13g2_tiehi \shift_storage.storage[1548]$_SDFFE_PN0P__1487  (.L_HI(net1487));
 sg13g2_tiehi \shift_storage.storage[1549]$_SDFFE_PN0P__1488  (.L_HI(net1488));
 sg13g2_tiehi \shift_storage.storage[154]$_SDFFE_PN0P__1489  (.L_HI(net1489));
 sg13g2_tiehi \shift_storage.storage[1550]$_SDFFE_PN0P__1490  (.L_HI(net1490));
 sg13g2_tiehi \shift_storage.storage[1551]$_SDFFE_PN0P__1491  (.L_HI(net1491));
 sg13g2_tiehi \shift_storage.storage[1552]$_SDFFE_PN0P__1492  (.L_HI(net1492));
 sg13g2_tiehi \shift_storage.storage[1553]$_SDFFE_PN0P__1493  (.L_HI(net1493));
 sg13g2_tiehi \shift_storage.storage[1554]$_SDFFE_PN0P__1494  (.L_HI(net1494));
 sg13g2_tiehi \shift_storage.storage[1555]$_SDFFE_PN0P__1495  (.L_HI(net1495));
 sg13g2_tiehi \shift_storage.storage[1556]$_SDFFE_PN0P__1496  (.L_HI(net1496));
 sg13g2_tiehi \shift_storage.storage[1557]$_SDFFE_PN0P__1497  (.L_HI(net1497));
 sg13g2_tiehi \shift_storage.storage[1558]$_SDFFE_PN0P__1498  (.L_HI(net1498));
 sg13g2_tiehi \shift_storage.storage[1559]$_SDFFE_PN0P__1499  (.L_HI(net1499));
 sg13g2_tiehi \shift_storage.storage[155]$_SDFFE_PN0P__1500  (.L_HI(net1500));
 sg13g2_tiehi \shift_storage.storage[1560]$_SDFFE_PN0P__1501  (.L_HI(net1501));
 sg13g2_tiehi \shift_storage.storage[1561]$_SDFFE_PN0P__1502  (.L_HI(net1502));
 sg13g2_tiehi \shift_storage.storage[1562]$_SDFFE_PN0P__1503  (.L_HI(net1503));
 sg13g2_tiehi \shift_storage.storage[1563]$_SDFFE_PN0P__1504  (.L_HI(net1504));
 sg13g2_tiehi \shift_storage.storage[1564]$_SDFFE_PN0P__1505  (.L_HI(net1505));
 sg13g2_tiehi \shift_storage.storage[1565]$_SDFFE_PN0P__1506  (.L_HI(net1506));
 sg13g2_tiehi \shift_storage.storage[1566]$_SDFFE_PN0P__1507  (.L_HI(net1507));
 sg13g2_tiehi \shift_storage.storage[1567]$_SDFFE_PN0P__1508  (.L_HI(net1508));
 sg13g2_tiehi \shift_storage.storage[1568]$_SDFFE_PN0P__1509  (.L_HI(net1509));
 sg13g2_tiehi \shift_storage.storage[1569]$_SDFFE_PN0P__1510  (.L_HI(net1510));
 sg13g2_tiehi \shift_storage.storage[156]$_SDFFE_PN0P__1511  (.L_HI(net1511));
 sg13g2_tiehi \shift_storage.storage[1570]$_SDFFE_PN0P__1512  (.L_HI(net1512));
 sg13g2_tiehi \shift_storage.storage[1571]$_SDFFE_PN0P__1513  (.L_HI(net1513));
 sg13g2_tiehi \shift_storage.storage[1572]$_SDFFE_PN0P__1514  (.L_HI(net1514));
 sg13g2_tiehi \shift_storage.storage[1573]$_SDFFE_PN0P__1515  (.L_HI(net1515));
 sg13g2_tiehi \shift_storage.storage[1574]$_SDFFE_PN0P__1516  (.L_HI(net1516));
 sg13g2_tiehi \shift_storage.storage[1575]$_SDFFE_PN0P__1517  (.L_HI(net1517));
 sg13g2_tiehi \shift_storage.storage[1576]$_SDFFE_PN0P__1518  (.L_HI(net1518));
 sg13g2_tiehi \shift_storage.storage[1577]$_SDFFE_PN0P__1519  (.L_HI(net1519));
 sg13g2_tiehi \shift_storage.storage[1578]$_SDFFE_PN0P__1520  (.L_HI(net1520));
 sg13g2_tiehi \shift_storage.storage[1579]$_SDFFE_PN0P__1521  (.L_HI(net1521));
 sg13g2_tiehi \shift_storage.storage[157]$_SDFFE_PN0P__1522  (.L_HI(net1522));
 sg13g2_tiehi \shift_storage.storage[1580]$_SDFFE_PN0P__1523  (.L_HI(net1523));
 sg13g2_tiehi \shift_storage.storage[1581]$_SDFFE_PN0P__1524  (.L_HI(net1524));
 sg13g2_tiehi \shift_storage.storage[1582]$_SDFFE_PN0P__1525  (.L_HI(net1525));
 sg13g2_tiehi \shift_storage.storage[1583]$_SDFFE_PN0P__1526  (.L_HI(net1526));
 sg13g2_tiehi \shift_storage.storage[1584]$_SDFFE_PN0P__1527  (.L_HI(net1527));
 sg13g2_tiehi \shift_storage.storage[1585]$_SDFFE_PN0P__1528  (.L_HI(net1528));
 sg13g2_tiehi \shift_storage.storage[1586]$_SDFFE_PN0P__1529  (.L_HI(net1529));
 sg13g2_tiehi \shift_storage.storage[1587]$_SDFFE_PN0P__1530  (.L_HI(net1530));
 sg13g2_tiehi \shift_storage.storage[1588]$_SDFFE_PN0P__1531  (.L_HI(net1531));
 sg13g2_tiehi \shift_storage.storage[1589]$_SDFFE_PN0P__1532  (.L_HI(net1532));
 sg13g2_tiehi \shift_storage.storage[158]$_SDFFE_PN0P__1533  (.L_HI(net1533));
 sg13g2_tiehi \shift_storage.storage[1590]$_SDFFE_PN0P__1534  (.L_HI(net1534));
 sg13g2_tiehi \shift_storage.storage[1591]$_SDFFE_PN0P__1535  (.L_HI(net1535));
 sg13g2_tiehi \shift_storage.storage[1592]$_SDFFE_PN0P__1536  (.L_HI(net1536));
 sg13g2_tiehi \shift_storage.storage[1593]$_SDFFE_PN0P__1537  (.L_HI(net1537));
 sg13g2_tiehi \shift_storage.storage[1594]$_SDFFE_PN0P__1538  (.L_HI(net1538));
 sg13g2_tiehi \shift_storage.storage[1595]$_SDFFE_PN0P__1539  (.L_HI(net1539));
 sg13g2_tiehi \shift_storage.storage[1596]$_SDFFE_PN0P__1540  (.L_HI(net1540));
 sg13g2_tiehi \shift_storage.storage[1597]$_SDFFE_PN0P__1541  (.L_HI(net1541));
 sg13g2_tiehi \shift_storage.storage[1598]$_SDFFE_PN0P__1542  (.L_HI(net1542));
 sg13g2_tiehi \shift_storage.storage[1599]$_SDFFE_PN0P__1543  (.L_HI(net1543));
 sg13g2_tiehi \shift_storage.storage[159]$_SDFFE_PN0P__1544  (.L_HI(net1544));
 sg13g2_tiehi \shift_storage.storage[15]$_SDFFE_PN0P__1545  (.L_HI(net1545));
 sg13g2_tiehi \shift_storage.storage[160]$_SDFFE_PN0P__1546  (.L_HI(net1546));
 sg13g2_tiehi \shift_storage.storage[161]$_SDFFE_PN0P__1547  (.L_HI(net1547));
 sg13g2_tiehi \shift_storage.storage[162]$_SDFFE_PN0P__1548  (.L_HI(net1548));
 sg13g2_tiehi \shift_storage.storage[163]$_SDFFE_PN0P__1549  (.L_HI(net1549));
 sg13g2_tiehi \shift_storage.storage[164]$_SDFFE_PN0P__1550  (.L_HI(net1550));
 sg13g2_tiehi \shift_storage.storage[165]$_SDFFE_PN0P__1551  (.L_HI(net1551));
 sg13g2_tiehi \shift_storage.storage[166]$_SDFFE_PN0P__1552  (.L_HI(net1552));
 sg13g2_tiehi \shift_storage.storage[167]$_SDFFE_PN0P__1553  (.L_HI(net1553));
 sg13g2_tiehi \shift_storage.storage[168]$_SDFFE_PN0P__1554  (.L_HI(net1554));
 sg13g2_tiehi \shift_storage.storage[169]$_SDFFE_PN0P__1555  (.L_HI(net1555));
 sg13g2_tiehi \shift_storage.storage[16]$_SDFFE_PN0P__1556  (.L_HI(net1556));
 sg13g2_tiehi \shift_storage.storage[170]$_SDFFE_PN0P__1557  (.L_HI(net1557));
 sg13g2_tiehi \shift_storage.storage[171]$_SDFFE_PN0P__1558  (.L_HI(net1558));
 sg13g2_tiehi \shift_storage.storage[172]$_SDFFE_PN0P__1559  (.L_HI(net1559));
 sg13g2_tiehi \shift_storage.storage[173]$_SDFFE_PN0P__1560  (.L_HI(net1560));
 sg13g2_tiehi \shift_storage.storage[174]$_SDFFE_PN0P__1561  (.L_HI(net1561));
 sg13g2_tiehi \shift_storage.storage[175]$_SDFFE_PN0P__1562  (.L_HI(net1562));
 sg13g2_tiehi \shift_storage.storage[176]$_SDFFE_PN0P__1563  (.L_HI(net1563));
 sg13g2_tiehi \shift_storage.storage[177]$_SDFFE_PN0P__1564  (.L_HI(net1564));
 sg13g2_tiehi \shift_storage.storage[178]$_SDFFE_PN0P__1565  (.L_HI(net1565));
 sg13g2_tiehi \shift_storage.storage[179]$_SDFFE_PN0P__1566  (.L_HI(net1566));
 sg13g2_tiehi \shift_storage.storage[17]$_SDFFE_PN0P__1567  (.L_HI(net1567));
 sg13g2_tiehi \shift_storage.storage[180]$_SDFFE_PN0P__1568  (.L_HI(net1568));
 sg13g2_tiehi \shift_storage.storage[181]$_SDFFE_PN0P__1569  (.L_HI(net1569));
 sg13g2_tiehi \shift_storage.storage[182]$_SDFFE_PN0P__1570  (.L_HI(net1570));
 sg13g2_tiehi \shift_storage.storage[183]$_SDFFE_PN0P__1571  (.L_HI(net1571));
 sg13g2_tiehi \shift_storage.storage[184]$_SDFFE_PN0P__1572  (.L_HI(net1572));
 sg13g2_tiehi \shift_storage.storage[185]$_SDFFE_PN0P__1573  (.L_HI(net1573));
 sg13g2_tiehi \shift_storage.storage[186]$_SDFFE_PN0P__1574  (.L_HI(net1574));
 sg13g2_tiehi \shift_storage.storage[187]$_SDFFE_PN0P__1575  (.L_HI(net1575));
 sg13g2_tiehi \shift_storage.storage[188]$_SDFFE_PN0P__1576  (.L_HI(net1576));
 sg13g2_tiehi \shift_storage.storage[189]$_SDFFE_PN0P__1577  (.L_HI(net1577));
 sg13g2_tiehi \shift_storage.storage[18]$_SDFFE_PN0P__1578  (.L_HI(net1578));
 sg13g2_tiehi \shift_storage.storage[190]$_SDFFE_PN0P__1579  (.L_HI(net1579));
 sg13g2_tiehi \shift_storage.storage[191]$_SDFFE_PN0P__1580  (.L_HI(net1580));
 sg13g2_tiehi \shift_storage.storage[192]$_SDFFE_PN0P__1581  (.L_HI(net1581));
 sg13g2_tiehi \shift_storage.storage[193]$_SDFFE_PN0P__1582  (.L_HI(net1582));
 sg13g2_tiehi \shift_storage.storage[194]$_SDFFE_PN0P__1583  (.L_HI(net1583));
 sg13g2_tiehi \shift_storage.storage[195]$_SDFFE_PN0P__1584  (.L_HI(net1584));
 sg13g2_tiehi \shift_storage.storage[196]$_SDFFE_PN0P__1585  (.L_HI(net1585));
 sg13g2_tiehi \shift_storage.storage[197]$_SDFFE_PN0P__1586  (.L_HI(net1586));
 sg13g2_tiehi \shift_storage.storage[198]$_SDFFE_PN0P__1587  (.L_HI(net1587));
 sg13g2_tiehi \shift_storage.storage[199]$_SDFFE_PN0P__1588  (.L_HI(net1588));
 sg13g2_tiehi \shift_storage.storage[19]$_SDFFE_PN0P__1589  (.L_HI(net1589));
 sg13g2_tiehi \shift_storage.storage[1]$_SDFFE_PN0P__1590  (.L_HI(net1590));
 sg13g2_tiehi \shift_storage.storage[200]$_SDFFE_PN0P__1591  (.L_HI(net1591));
 sg13g2_tiehi \shift_storage.storage[201]$_SDFFE_PN0P__1592  (.L_HI(net1592));
 sg13g2_tiehi \shift_storage.storage[202]$_SDFFE_PN0P__1593  (.L_HI(net1593));
 sg13g2_tiehi \shift_storage.storage[203]$_SDFFE_PN0P__1594  (.L_HI(net1594));
 sg13g2_tiehi \shift_storage.storage[204]$_SDFFE_PN0P__1595  (.L_HI(net1595));
 sg13g2_tiehi \shift_storage.storage[205]$_SDFFE_PN0P__1596  (.L_HI(net1596));
 sg13g2_tiehi \shift_storage.storage[206]$_SDFFE_PN0P__1597  (.L_HI(net1597));
 sg13g2_tiehi \shift_storage.storage[207]$_SDFFE_PN0P__1598  (.L_HI(net1598));
 sg13g2_tiehi \shift_storage.storage[208]$_SDFFE_PN0P__1599  (.L_HI(net1599));
 sg13g2_tiehi \shift_storage.storage[209]$_SDFFE_PN0P__1600  (.L_HI(net1600));
 sg13g2_tiehi \shift_storage.storage[20]$_SDFFE_PN0P__1601  (.L_HI(net1601));
 sg13g2_tiehi \shift_storage.storage[210]$_SDFFE_PN0P__1602  (.L_HI(net1602));
 sg13g2_tiehi \shift_storage.storage[211]$_SDFFE_PN0P__1603  (.L_HI(net1603));
 sg13g2_tiehi \shift_storage.storage[212]$_SDFFE_PN0P__1604  (.L_HI(net1604));
 sg13g2_tiehi \shift_storage.storage[213]$_SDFFE_PN0P__1605  (.L_HI(net1605));
 sg13g2_tiehi \shift_storage.storage[214]$_SDFFE_PN0P__1606  (.L_HI(net1606));
 sg13g2_tiehi \shift_storage.storage[215]$_SDFFE_PN0P__1607  (.L_HI(net1607));
 sg13g2_tiehi \shift_storage.storage[216]$_SDFFE_PN0P__1608  (.L_HI(net1608));
 sg13g2_tiehi \shift_storage.storage[217]$_SDFFE_PN0P__1609  (.L_HI(net1609));
 sg13g2_tiehi \shift_storage.storage[218]$_SDFFE_PN0P__1610  (.L_HI(net1610));
 sg13g2_tiehi \shift_storage.storage[219]$_SDFFE_PN0P__1611  (.L_HI(net1611));
 sg13g2_tiehi \shift_storage.storage[21]$_SDFFE_PN0P__1612  (.L_HI(net1612));
 sg13g2_tiehi \shift_storage.storage[220]$_SDFFE_PN0P__1613  (.L_HI(net1613));
 sg13g2_tiehi \shift_storage.storage[221]$_SDFFE_PN0P__1614  (.L_HI(net1614));
 sg13g2_tiehi \shift_storage.storage[222]$_SDFFE_PN0P__1615  (.L_HI(net1615));
 sg13g2_tiehi \shift_storage.storage[223]$_SDFFE_PN0P__1616  (.L_HI(net1616));
 sg13g2_tiehi \shift_storage.storage[224]$_SDFFE_PN0P__1617  (.L_HI(net1617));
 sg13g2_tiehi \shift_storage.storage[225]$_SDFFE_PN0P__1618  (.L_HI(net1618));
 sg13g2_tiehi \shift_storage.storage[226]$_SDFFE_PN0P__1619  (.L_HI(net1619));
 sg13g2_tiehi \shift_storage.storage[227]$_SDFFE_PN0P__1620  (.L_HI(net1620));
 sg13g2_tiehi \shift_storage.storage[228]$_SDFFE_PN0P__1621  (.L_HI(net1621));
 sg13g2_tiehi \shift_storage.storage[229]$_SDFFE_PN0P__1622  (.L_HI(net1622));
 sg13g2_tiehi \shift_storage.storage[22]$_SDFFE_PN0P__1623  (.L_HI(net1623));
 sg13g2_tiehi \shift_storage.storage[230]$_SDFFE_PN0P__1624  (.L_HI(net1624));
 sg13g2_tiehi \shift_storage.storage[231]$_SDFFE_PN0P__1625  (.L_HI(net1625));
 sg13g2_tiehi \shift_storage.storage[232]$_SDFFE_PN0P__1626  (.L_HI(net1626));
 sg13g2_tiehi \shift_storage.storage[233]$_SDFFE_PN0P__1627  (.L_HI(net1627));
 sg13g2_tiehi \shift_storage.storage[234]$_SDFFE_PN0P__1628  (.L_HI(net1628));
 sg13g2_tiehi \shift_storage.storage[235]$_SDFFE_PN0P__1629  (.L_HI(net1629));
 sg13g2_tiehi \shift_storage.storage[236]$_SDFFE_PN0P__1630  (.L_HI(net1630));
 sg13g2_tiehi \shift_storage.storage[237]$_SDFFE_PN0P__1631  (.L_HI(net1631));
 sg13g2_tiehi \shift_storage.storage[238]$_SDFFE_PN0P__1632  (.L_HI(net1632));
 sg13g2_tiehi \shift_storage.storage[239]$_SDFFE_PN0P__1633  (.L_HI(net1633));
 sg13g2_tiehi \shift_storage.storage[23]$_SDFFE_PN0P__1634  (.L_HI(net1634));
 sg13g2_tiehi \shift_storage.storage[240]$_SDFFE_PN0P__1635  (.L_HI(net1635));
 sg13g2_tiehi \shift_storage.storage[241]$_SDFFE_PN0P__1636  (.L_HI(net1636));
 sg13g2_tiehi \shift_storage.storage[242]$_SDFFE_PN0P__1637  (.L_HI(net1637));
 sg13g2_tiehi \shift_storage.storage[243]$_SDFFE_PN0P__1638  (.L_HI(net1638));
 sg13g2_tiehi \shift_storage.storage[244]$_SDFFE_PN0P__1639  (.L_HI(net1639));
 sg13g2_tiehi \shift_storage.storage[245]$_SDFFE_PN0P__1640  (.L_HI(net1640));
 sg13g2_tiehi \shift_storage.storage[246]$_SDFFE_PN0P__1641  (.L_HI(net1641));
 sg13g2_tiehi \shift_storage.storage[247]$_SDFFE_PN0P__1642  (.L_HI(net1642));
 sg13g2_tiehi \shift_storage.storage[248]$_SDFFE_PN0P__1643  (.L_HI(net1643));
 sg13g2_tiehi \shift_storage.storage[249]$_SDFFE_PN0P__1644  (.L_HI(net1644));
 sg13g2_tiehi \shift_storage.storage[24]$_SDFFE_PN0P__1645  (.L_HI(net1645));
 sg13g2_tiehi \shift_storage.storage[250]$_SDFFE_PN0P__1646  (.L_HI(net1646));
 sg13g2_tiehi \shift_storage.storage[251]$_SDFFE_PN0P__1647  (.L_HI(net1647));
 sg13g2_tiehi \shift_storage.storage[252]$_SDFFE_PN0P__1648  (.L_HI(net1648));
 sg13g2_tiehi \shift_storage.storage[253]$_SDFFE_PN0P__1649  (.L_HI(net1649));
 sg13g2_tiehi \shift_storage.storage[254]$_SDFFE_PN0P__1650  (.L_HI(net1650));
 sg13g2_tiehi \shift_storage.storage[255]$_SDFFE_PN0P__1651  (.L_HI(net1651));
 sg13g2_tiehi \shift_storage.storage[256]$_SDFFE_PN0P__1652  (.L_HI(net1652));
 sg13g2_tiehi \shift_storage.storage[257]$_SDFFE_PN0P__1653  (.L_HI(net1653));
 sg13g2_tiehi \shift_storage.storage[258]$_SDFFE_PN0P__1654  (.L_HI(net1654));
 sg13g2_tiehi \shift_storage.storage[259]$_SDFFE_PN0P__1655  (.L_HI(net1655));
 sg13g2_tiehi \shift_storage.storage[25]$_SDFFE_PN0P__1656  (.L_HI(net1656));
 sg13g2_tiehi \shift_storage.storage[260]$_SDFFE_PN0P__1657  (.L_HI(net1657));
 sg13g2_tiehi \shift_storage.storage[261]$_SDFFE_PN0P__1658  (.L_HI(net1658));
 sg13g2_tiehi \shift_storage.storage[262]$_SDFFE_PN0P__1659  (.L_HI(net1659));
 sg13g2_tiehi \shift_storage.storage[263]$_SDFFE_PN0P__1660  (.L_HI(net1660));
 sg13g2_tiehi \shift_storage.storage[264]$_SDFFE_PN0P__1661  (.L_HI(net1661));
 sg13g2_tiehi \shift_storage.storage[265]$_SDFFE_PN0P__1662  (.L_HI(net1662));
 sg13g2_tiehi \shift_storage.storage[266]$_SDFFE_PN0P__1663  (.L_HI(net1663));
 sg13g2_tiehi \shift_storage.storage[267]$_SDFFE_PN0P__1664  (.L_HI(net1664));
 sg13g2_tiehi \shift_storage.storage[268]$_SDFFE_PN0P__1665  (.L_HI(net1665));
 sg13g2_tiehi \shift_storage.storage[269]$_SDFFE_PN0P__1666  (.L_HI(net1666));
 sg13g2_tiehi \shift_storage.storage[26]$_SDFFE_PN0P__1667  (.L_HI(net1667));
 sg13g2_tiehi \shift_storage.storage[270]$_SDFFE_PN0P__1668  (.L_HI(net1668));
 sg13g2_tiehi \shift_storage.storage[271]$_SDFFE_PN0P__1669  (.L_HI(net1669));
 sg13g2_tiehi \shift_storage.storage[272]$_SDFFE_PN0P__1670  (.L_HI(net1670));
 sg13g2_tiehi \shift_storage.storage[273]$_SDFFE_PN0P__1671  (.L_HI(net1671));
 sg13g2_tiehi \shift_storage.storage[274]$_SDFFE_PN0P__1672  (.L_HI(net1672));
 sg13g2_tiehi \shift_storage.storage[275]$_SDFFE_PN0P__1673  (.L_HI(net1673));
 sg13g2_tiehi \shift_storage.storage[276]$_SDFFE_PN0P__1674  (.L_HI(net1674));
 sg13g2_tiehi \shift_storage.storage[277]$_SDFFE_PN0P__1675  (.L_HI(net1675));
 sg13g2_tiehi \shift_storage.storage[278]$_SDFFE_PN0P__1676  (.L_HI(net1676));
 sg13g2_tiehi \shift_storage.storage[279]$_SDFFE_PN0P__1677  (.L_HI(net1677));
 sg13g2_tiehi \shift_storage.storage[27]$_SDFFE_PN0P__1678  (.L_HI(net1678));
 sg13g2_tiehi \shift_storage.storage[280]$_SDFFE_PN0P__1679  (.L_HI(net1679));
 sg13g2_tiehi \shift_storage.storage[281]$_SDFFE_PN0P__1680  (.L_HI(net1680));
 sg13g2_tiehi \shift_storage.storage[282]$_SDFFE_PN0P__1681  (.L_HI(net1681));
 sg13g2_tiehi \shift_storage.storage[283]$_SDFFE_PN0P__1682  (.L_HI(net1682));
 sg13g2_tiehi \shift_storage.storage[284]$_SDFFE_PN0P__1683  (.L_HI(net1683));
 sg13g2_tiehi \shift_storage.storage[285]$_SDFFE_PN0P__1684  (.L_HI(net1684));
 sg13g2_tiehi \shift_storage.storage[286]$_SDFFE_PN0P__1685  (.L_HI(net1685));
 sg13g2_tiehi \shift_storage.storage[287]$_SDFFE_PN0P__1686  (.L_HI(net1686));
 sg13g2_tiehi \shift_storage.storage[288]$_SDFFE_PN0P__1687  (.L_HI(net1687));
 sg13g2_tiehi \shift_storage.storage[289]$_SDFFE_PN0P__1688  (.L_HI(net1688));
 sg13g2_tiehi \shift_storage.storage[28]$_SDFFE_PN0P__1689  (.L_HI(net1689));
 sg13g2_tiehi \shift_storage.storage[290]$_SDFFE_PN0P__1690  (.L_HI(net1690));
 sg13g2_tiehi \shift_storage.storage[291]$_SDFFE_PN0P__1691  (.L_HI(net1691));
 sg13g2_tiehi \shift_storage.storage[292]$_SDFFE_PN0P__1692  (.L_HI(net1692));
 sg13g2_tiehi \shift_storage.storage[293]$_SDFFE_PN0P__1693  (.L_HI(net1693));
 sg13g2_tiehi \shift_storage.storage[294]$_SDFFE_PN0P__1694  (.L_HI(net1694));
 sg13g2_tiehi \shift_storage.storage[295]$_SDFFE_PN0P__1695  (.L_HI(net1695));
 sg13g2_tiehi \shift_storage.storage[296]$_SDFFE_PN0P__1696  (.L_HI(net1696));
 sg13g2_tiehi \shift_storage.storage[297]$_SDFFE_PN0P__1697  (.L_HI(net1697));
 sg13g2_tiehi \shift_storage.storage[298]$_SDFFE_PN0P__1698  (.L_HI(net1698));
 sg13g2_tiehi \shift_storage.storage[299]$_SDFFE_PN0P__1699  (.L_HI(net1699));
 sg13g2_tiehi \shift_storage.storage[29]$_SDFFE_PN0P__1700  (.L_HI(net1700));
 sg13g2_tiehi \shift_storage.storage[2]$_SDFFE_PN0P__1701  (.L_HI(net1701));
 sg13g2_tiehi \shift_storage.storage[300]$_SDFFE_PN0P__1702  (.L_HI(net1702));
 sg13g2_tiehi \shift_storage.storage[301]$_SDFFE_PN0P__1703  (.L_HI(net1703));
 sg13g2_tiehi \shift_storage.storage[302]$_SDFFE_PN0P__1704  (.L_HI(net1704));
 sg13g2_tiehi \shift_storage.storage[303]$_SDFFE_PN0P__1705  (.L_HI(net1705));
 sg13g2_tiehi \shift_storage.storage[304]$_SDFFE_PN0P__1706  (.L_HI(net1706));
 sg13g2_tiehi \shift_storage.storage[305]$_SDFFE_PN0P__1707  (.L_HI(net1707));
 sg13g2_tiehi \shift_storage.storage[306]$_SDFFE_PN0P__1708  (.L_HI(net1708));
 sg13g2_tiehi \shift_storage.storage[307]$_SDFFE_PN0P__1709  (.L_HI(net1709));
 sg13g2_tiehi \shift_storage.storage[308]$_SDFFE_PN0P__1710  (.L_HI(net1710));
 sg13g2_tiehi \shift_storage.storage[309]$_SDFFE_PN0P__1711  (.L_HI(net1711));
 sg13g2_tiehi \shift_storage.storage[30]$_SDFFE_PN0P__1712  (.L_HI(net1712));
 sg13g2_tiehi \shift_storage.storage[310]$_SDFFE_PN0P__1713  (.L_HI(net1713));
 sg13g2_tiehi \shift_storage.storage[311]$_SDFFE_PN0P__1714  (.L_HI(net1714));
 sg13g2_tiehi \shift_storage.storage[312]$_SDFFE_PN0P__1715  (.L_HI(net1715));
 sg13g2_tiehi \shift_storage.storage[313]$_SDFFE_PN0P__1716  (.L_HI(net1716));
 sg13g2_tiehi \shift_storage.storage[314]$_SDFFE_PN0P__1717  (.L_HI(net1717));
 sg13g2_tiehi \shift_storage.storage[315]$_SDFFE_PN0P__1718  (.L_HI(net1718));
 sg13g2_tiehi \shift_storage.storage[316]$_SDFFE_PN0P__1719  (.L_HI(net1719));
 sg13g2_tiehi \shift_storage.storage[317]$_SDFFE_PN0P__1720  (.L_HI(net1720));
 sg13g2_tiehi \shift_storage.storage[318]$_SDFFE_PN0P__1721  (.L_HI(net1721));
 sg13g2_tiehi \shift_storage.storage[319]$_SDFFE_PN0P__1722  (.L_HI(net1722));
 sg13g2_tiehi \shift_storage.storage[31]$_SDFFE_PN0P__1723  (.L_HI(net1723));
 sg13g2_tiehi \shift_storage.storage[320]$_SDFFE_PN0P__1724  (.L_HI(net1724));
 sg13g2_tiehi \shift_storage.storage[321]$_SDFFE_PN0P__1725  (.L_HI(net1725));
 sg13g2_tiehi \shift_storage.storage[322]$_SDFFE_PN0P__1726  (.L_HI(net1726));
 sg13g2_tiehi \shift_storage.storage[323]$_SDFFE_PN0P__1727  (.L_HI(net1727));
 sg13g2_tiehi \shift_storage.storage[324]$_SDFFE_PN0P__1728  (.L_HI(net1728));
 sg13g2_tiehi \shift_storage.storage[325]$_SDFFE_PN0P__1729  (.L_HI(net1729));
 sg13g2_tiehi \shift_storage.storage[326]$_SDFFE_PN0P__1730  (.L_HI(net1730));
 sg13g2_tiehi \shift_storage.storage[327]$_SDFFE_PN0P__1731  (.L_HI(net1731));
 sg13g2_tiehi \shift_storage.storage[328]$_SDFFE_PN0P__1732  (.L_HI(net1732));
 sg13g2_tiehi \shift_storage.storage[329]$_SDFFE_PN0P__1733  (.L_HI(net1733));
 sg13g2_tiehi \shift_storage.storage[32]$_SDFFE_PN0P__1734  (.L_HI(net1734));
 sg13g2_tiehi \shift_storage.storage[330]$_SDFFE_PN0P__1735  (.L_HI(net1735));
 sg13g2_tiehi \shift_storage.storage[331]$_SDFFE_PN0P__1736  (.L_HI(net1736));
 sg13g2_tiehi \shift_storage.storage[332]$_SDFFE_PN0P__1737  (.L_HI(net1737));
 sg13g2_tiehi \shift_storage.storage[333]$_SDFFE_PN0P__1738  (.L_HI(net1738));
 sg13g2_tiehi \shift_storage.storage[334]$_SDFFE_PN0P__1739  (.L_HI(net1739));
 sg13g2_tiehi \shift_storage.storage[335]$_SDFFE_PN0P__1740  (.L_HI(net1740));
 sg13g2_tiehi \shift_storage.storage[336]$_SDFFE_PN0P__1741  (.L_HI(net1741));
 sg13g2_tiehi \shift_storage.storage[337]$_SDFFE_PN0P__1742  (.L_HI(net1742));
 sg13g2_tiehi \shift_storage.storage[338]$_SDFFE_PN0P__1743  (.L_HI(net1743));
 sg13g2_tiehi \shift_storage.storage[339]$_SDFFE_PN0P__1744  (.L_HI(net1744));
 sg13g2_tiehi \shift_storage.storage[33]$_SDFFE_PN0P__1745  (.L_HI(net1745));
 sg13g2_tiehi \shift_storage.storage[340]$_SDFFE_PN0P__1746  (.L_HI(net1746));
 sg13g2_tiehi \shift_storage.storage[341]$_SDFFE_PN0P__1747  (.L_HI(net1747));
 sg13g2_tiehi \shift_storage.storage[342]$_SDFFE_PN0P__1748  (.L_HI(net1748));
 sg13g2_tiehi \shift_storage.storage[343]$_SDFFE_PN0P__1749  (.L_HI(net1749));
 sg13g2_tiehi \shift_storage.storage[344]$_SDFFE_PN0P__1750  (.L_HI(net1750));
 sg13g2_tiehi \shift_storage.storage[345]$_SDFFE_PN0P__1751  (.L_HI(net1751));
 sg13g2_tiehi \shift_storage.storage[346]$_SDFFE_PN0P__1752  (.L_HI(net1752));
 sg13g2_tiehi \shift_storage.storage[347]$_SDFFE_PN0P__1753  (.L_HI(net1753));
 sg13g2_tiehi \shift_storage.storage[348]$_SDFFE_PN0P__1754  (.L_HI(net1754));
 sg13g2_tiehi \shift_storage.storage[349]$_SDFFE_PN0P__1755  (.L_HI(net1755));
 sg13g2_tiehi \shift_storage.storage[34]$_SDFFE_PN0P__1756  (.L_HI(net1756));
 sg13g2_tiehi \shift_storage.storage[350]$_SDFFE_PN0P__1757  (.L_HI(net1757));
 sg13g2_tiehi \shift_storage.storage[351]$_SDFFE_PN0P__1758  (.L_HI(net1758));
 sg13g2_tiehi \shift_storage.storage[352]$_SDFFE_PN0P__1759  (.L_HI(net1759));
 sg13g2_tiehi \shift_storage.storage[353]$_SDFFE_PN0P__1760  (.L_HI(net1760));
 sg13g2_tiehi \shift_storage.storage[354]$_SDFFE_PN0P__1761  (.L_HI(net1761));
 sg13g2_tiehi \shift_storage.storage[355]$_SDFFE_PN0P__1762  (.L_HI(net1762));
 sg13g2_tiehi \shift_storage.storage[356]$_SDFFE_PN0P__1763  (.L_HI(net1763));
 sg13g2_tiehi \shift_storage.storage[357]$_SDFFE_PN0P__1764  (.L_HI(net1764));
 sg13g2_tiehi \shift_storage.storage[358]$_SDFFE_PN0P__1765  (.L_HI(net1765));
 sg13g2_tiehi \shift_storage.storage[359]$_SDFFE_PN0P__1766  (.L_HI(net1766));
 sg13g2_tiehi \shift_storage.storage[35]$_SDFFE_PN0P__1767  (.L_HI(net1767));
 sg13g2_tiehi \shift_storage.storage[360]$_SDFFE_PN0P__1768  (.L_HI(net1768));
 sg13g2_tiehi \shift_storage.storage[361]$_SDFFE_PN0P__1769  (.L_HI(net1769));
 sg13g2_tiehi \shift_storage.storage[362]$_SDFFE_PN0P__1770  (.L_HI(net1770));
 sg13g2_tiehi \shift_storage.storage[363]$_SDFFE_PN0P__1771  (.L_HI(net1771));
 sg13g2_tiehi \shift_storage.storage[364]$_SDFFE_PN0P__1772  (.L_HI(net1772));
 sg13g2_tiehi \shift_storage.storage[365]$_SDFFE_PN0P__1773  (.L_HI(net1773));
 sg13g2_tiehi \shift_storage.storage[366]$_SDFFE_PN0P__1774  (.L_HI(net1774));
 sg13g2_tiehi \shift_storage.storage[367]$_SDFFE_PN0P__1775  (.L_HI(net1775));
 sg13g2_tiehi \shift_storage.storage[368]$_SDFFE_PN0P__1776  (.L_HI(net1776));
 sg13g2_tiehi \shift_storage.storage[369]$_SDFFE_PN0P__1777  (.L_HI(net1777));
 sg13g2_tiehi \shift_storage.storage[36]$_SDFFE_PN0P__1778  (.L_HI(net1778));
 sg13g2_tiehi \shift_storage.storage[370]$_SDFFE_PN0P__1779  (.L_HI(net1779));
 sg13g2_tiehi \shift_storage.storage[371]$_SDFFE_PN0P__1780  (.L_HI(net1780));
 sg13g2_tiehi \shift_storage.storage[372]$_SDFFE_PN0P__1781  (.L_HI(net1781));
 sg13g2_tiehi \shift_storage.storage[373]$_SDFFE_PN0P__1782  (.L_HI(net1782));
 sg13g2_tiehi \shift_storage.storage[374]$_SDFFE_PN0P__1783  (.L_HI(net1783));
 sg13g2_tiehi \shift_storage.storage[375]$_SDFFE_PN0P__1784  (.L_HI(net1784));
 sg13g2_tiehi \shift_storage.storage[376]$_SDFFE_PN0P__1785  (.L_HI(net1785));
 sg13g2_tiehi \shift_storage.storage[377]$_SDFFE_PN0P__1786  (.L_HI(net1786));
 sg13g2_tiehi \shift_storage.storage[378]$_SDFFE_PN0P__1787  (.L_HI(net1787));
 sg13g2_tiehi \shift_storage.storage[379]$_SDFFE_PN0P__1788  (.L_HI(net1788));
 sg13g2_tiehi \shift_storage.storage[37]$_SDFFE_PN0P__1789  (.L_HI(net1789));
 sg13g2_tiehi \shift_storage.storage[380]$_SDFFE_PN0P__1790  (.L_HI(net1790));
 sg13g2_tiehi \shift_storage.storage[381]$_SDFFE_PN0P__1791  (.L_HI(net1791));
 sg13g2_tiehi \shift_storage.storage[382]$_SDFFE_PN0P__1792  (.L_HI(net1792));
 sg13g2_tiehi \shift_storage.storage[383]$_SDFFE_PN0P__1793  (.L_HI(net1793));
 sg13g2_tiehi \shift_storage.storage[384]$_SDFFE_PN0P__1794  (.L_HI(net1794));
 sg13g2_tiehi \shift_storage.storage[385]$_SDFFE_PN0P__1795  (.L_HI(net1795));
 sg13g2_tiehi \shift_storage.storage[386]$_SDFFE_PN0P__1796  (.L_HI(net1796));
 sg13g2_tiehi \shift_storage.storage[387]$_SDFFE_PN0P__1797  (.L_HI(net1797));
 sg13g2_tiehi \shift_storage.storage[388]$_SDFFE_PN0P__1798  (.L_HI(net1798));
 sg13g2_tiehi \shift_storage.storage[389]$_SDFFE_PN0P__1799  (.L_HI(net1799));
 sg13g2_tiehi \shift_storage.storage[38]$_SDFFE_PN0P__1800  (.L_HI(net1800));
 sg13g2_tiehi \shift_storage.storage[390]$_SDFFE_PN0P__1801  (.L_HI(net1801));
 sg13g2_tiehi \shift_storage.storage[391]$_SDFFE_PN0P__1802  (.L_HI(net1802));
 sg13g2_tiehi \shift_storage.storage[392]$_SDFFE_PN0P__1803  (.L_HI(net1803));
 sg13g2_tiehi \shift_storage.storage[393]$_SDFFE_PN0P__1804  (.L_HI(net1804));
 sg13g2_tiehi \shift_storage.storage[394]$_SDFFE_PN0P__1805  (.L_HI(net1805));
 sg13g2_tiehi \shift_storage.storage[395]$_SDFFE_PN0P__1806  (.L_HI(net1806));
 sg13g2_tiehi \shift_storage.storage[396]$_SDFFE_PN0P__1807  (.L_HI(net1807));
 sg13g2_tiehi \shift_storage.storage[397]$_SDFFE_PN0P__1808  (.L_HI(net1808));
 sg13g2_tiehi \shift_storage.storage[398]$_SDFFE_PN0P__1809  (.L_HI(net1809));
 sg13g2_tiehi \shift_storage.storage[399]$_SDFFE_PN0P__1810  (.L_HI(net1810));
 sg13g2_tiehi \shift_storage.storage[39]$_SDFFE_PN0P__1811  (.L_HI(net1811));
 sg13g2_tiehi \shift_storage.storage[3]$_SDFFE_PN0P__1812  (.L_HI(net1812));
 sg13g2_tiehi \shift_storage.storage[400]$_SDFFE_PN0P__1813  (.L_HI(net1813));
 sg13g2_tiehi \shift_storage.storage[401]$_SDFFE_PN0P__1814  (.L_HI(net1814));
 sg13g2_tiehi \shift_storage.storage[402]$_SDFFE_PN0P__1815  (.L_HI(net1815));
 sg13g2_tiehi \shift_storage.storage[403]$_SDFFE_PN0P__1816  (.L_HI(net1816));
 sg13g2_tiehi \shift_storage.storage[404]$_SDFFE_PN0P__1817  (.L_HI(net1817));
 sg13g2_tiehi \shift_storage.storage[405]$_SDFFE_PN0P__1818  (.L_HI(net1818));
 sg13g2_tiehi \shift_storage.storage[406]$_SDFFE_PN0P__1819  (.L_HI(net1819));
 sg13g2_tiehi \shift_storage.storage[407]$_SDFFE_PN0P__1820  (.L_HI(net1820));
 sg13g2_tiehi \shift_storage.storage[408]$_SDFFE_PN0P__1821  (.L_HI(net1821));
 sg13g2_tiehi \shift_storage.storage[409]$_SDFFE_PN0P__1822  (.L_HI(net1822));
 sg13g2_tiehi \shift_storage.storage[40]$_SDFFE_PN0P__1823  (.L_HI(net1823));
 sg13g2_tiehi \shift_storage.storage[410]$_SDFFE_PN0P__1824  (.L_HI(net1824));
 sg13g2_tiehi \shift_storage.storage[411]$_SDFFE_PN0P__1825  (.L_HI(net1825));
 sg13g2_tiehi \shift_storage.storage[412]$_SDFFE_PN0P__1826  (.L_HI(net1826));
 sg13g2_tiehi \shift_storage.storage[413]$_SDFFE_PN0P__1827  (.L_HI(net1827));
 sg13g2_tiehi \shift_storage.storage[414]$_SDFFE_PN0P__1828  (.L_HI(net1828));
 sg13g2_tiehi \shift_storage.storage[415]$_SDFFE_PN0P__1829  (.L_HI(net1829));
 sg13g2_tiehi \shift_storage.storage[416]$_SDFFE_PN0P__1830  (.L_HI(net1830));
 sg13g2_tiehi \shift_storage.storage[417]$_SDFFE_PN0P__1831  (.L_HI(net1831));
 sg13g2_tiehi \shift_storage.storage[418]$_SDFFE_PN0P__1832  (.L_HI(net1832));
 sg13g2_tiehi \shift_storage.storage[419]$_SDFFE_PN0P__1833  (.L_HI(net1833));
 sg13g2_tiehi \shift_storage.storage[41]$_SDFFE_PN0P__1834  (.L_HI(net1834));
 sg13g2_tiehi \shift_storage.storage[420]$_SDFFE_PN0P__1835  (.L_HI(net1835));
 sg13g2_tiehi \shift_storage.storage[421]$_SDFFE_PN0P__1836  (.L_HI(net1836));
 sg13g2_tiehi \shift_storage.storage[422]$_SDFFE_PN0P__1837  (.L_HI(net1837));
 sg13g2_tiehi \shift_storage.storage[423]$_SDFFE_PN0P__1838  (.L_HI(net1838));
 sg13g2_tiehi \shift_storage.storage[424]$_SDFFE_PN0P__1839  (.L_HI(net1839));
 sg13g2_tiehi \shift_storage.storage[425]$_SDFFE_PN0P__1840  (.L_HI(net1840));
 sg13g2_tiehi \shift_storage.storage[426]$_SDFFE_PN0P__1841  (.L_HI(net1841));
 sg13g2_tiehi \shift_storage.storage[427]$_SDFFE_PN0P__1842  (.L_HI(net1842));
 sg13g2_tiehi \shift_storage.storage[428]$_SDFFE_PN0P__1843  (.L_HI(net1843));
 sg13g2_tiehi \shift_storage.storage[429]$_SDFFE_PN0P__1844  (.L_HI(net1844));
 sg13g2_tiehi \shift_storage.storage[42]$_SDFFE_PN0P__1845  (.L_HI(net1845));
 sg13g2_tiehi \shift_storage.storage[430]$_SDFFE_PN0P__1846  (.L_HI(net1846));
 sg13g2_tiehi \shift_storage.storage[431]$_SDFFE_PN0P__1847  (.L_HI(net1847));
 sg13g2_tiehi \shift_storage.storage[432]$_SDFFE_PN0P__1848  (.L_HI(net1848));
 sg13g2_tiehi \shift_storage.storage[433]$_SDFFE_PN0P__1849  (.L_HI(net1849));
 sg13g2_tiehi \shift_storage.storage[434]$_SDFFE_PN0P__1850  (.L_HI(net1850));
 sg13g2_tiehi \shift_storage.storage[435]$_SDFFE_PN0P__1851  (.L_HI(net1851));
 sg13g2_tiehi \shift_storage.storage[436]$_SDFFE_PN0P__1852  (.L_HI(net1852));
 sg13g2_tiehi \shift_storage.storage[437]$_SDFFE_PN0P__1853  (.L_HI(net1853));
 sg13g2_tiehi \shift_storage.storage[438]$_SDFFE_PN0P__1854  (.L_HI(net1854));
 sg13g2_tiehi \shift_storage.storage[439]$_SDFFE_PN0P__1855  (.L_HI(net1855));
 sg13g2_tiehi \shift_storage.storage[43]$_SDFFE_PN0P__1856  (.L_HI(net1856));
 sg13g2_tiehi \shift_storage.storage[440]$_SDFFE_PN0P__1857  (.L_HI(net1857));
 sg13g2_tiehi \shift_storage.storage[441]$_SDFFE_PN0P__1858  (.L_HI(net1858));
 sg13g2_tiehi \shift_storage.storage[442]$_SDFFE_PN0P__1859  (.L_HI(net1859));
 sg13g2_tiehi \shift_storage.storage[443]$_SDFFE_PN0P__1860  (.L_HI(net1860));
 sg13g2_tiehi \shift_storage.storage[444]$_SDFFE_PN0P__1861  (.L_HI(net1861));
 sg13g2_tiehi \shift_storage.storage[445]$_SDFFE_PN0P__1862  (.L_HI(net1862));
 sg13g2_tiehi \shift_storage.storage[446]$_SDFFE_PN0P__1863  (.L_HI(net1863));
 sg13g2_tiehi \shift_storage.storage[447]$_SDFFE_PN0P__1864  (.L_HI(net1864));
 sg13g2_tiehi \shift_storage.storage[448]$_SDFFE_PN0P__1865  (.L_HI(net1865));
 sg13g2_tiehi \shift_storage.storage[449]$_SDFFE_PN0P__1866  (.L_HI(net1866));
 sg13g2_tiehi \shift_storage.storage[44]$_SDFFE_PN0P__1867  (.L_HI(net1867));
 sg13g2_tiehi \shift_storage.storage[450]$_SDFFE_PN0P__1868  (.L_HI(net1868));
 sg13g2_tiehi \shift_storage.storage[451]$_SDFFE_PN0P__1869  (.L_HI(net1869));
 sg13g2_tiehi \shift_storage.storage[452]$_SDFFE_PN0P__1870  (.L_HI(net1870));
 sg13g2_tiehi \shift_storage.storage[453]$_SDFFE_PN0P__1871  (.L_HI(net1871));
 sg13g2_tiehi \shift_storage.storage[454]$_SDFFE_PN0P__1872  (.L_HI(net1872));
 sg13g2_tiehi \shift_storage.storage[455]$_SDFFE_PN0P__1873  (.L_HI(net1873));
 sg13g2_tiehi \shift_storage.storage[456]$_SDFFE_PN0P__1874  (.L_HI(net1874));
 sg13g2_tiehi \shift_storage.storage[457]$_SDFFE_PN0P__1875  (.L_HI(net1875));
 sg13g2_tiehi \shift_storage.storage[458]$_SDFFE_PN0P__1876  (.L_HI(net1876));
 sg13g2_tiehi \shift_storage.storage[459]$_SDFFE_PN0P__1877  (.L_HI(net1877));
 sg13g2_tiehi \shift_storage.storage[45]$_SDFFE_PN0P__1878  (.L_HI(net1878));
 sg13g2_tiehi \shift_storage.storage[460]$_SDFFE_PN0P__1879  (.L_HI(net1879));
 sg13g2_tiehi \shift_storage.storage[461]$_SDFFE_PN0P__1880  (.L_HI(net1880));
 sg13g2_tiehi \shift_storage.storage[462]$_SDFFE_PN0P__1881  (.L_HI(net1881));
 sg13g2_tiehi \shift_storage.storage[463]$_SDFFE_PN0P__1882  (.L_HI(net1882));
 sg13g2_tiehi \shift_storage.storage[464]$_SDFFE_PN0P__1883  (.L_HI(net1883));
 sg13g2_tiehi \shift_storage.storage[465]$_SDFFE_PN0P__1884  (.L_HI(net1884));
 sg13g2_tiehi \shift_storage.storage[466]$_SDFFE_PN0P__1885  (.L_HI(net1885));
 sg13g2_tiehi \shift_storage.storage[467]$_SDFFE_PN0P__1886  (.L_HI(net1886));
 sg13g2_tiehi \shift_storage.storage[468]$_SDFFE_PN0P__1887  (.L_HI(net1887));
 sg13g2_tiehi \shift_storage.storage[469]$_SDFFE_PN0P__1888  (.L_HI(net1888));
 sg13g2_tiehi \shift_storage.storage[46]$_SDFFE_PN0P__1889  (.L_HI(net1889));
 sg13g2_tiehi \shift_storage.storage[470]$_SDFFE_PN0P__1890  (.L_HI(net1890));
 sg13g2_tiehi \shift_storage.storage[471]$_SDFFE_PN0P__1891  (.L_HI(net1891));
 sg13g2_tiehi \shift_storage.storage[472]$_SDFFE_PN0P__1892  (.L_HI(net1892));
 sg13g2_tiehi \shift_storage.storage[473]$_SDFFE_PN0P__1893  (.L_HI(net1893));
 sg13g2_tiehi \shift_storage.storage[474]$_SDFFE_PN0P__1894  (.L_HI(net1894));
 sg13g2_tiehi \shift_storage.storage[475]$_SDFFE_PN0P__1895  (.L_HI(net1895));
 sg13g2_tiehi \shift_storage.storage[476]$_SDFFE_PN0P__1896  (.L_HI(net1896));
 sg13g2_tiehi \shift_storage.storage[477]$_SDFFE_PN0P__1897  (.L_HI(net1897));
 sg13g2_tiehi \shift_storage.storage[478]$_SDFFE_PN0P__1898  (.L_HI(net1898));
 sg13g2_tiehi \shift_storage.storage[479]$_SDFFE_PN0P__1899  (.L_HI(net1899));
 sg13g2_tiehi \shift_storage.storage[47]$_SDFFE_PN0P__1900  (.L_HI(net1900));
 sg13g2_tiehi \shift_storage.storage[480]$_SDFFE_PN0P__1901  (.L_HI(net1901));
 sg13g2_tiehi \shift_storage.storage[481]$_SDFFE_PN0P__1902  (.L_HI(net1902));
 sg13g2_tiehi \shift_storage.storage[482]$_SDFFE_PN0P__1903  (.L_HI(net1903));
 sg13g2_tiehi \shift_storage.storage[483]$_SDFFE_PN0P__1904  (.L_HI(net1904));
 sg13g2_tiehi \shift_storage.storage[484]$_SDFFE_PN0P__1905  (.L_HI(net1905));
 sg13g2_tiehi \shift_storage.storage[485]$_SDFFE_PN0P__1906  (.L_HI(net1906));
 sg13g2_tiehi \shift_storage.storage[486]$_SDFFE_PN0P__1907  (.L_HI(net1907));
 sg13g2_tiehi \shift_storage.storage[487]$_SDFFE_PN0P__1908  (.L_HI(net1908));
 sg13g2_tiehi \shift_storage.storage[488]$_SDFFE_PN0P__1909  (.L_HI(net1909));
 sg13g2_tiehi \shift_storage.storage[489]$_SDFFE_PN0P__1910  (.L_HI(net1910));
 sg13g2_tiehi \shift_storage.storage[48]$_SDFFE_PN0P__1911  (.L_HI(net1911));
 sg13g2_tiehi \shift_storage.storage[490]$_SDFFE_PN0P__1912  (.L_HI(net1912));
 sg13g2_tiehi \shift_storage.storage[491]$_SDFFE_PN0P__1913  (.L_HI(net1913));
 sg13g2_tiehi \shift_storage.storage[492]$_SDFFE_PN0P__1914  (.L_HI(net1914));
 sg13g2_tiehi \shift_storage.storage[493]$_SDFFE_PN0P__1915  (.L_HI(net1915));
 sg13g2_tiehi \shift_storage.storage[494]$_SDFFE_PN0P__1916  (.L_HI(net1916));
 sg13g2_tiehi \shift_storage.storage[495]$_SDFFE_PN0P__1917  (.L_HI(net1917));
 sg13g2_tiehi \shift_storage.storage[496]$_SDFFE_PN0P__1918  (.L_HI(net1918));
 sg13g2_tiehi \shift_storage.storage[497]$_SDFFE_PN0P__1919  (.L_HI(net1919));
 sg13g2_tiehi \shift_storage.storage[498]$_SDFFE_PN0P__1920  (.L_HI(net1920));
 sg13g2_tiehi \shift_storage.storage[499]$_SDFFE_PN0P__1921  (.L_HI(net1921));
 sg13g2_tiehi \shift_storage.storage[49]$_SDFFE_PN0P__1922  (.L_HI(net1922));
 sg13g2_tiehi \shift_storage.storage[4]$_SDFFE_PN0P__1923  (.L_HI(net1923));
 sg13g2_tiehi \shift_storage.storage[500]$_SDFFE_PN0P__1924  (.L_HI(net1924));
 sg13g2_tiehi \shift_storage.storage[501]$_SDFFE_PN0P__1925  (.L_HI(net1925));
 sg13g2_tiehi \shift_storage.storage[502]$_SDFFE_PN0P__1926  (.L_HI(net1926));
 sg13g2_tiehi \shift_storage.storage[503]$_SDFFE_PN0P__1927  (.L_HI(net1927));
 sg13g2_tiehi \shift_storage.storage[504]$_SDFFE_PN0P__1928  (.L_HI(net1928));
 sg13g2_tiehi \shift_storage.storage[505]$_SDFFE_PN0P__1929  (.L_HI(net1929));
 sg13g2_tiehi \shift_storage.storage[506]$_SDFFE_PN0P__1930  (.L_HI(net1930));
 sg13g2_tiehi \shift_storage.storage[507]$_SDFFE_PN0P__1931  (.L_HI(net1931));
 sg13g2_tiehi \shift_storage.storage[508]$_SDFFE_PN0P__1932  (.L_HI(net1932));
 sg13g2_tiehi \shift_storage.storage[509]$_SDFFE_PN0P__1933  (.L_HI(net1933));
 sg13g2_tiehi \shift_storage.storage[50]$_SDFFE_PN0P__1934  (.L_HI(net1934));
 sg13g2_tiehi \shift_storage.storage[510]$_SDFFE_PN0P__1935  (.L_HI(net1935));
 sg13g2_tiehi \shift_storage.storage[511]$_SDFFE_PN0P__1936  (.L_HI(net1936));
 sg13g2_tiehi \shift_storage.storage[512]$_SDFFE_PN0P__1937  (.L_HI(net1937));
 sg13g2_tiehi \shift_storage.storage[513]$_SDFFE_PN0P__1938  (.L_HI(net1938));
 sg13g2_tiehi \shift_storage.storage[514]$_SDFFE_PN0P__1939  (.L_HI(net1939));
 sg13g2_tiehi \shift_storage.storage[515]$_SDFFE_PN0P__1940  (.L_HI(net1940));
 sg13g2_tiehi \shift_storage.storage[516]$_SDFFE_PN0P__1941  (.L_HI(net1941));
 sg13g2_tiehi \shift_storage.storage[517]$_SDFFE_PN0P__1942  (.L_HI(net1942));
 sg13g2_tiehi \shift_storage.storage[518]$_SDFFE_PN0P__1943  (.L_HI(net1943));
 sg13g2_tiehi \shift_storage.storage[519]$_SDFFE_PN0P__1944  (.L_HI(net1944));
 sg13g2_tiehi \shift_storage.storage[51]$_SDFFE_PN0P__1945  (.L_HI(net1945));
 sg13g2_tiehi \shift_storage.storage[520]$_SDFFE_PN0P__1946  (.L_HI(net1946));
 sg13g2_tiehi \shift_storage.storage[521]$_SDFFE_PN0P__1947  (.L_HI(net1947));
 sg13g2_tiehi \shift_storage.storage[522]$_SDFFE_PN0P__1948  (.L_HI(net1948));
 sg13g2_tiehi \shift_storage.storage[523]$_SDFFE_PN0P__1949  (.L_HI(net1949));
 sg13g2_tiehi \shift_storage.storage[524]$_SDFFE_PN0P__1950  (.L_HI(net1950));
 sg13g2_tiehi \shift_storage.storage[525]$_SDFFE_PN0P__1951  (.L_HI(net1951));
 sg13g2_tiehi \shift_storage.storage[526]$_SDFFE_PN0P__1952  (.L_HI(net1952));
 sg13g2_tiehi \shift_storage.storage[527]$_SDFFE_PN0P__1953  (.L_HI(net1953));
 sg13g2_tiehi \shift_storage.storage[528]$_SDFFE_PN0P__1954  (.L_HI(net1954));
 sg13g2_tiehi \shift_storage.storage[529]$_SDFFE_PN0P__1955  (.L_HI(net1955));
 sg13g2_tiehi \shift_storage.storage[52]$_SDFFE_PN0P__1956  (.L_HI(net1956));
 sg13g2_tiehi \shift_storage.storage[530]$_SDFFE_PN0P__1957  (.L_HI(net1957));
 sg13g2_tiehi \shift_storage.storage[531]$_SDFFE_PN0P__1958  (.L_HI(net1958));
 sg13g2_tiehi \shift_storage.storage[532]$_SDFFE_PN0P__1959  (.L_HI(net1959));
 sg13g2_tiehi \shift_storage.storage[533]$_SDFFE_PN0P__1960  (.L_HI(net1960));
 sg13g2_tiehi \shift_storage.storage[534]$_SDFFE_PN0P__1961  (.L_HI(net1961));
 sg13g2_tiehi \shift_storage.storage[535]$_SDFFE_PN0P__1962  (.L_HI(net1962));
 sg13g2_tiehi \shift_storage.storage[536]$_SDFFE_PN0P__1963  (.L_HI(net1963));
 sg13g2_tiehi \shift_storage.storage[537]$_SDFFE_PN0P__1964  (.L_HI(net1964));
 sg13g2_tiehi \shift_storage.storage[538]$_SDFFE_PN0P__1965  (.L_HI(net1965));
 sg13g2_tiehi \shift_storage.storage[539]$_SDFFE_PN0P__1966  (.L_HI(net1966));
 sg13g2_tiehi \shift_storage.storage[53]$_SDFFE_PN0P__1967  (.L_HI(net1967));
 sg13g2_tiehi \shift_storage.storage[540]$_SDFFE_PN0P__1968  (.L_HI(net1968));
 sg13g2_tiehi \shift_storage.storage[541]$_SDFFE_PN0P__1969  (.L_HI(net1969));
 sg13g2_tiehi \shift_storage.storage[542]$_SDFFE_PN0P__1970  (.L_HI(net1970));
 sg13g2_tiehi \shift_storage.storage[543]$_SDFFE_PN0P__1971  (.L_HI(net1971));
 sg13g2_tiehi \shift_storage.storage[544]$_SDFFE_PN0P__1972  (.L_HI(net1972));
 sg13g2_tiehi \shift_storage.storage[545]$_SDFFE_PN0P__1973  (.L_HI(net1973));
 sg13g2_tiehi \shift_storage.storage[546]$_SDFFE_PN0P__1974  (.L_HI(net1974));
 sg13g2_tiehi \shift_storage.storage[547]$_SDFFE_PN0P__1975  (.L_HI(net1975));
 sg13g2_tiehi \shift_storage.storage[548]$_SDFFE_PN0P__1976  (.L_HI(net1976));
 sg13g2_tiehi \shift_storage.storage[549]$_SDFFE_PN0P__1977  (.L_HI(net1977));
 sg13g2_tiehi \shift_storage.storage[54]$_SDFFE_PN0P__1978  (.L_HI(net1978));
 sg13g2_tiehi \shift_storage.storage[550]$_SDFFE_PN0P__1979  (.L_HI(net1979));
 sg13g2_tiehi \shift_storage.storage[551]$_SDFFE_PN0P__1980  (.L_HI(net1980));
 sg13g2_tiehi \shift_storage.storage[552]$_SDFFE_PN0P__1981  (.L_HI(net1981));
 sg13g2_tiehi \shift_storage.storage[553]$_SDFFE_PN0P__1982  (.L_HI(net1982));
 sg13g2_tiehi \shift_storage.storage[554]$_SDFFE_PN0P__1983  (.L_HI(net1983));
 sg13g2_tiehi \shift_storage.storage[555]$_SDFFE_PN0P__1984  (.L_HI(net1984));
 sg13g2_tiehi \shift_storage.storage[556]$_SDFFE_PN0P__1985  (.L_HI(net1985));
 sg13g2_tiehi \shift_storage.storage[557]$_SDFFE_PN0P__1986  (.L_HI(net1986));
 sg13g2_tiehi \shift_storage.storage[558]$_SDFFE_PN0P__1987  (.L_HI(net1987));
 sg13g2_tiehi \shift_storage.storage[559]$_SDFFE_PN0P__1988  (.L_HI(net1988));
 sg13g2_tiehi \shift_storage.storage[55]$_SDFFE_PN0P__1989  (.L_HI(net1989));
 sg13g2_tiehi \shift_storage.storage[560]$_SDFFE_PN0P__1990  (.L_HI(net1990));
 sg13g2_tiehi \shift_storage.storage[561]$_SDFFE_PN0P__1991  (.L_HI(net1991));
 sg13g2_tiehi \shift_storage.storage[562]$_SDFFE_PN0P__1992  (.L_HI(net1992));
 sg13g2_tiehi \shift_storage.storage[563]$_SDFFE_PN0P__1993  (.L_HI(net1993));
 sg13g2_tiehi \shift_storage.storage[564]$_SDFFE_PN0P__1994  (.L_HI(net1994));
 sg13g2_tiehi \shift_storage.storage[565]$_SDFFE_PN0P__1995  (.L_HI(net1995));
 sg13g2_tiehi \shift_storage.storage[566]$_SDFFE_PN0P__1996  (.L_HI(net1996));
 sg13g2_tiehi \shift_storage.storage[567]$_SDFFE_PN0P__1997  (.L_HI(net1997));
 sg13g2_tiehi \shift_storage.storage[568]$_SDFFE_PN0P__1998  (.L_HI(net1998));
 sg13g2_tiehi \shift_storage.storage[569]$_SDFFE_PN0P__1999  (.L_HI(net1999));
 sg13g2_tiehi \shift_storage.storage[56]$_SDFFE_PN0P__2000  (.L_HI(net2000));
 sg13g2_tiehi \shift_storage.storage[570]$_SDFFE_PN0P__2001  (.L_HI(net2001));
 sg13g2_tiehi \shift_storage.storage[571]$_SDFFE_PN0P__2002  (.L_HI(net2002));
 sg13g2_tiehi \shift_storage.storage[572]$_SDFFE_PN0P__2003  (.L_HI(net2003));
 sg13g2_tiehi \shift_storage.storage[573]$_SDFFE_PN0P__2004  (.L_HI(net2004));
 sg13g2_tiehi \shift_storage.storage[574]$_SDFFE_PN0P__2005  (.L_HI(net2005));
 sg13g2_tiehi \shift_storage.storage[575]$_SDFFE_PN0P__2006  (.L_HI(net2006));
 sg13g2_tiehi \shift_storage.storage[576]$_SDFFE_PN0P__2007  (.L_HI(net2007));
 sg13g2_tiehi \shift_storage.storage[577]$_SDFFE_PN0P__2008  (.L_HI(net2008));
 sg13g2_tiehi \shift_storage.storage[578]$_SDFFE_PN0P__2009  (.L_HI(net2009));
 sg13g2_tiehi \shift_storage.storage[579]$_SDFFE_PN0P__2010  (.L_HI(net2010));
 sg13g2_tiehi \shift_storage.storage[57]$_SDFFE_PN0P__2011  (.L_HI(net2011));
 sg13g2_tiehi \shift_storage.storage[580]$_SDFFE_PN0P__2012  (.L_HI(net2012));
 sg13g2_tiehi \shift_storage.storage[581]$_SDFFE_PN0P__2013  (.L_HI(net2013));
 sg13g2_tiehi \shift_storage.storage[582]$_SDFFE_PN0P__2014  (.L_HI(net2014));
 sg13g2_tiehi \shift_storage.storage[583]$_SDFFE_PN0P__2015  (.L_HI(net2015));
 sg13g2_tiehi \shift_storage.storage[584]$_SDFFE_PN0P__2016  (.L_HI(net2016));
 sg13g2_tiehi \shift_storage.storage[585]$_SDFFE_PN0P__2017  (.L_HI(net2017));
 sg13g2_tiehi \shift_storage.storage[586]$_SDFFE_PN0P__2018  (.L_HI(net2018));
 sg13g2_tiehi \shift_storage.storage[587]$_SDFFE_PN0P__2019  (.L_HI(net2019));
 sg13g2_tiehi \shift_storage.storage[588]$_SDFFE_PN0P__2020  (.L_HI(net2020));
 sg13g2_tiehi \shift_storage.storage[589]$_SDFFE_PN0P__2021  (.L_HI(net2021));
 sg13g2_tiehi \shift_storage.storage[58]$_SDFFE_PN0P__2022  (.L_HI(net2022));
 sg13g2_tiehi \shift_storage.storage[590]$_SDFFE_PN0P__2023  (.L_HI(net2023));
 sg13g2_tiehi \shift_storage.storage[591]$_SDFFE_PN0P__2024  (.L_HI(net2024));
 sg13g2_tiehi \shift_storage.storage[592]$_SDFFE_PN0P__2025  (.L_HI(net2025));
 sg13g2_tiehi \shift_storage.storage[593]$_SDFFE_PN0P__2026  (.L_HI(net2026));
 sg13g2_tiehi \shift_storage.storage[594]$_SDFFE_PN0P__2027  (.L_HI(net2027));
 sg13g2_tiehi \shift_storage.storage[595]$_SDFFE_PN0P__2028  (.L_HI(net2028));
 sg13g2_tiehi \shift_storage.storage[596]$_SDFFE_PN0P__2029  (.L_HI(net2029));
 sg13g2_tiehi \shift_storage.storage[597]$_SDFFE_PN0P__2030  (.L_HI(net2030));
 sg13g2_tiehi \shift_storage.storage[598]$_SDFFE_PN0P__2031  (.L_HI(net2031));
 sg13g2_tiehi \shift_storage.storage[599]$_SDFFE_PN0P__2032  (.L_HI(net2032));
 sg13g2_tiehi \shift_storage.storage[59]$_SDFFE_PN0P__2033  (.L_HI(net2033));
 sg13g2_tiehi \shift_storage.storage[5]$_SDFFE_PN0P__2034  (.L_HI(net2034));
 sg13g2_tiehi \shift_storage.storage[600]$_SDFFE_PN0P__2035  (.L_HI(net2035));
 sg13g2_tiehi \shift_storage.storage[601]$_SDFFE_PN0P__2036  (.L_HI(net2036));
 sg13g2_tiehi \shift_storage.storage[602]$_SDFFE_PN0P__2037  (.L_HI(net2037));
 sg13g2_tiehi \shift_storage.storage[603]$_SDFFE_PN0P__2038  (.L_HI(net2038));
 sg13g2_tiehi \shift_storage.storage[604]$_SDFFE_PN0P__2039  (.L_HI(net2039));
 sg13g2_tiehi \shift_storage.storage[605]$_SDFFE_PN0P__2040  (.L_HI(net2040));
 sg13g2_tiehi \shift_storage.storage[606]$_SDFFE_PN0P__2041  (.L_HI(net2041));
 sg13g2_tiehi \shift_storage.storage[607]$_SDFFE_PN0P__2042  (.L_HI(net2042));
 sg13g2_tiehi \shift_storage.storage[608]$_SDFFE_PN0P__2043  (.L_HI(net2043));
 sg13g2_tiehi \shift_storage.storage[609]$_SDFFE_PN0P__2044  (.L_HI(net2044));
 sg13g2_tiehi \shift_storage.storage[60]$_SDFFE_PN0P__2045  (.L_HI(net2045));
 sg13g2_tiehi \shift_storage.storage[610]$_SDFFE_PN0P__2046  (.L_HI(net2046));
 sg13g2_tiehi \shift_storage.storage[611]$_SDFFE_PN0P__2047  (.L_HI(net2047));
 sg13g2_tiehi \shift_storage.storage[612]$_SDFFE_PN0P__2048  (.L_HI(net2048));
 sg13g2_tiehi \shift_storage.storage[613]$_SDFFE_PN0P__2049  (.L_HI(net2049));
 sg13g2_tiehi \shift_storage.storage[614]$_SDFFE_PN0P__2050  (.L_HI(net2050));
 sg13g2_tiehi \shift_storage.storage[615]$_SDFFE_PN0P__2051  (.L_HI(net2051));
 sg13g2_tiehi \shift_storage.storage[616]$_SDFFE_PN0P__2052  (.L_HI(net2052));
 sg13g2_tiehi \shift_storage.storage[617]$_SDFFE_PN0P__2053  (.L_HI(net2053));
 sg13g2_tiehi \shift_storage.storage[618]$_SDFFE_PN0P__2054  (.L_HI(net2054));
 sg13g2_tiehi \shift_storage.storage[619]$_SDFFE_PN0P__2055  (.L_HI(net2055));
 sg13g2_tiehi \shift_storage.storage[61]$_SDFFE_PN0P__2056  (.L_HI(net2056));
 sg13g2_tiehi \shift_storage.storage[620]$_SDFFE_PN0P__2057  (.L_HI(net2057));
 sg13g2_tiehi \shift_storage.storage[621]$_SDFFE_PN0P__2058  (.L_HI(net2058));
 sg13g2_tiehi \shift_storage.storage[622]$_SDFFE_PN0P__2059  (.L_HI(net2059));
 sg13g2_tiehi \shift_storage.storage[623]$_SDFFE_PN0P__2060  (.L_HI(net2060));
 sg13g2_tiehi \shift_storage.storage[624]$_SDFFE_PN0P__2061  (.L_HI(net2061));
 sg13g2_tiehi \shift_storage.storage[625]$_SDFFE_PN0P__2062  (.L_HI(net2062));
 sg13g2_tiehi \shift_storage.storage[626]$_SDFFE_PN0P__2063  (.L_HI(net2063));
 sg13g2_tiehi \shift_storage.storage[627]$_SDFFE_PN0P__2064  (.L_HI(net2064));
 sg13g2_tiehi \shift_storage.storage[628]$_SDFFE_PN0P__2065  (.L_HI(net2065));
 sg13g2_tiehi \shift_storage.storage[629]$_SDFFE_PN0P__2066  (.L_HI(net2066));
 sg13g2_tiehi \shift_storage.storage[62]$_SDFFE_PN0P__2067  (.L_HI(net2067));
 sg13g2_tiehi \shift_storage.storage[630]$_SDFFE_PN0P__2068  (.L_HI(net2068));
 sg13g2_tiehi \shift_storage.storage[631]$_SDFFE_PN0P__2069  (.L_HI(net2069));
 sg13g2_tiehi \shift_storage.storage[632]$_SDFFE_PN0P__2070  (.L_HI(net2070));
 sg13g2_tiehi \shift_storage.storage[633]$_SDFFE_PN0P__2071  (.L_HI(net2071));
 sg13g2_tiehi \shift_storage.storage[634]$_SDFFE_PN0P__2072  (.L_HI(net2072));
 sg13g2_tiehi \shift_storage.storage[635]$_SDFFE_PN0P__2073  (.L_HI(net2073));
 sg13g2_tiehi \shift_storage.storage[636]$_SDFFE_PN0P__2074  (.L_HI(net2074));
 sg13g2_tiehi \shift_storage.storage[637]$_SDFFE_PN0P__2075  (.L_HI(net2075));
 sg13g2_tiehi \shift_storage.storage[638]$_SDFFE_PN0P__2076  (.L_HI(net2076));
 sg13g2_tiehi \shift_storage.storage[639]$_SDFFE_PN0P__2077  (.L_HI(net2077));
 sg13g2_tiehi \shift_storage.storage[63]$_SDFFE_PN0P__2078  (.L_HI(net2078));
 sg13g2_tiehi \shift_storage.storage[640]$_SDFFE_PN0P__2079  (.L_HI(net2079));
 sg13g2_tiehi \shift_storage.storage[641]$_SDFFE_PN0P__2080  (.L_HI(net2080));
 sg13g2_tiehi \shift_storage.storage[642]$_SDFFE_PN0P__2081  (.L_HI(net2081));
 sg13g2_tiehi \shift_storage.storage[643]$_SDFFE_PN0P__2082  (.L_HI(net2082));
 sg13g2_tiehi \shift_storage.storage[644]$_SDFFE_PN0P__2083  (.L_HI(net2083));
 sg13g2_tiehi \shift_storage.storage[645]$_SDFFE_PN0P__2084  (.L_HI(net2084));
 sg13g2_tiehi \shift_storage.storage[646]$_SDFFE_PN0P__2085  (.L_HI(net2085));
 sg13g2_tiehi \shift_storage.storage[647]$_SDFFE_PN0P__2086  (.L_HI(net2086));
 sg13g2_tiehi \shift_storage.storage[648]$_SDFFE_PN0P__2087  (.L_HI(net2087));
 sg13g2_tiehi \shift_storage.storage[649]$_SDFFE_PN0P__2088  (.L_HI(net2088));
 sg13g2_tiehi \shift_storage.storage[64]$_SDFFE_PN0P__2089  (.L_HI(net2089));
 sg13g2_tiehi \shift_storage.storage[650]$_SDFFE_PN0P__2090  (.L_HI(net2090));
 sg13g2_tiehi \shift_storage.storage[651]$_SDFFE_PN0P__2091  (.L_HI(net2091));
 sg13g2_tiehi \shift_storage.storage[652]$_SDFFE_PN0P__2092  (.L_HI(net2092));
 sg13g2_tiehi \shift_storage.storage[653]$_SDFFE_PN0P__2093  (.L_HI(net2093));
 sg13g2_tiehi \shift_storage.storage[654]$_SDFFE_PN0P__2094  (.L_HI(net2094));
 sg13g2_tiehi \shift_storage.storage[655]$_SDFFE_PN0P__2095  (.L_HI(net2095));
 sg13g2_tiehi \shift_storage.storage[656]$_SDFFE_PN0P__2096  (.L_HI(net2096));
 sg13g2_tiehi \shift_storage.storage[657]$_SDFFE_PN0P__2097  (.L_HI(net2097));
 sg13g2_tiehi \shift_storage.storage[658]$_SDFFE_PN0P__2098  (.L_HI(net2098));
 sg13g2_tiehi \shift_storage.storage[659]$_SDFFE_PN0P__2099  (.L_HI(net2099));
 sg13g2_tiehi \shift_storage.storage[65]$_SDFFE_PN0P__2100  (.L_HI(net2100));
 sg13g2_tiehi \shift_storage.storage[660]$_SDFFE_PN0P__2101  (.L_HI(net2101));
 sg13g2_tiehi \shift_storage.storage[661]$_SDFFE_PN0P__2102  (.L_HI(net2102));
 sg13g2_tiehi \shift_storage.storage[662]$_SDFFE_PN0P__2103  (.L_HI(net2103));
 sg13g2_tiehi \shift_storage.storage[663]$_SDFFE_PN0P__2104  (.L_HI(net2104));
 sg13g2_tiehi \shift_storage.storage[664]$_SDFFE_PN0P__2105  (.L_HI(net2105));
 sg13g2_tiehi \shift_storage.storage[665]$_SDFFE_PN0P__2106  (.L_HI(net2106));
 sg13g2_tiehi \shift_storage.storage[666]$_SDFFE_PN0P__2107  (.L_HI(net2107));
 sg13g2_tiehi \shift_storage.storage[667]$_SDFFE_PN0P__2108  (.L_HI(net2108));
 sg13g2_tiehi \shift_storage.storage[668]$_SDFFE_PN0P__2109  (.L_HI(net2109));
 sg13g2_tiehi \shift_storage.storage[669]$_SDFFE_PN0P__2110  (.L_HI(net2110));
 sg13g2_tiehi \shift_storage.storage[66]$_SDFFE_PN0P__2111  (.L_HI(net2111));
 sg13g2_tiehi \shift_storage.storage[670]$_SDFFE_PN0P__2112  (.L_HI(net2112));
 sg13g2_tiehi \shift_storage.storage[671]$_SDFFE_PN0P__2113  (.L_HI(net2113));
 sg13g2_tiehi \shift_storage.storage[672]$_SDFFE_PN0P__2114  (.L_HI(net2114));
 sg13g2_tiehi \shift_storage.storage[673]$_SDFFE_PN0P__2115  (.L_HI(net2115));
 sg13g2_tiehi \shift_storage.storage[674]$_SDFFE_PN0P__2116  (.L_HI(net2116));
 sg13g2_tiehi \shift_storage.storage[675]$_SDFFE_PN0P__2117  (.L_HI(net2117));
 sg13g2_tiehi \shift_storage.storage[676]$_SDFFE_PN0P__2118  (.L_HI(net2118));
 sg13g2_tiehi \shift_storage.storage[677]$_SDFFE_PN0P__2119  (.L_HI(net2119));
 sg13g2_tiehi \shift_storage.storage[678]$_SDFFE_PN0P__2120  (.L_HI(net2120));
 sg13g2_tiehi \shift_storage.storage[679]$_SDFFE_PN0P__2121  (.L_HI(net2121));
 sg13g2_tiehi \shift_storage.storage[67]$_SDFFE_PN0P__2122  (.L_HI(net2122));
 sg13g2_tiehi \shift_storage.storage[680]$_SDFFE_PN0P__2123  (.L_HI(net2123));
 sg13g2_tiehi \shift_storage.storage[681]$_SDFFE_PN0P__2124  (.L_HI(net2124));
 sg13g2_tiehi \shift_storage.storage[682]$_SDFFE_PN0P__2125  (.L_HI(net2125));
 sg13g2_tiehi \shift_storage.storage[683]$_SDFFE_PN0P__2126  (.L_HI(net2126));
 sg13g2_tiehi \shift_storage.storage[684]$_SDFFE_PN0P__2127  (.L_HI(net2127));
 sg13g2_tiehi \shift_storage.storage[685]$_SDFFE_PN0P__2128  (.L_HI(net2128));
 sg13g2_tiehi \shift_storage.storage[686]$_SDFFE_PN0P__2129  (.L_HI(net2129));
 sg13g2_tiehi \shift_storage.storage[687]$_SDFFE_PN0P__2130  (.L_HI(net2130));
 sg13g2_tiehi \shift_storage.storage[688]$_SDFFE_PN0P__2131  (.L_HI(net2131));
 sg13g2_tiehi \shift_storage.storage[689]$_SDFFE_PN0P__2132  (.L_HI(net2132));
 sg13g2_tiehi \shift_storage.storage[68]$_SDFFE_PN0P__2133  (.L_HI(net2133));
 sg13g2_tiehi \shift_storage.storage[690]$_SDFFE_PN0P__2134  (.L_HI(net2134));
 sg13g2_tiehi \shift_storage.storage[691]$_SDFFE_PN0P__2135  (.L_HI(net2135));
 sg13g2_tiehi \shift_storage.storage[692]$_SDFFE_PN0P__2136  (.L_HI(net2136));
 sg13g2_tiehi \shift_storage.storage[693]$_SDFFE_PN0P__2137  (.L_HI(net2137));
 sg13g2_tiehi \shift_storage.storage[694]$_SDFFE_PN0P__2138  (.L_HI(net2138));
 sg13g2_tiehi \shift_storage.storage[695]$_SDFFE_PN0P__2139  (.L_HI(net2139));
 sg13g2_tiehi \shift_storage.storage[696]$_SDFFE_PN0P__2140  (.L_HI(net2140));
 sg13g2_tiehi \shift_storage.storage[697]$_SDFFE_PN0P__2141  (.L_HI(net2141));
 sg13g2_tiehi \shift_storage.storage[698]$_SDFFE_PN0P__2142  (.L_HI(net2142));
 sg13g2_tiehi \shift_storage.storage[699]$_SDFFE_PN0P__2143  (.L_HI(net2143));
 sg13g2_tiehi \shift_storage.storage[69]$_SDFFE_PN0P__2144  (.L_HI(net2144));
 sg13g2_tiehi \shift_storage.storage[6]$_SDFFE_PN0P__2145  (.L_HI(net2145));
 sg13g2_tiehi \shift_storage.storage[700]$_SDFFE_PN0P__2146  (.L_HI(net2146));
 sg13g2_tiehi \shift_storage.storage[701]$_SDFFE_PN0P__2147  (.L_HI(net2147));
 sg13g2_tiehi \shift_storage.storage[702]$_SDFFE_PN0P__2148  (.L_HI(net2148));
 sg13g2_tiehi \shift_storage.storage[703]$_SDFFE_PN0P__2149  (.L_HI(net2149));
 sg13g2_tiehi \shift_storage.storage[704]$_SDFFE_PN0P__2150  (.L_HI(net2150));
 sg13g2_tiehi \shift_storage.storage[705]$_SDFFE_PN0P__2151  (.L_HI(net2151));
 sg13g2_tiehi \shift_storage.storage[706]$_SDFFE_PN0P__2152  (.L_HI(net2152));
 sg13g2_tiehi \shift_storage.storage[707]$_SDFFE_PN0P__2153  (.L_HI(net2153));
 sg13g2_tiehi \shift_storage.storage[708]$_SDFFE_PN0P__2154  (.L_HI(net2154));
 sg13g2_tiehi \shift_storage.storage[709]$_SDFFE_PN0P__2155  (.L_HI(net2155));
 sg13g2_tiehi \shift_storage.storage[70]$_SDFFE_PN0P__2156  (.L_HI(net2156));
 sg13g2_tiehi \shift_storage.storage[710]$_SDFFE_PN0P__2157  (.L_HI(net2157));
 sg13g2_tiehi \shift_storage.storage[711]$_SDFFE_PN0P__2158  (.L_HI(net2158));
 sg13g2_tiehi \shift_storage.storage[712]$_SDFFE_PN0P__2159  (.L_HI(net2159));
 sg13g2_tiehi \shift_storage.storage[713]$_SDFFE_PN0P__2160  (.L_HI(net2160));
 sg13g2_tiehi \shift_storage.storage[714]$_SDFFE_PN0P__2161  (.L_HI(net2161));
 sg13g2_tiehi \shift_storage.storage[715]$_SDFFE_PN0P__2162  (.L_HI(net2162));
 sg13g2_tiehi \shift_storage.storage[716]$_SDFFE_PN0P__2163  (.L_HI(net2163));
 sg13g2_tiehi \shift_storage.storage[717]$_SDFFE_PN0P__2164  (.L_HI(net2164));
 sg13g2_tiehi \shift_storage.storage[718]$_SDFFE_PN0P__2165  (.L_HI(net2165));
 sg13g2_tiehi \shift_storage.storage[719]$_SDFFE_PN0P__2166  (.L_HI(net2166));
 sg13g2_tiehi \shift_storage.storage[71]$_SDFFE_PN0P__2167  (.L_HI(net2167));
 sg13g2_tiehi \shift_storage.storage[720]$_SDFFE_PN0P__2168  (.L_HI(net2168));
 sg13g2_tiehi \shift_storage.storage[721]$_SDFFE_PN0P__2169  (.L_HI(net2169));
 sg13g2_tiehi \shift_storage.storage[722]$_SDFFE_PN0P__2170  (.L_HI(net2170));
 sg13g2_tiehi \shift_storage.storage[723]$_SDFFE_PN0P__2171  (.L_HI(net2171));
 sg13g2_tiehi \shift_storage.storage[724]$_SDFFE_PN0P__2172  (.L_HI(net2172));
 sg13g2_tiehi \shift_storage.storage[725]$_SDFFE_PN0P__2173  (.L_HI(net2173));
 sg13g2_tiehi \shift_storage.storage[726]$_SDFFE_PN0P__2174  (.L_HI(net2174));
 sg13g2_tiehi \shift_storage.storage[727]$_SDFFE_PN0P__2175  (.L_HI(net2175));
 sg13g2_tiehi \shift_storage.storage[728]$_SDFFE_PN0P__2176  (.L_HI(net2176));
 sg13g2_tiehi \shift_storage.storage[729]$_SDFFE_PN0P__2177  (.L_HI(net2177));
 sg13g2_tiehi \shift_storage.storage[72]$_SDFFE_PN0P__2178  (.L_HI(net2178));
 sg13g2_tiehi \shift_storage.storage[730]$_SDFFE_PN0P__2179  (.L_HI(net2179));
 sg13g2_tiehi \shift_storage.storage[731]$_SDFFE_PN0P__2180  (.L_HI(net2180));
 sg13g2_tiehi \shift_storage.storage[732]$_SDFFE_PN0P__2181  (.L_HI(net2181));
 sg13g2_tiehi \shift_storage.storage[733]$_SDFFE_PN0P__2182  (.L_HI(net2182));
 sg13g2_tiehi \shift_storage.storage[734]$_SDFFE_PN0P__2183  (.L_HI(net2183));
 sg13g2_tiehi \shift_storage.storage[735]$_SDFFE_PN0P__2184  (.L_HI(net2184));
 sg13g2_tiehi \shift_storage.storage[736]$_SDFFE_PN0P__2185  (.L_HI(net2185));
 sg13g2_tiehi \shift_storage.storage[737]$_SDFFE_PN0P__2186  (.L_HI(net2186));
 sg13g2_tiehi \shift_storage.storage[738]$_SDFFE_PN0P__2187  (.L_HI(net2187));
 sg13g2_tiehi \shift_storage.storage[739]$_SDFFE_PN0P__2188  (.L_HI(net2188));
 sg13g2_tiehi \shift_storage.storage[73]$_SDFFE_PN0P__2189  (.L_HI(net2189));
 sg13g2_tiehi \shift_storage.storage[740]$_SDFFE_PN0P__2190  (.L_HI(net2190));
 sg13g2_tiehi \shift_storage.storage[741]$_SDFFE_PN0P__2191  (.L_HI(net2191));
 sg13g2_tiehi \shift_storage.storage[742]$_SDFFE_PN0P__2192  (.L_HI(net2192));
 sg13g2_tiehi \shift_storage.storage[743]$_SDFFE_PN0P__2193  (.L_HI(net2193));
 sg13g2_tiehi \shift_storage.storage[744]$_SDFFE_PN0P__2194  (.L_HI(net2194));
 sg13g2_tiehi \shift_storage.storage[745]$_SDFFE_PN0P__2195  (.L_HI(net2195));
 sg13g2_tiehi \shift_storage.storage[746]$_SDFFE_PN0P__2196  (.L_HI(net2196));
 sg13g2_tiehi \shift_storage.storage[747]$_SDFFE_PN0P__2197  (.L_HI(net2197));
 sg13g2_tiehi \shift_storage.storage[748]$_SDFFE_PN0P__2198  (.L_HI(net2198));
 sg13g2_tiehi \shift_storage.storage[749]$_SDFFE_PN0P__2199  (.L_HI(net2199));
 sg13g2_tiehi \shift_storage.storage[74]$_SDFFE_PN0P__2200  (.L_HI(net2200));
 sg13g2_tiehi \shift_storage.storage[750]$_SDFFE_PN0P__2201  (.L_HI(net2201));
 sg13g2_tiehi \shift_storage.storage[751]$_SDFFE_PN0P__2202  (.L_HI(net2202));
 sg13g2_tiehi \shift_storage.storage[752]$_SDFFE_PN0P__2203  (.L_HI(net2203));
 sg13g2_tiehi \shift_storage.storage[753]$_SDFFE_PN0P__2204  (.L_HI(net2204));
 sg13g2_tiehi \shift_storage.storage[754]$_SDFFE_PN0P__2205  (.L_HI(net2205));
 sg13g2_tiehi \shift_storage.storage[755]$_SDFFE_PN0P__2206  (.L_HI(net2206));
 sg13g2_tiehi \shift_storage.storage[756]$_SDFFE_PN0P__2207  (.L_HI(net2207));
 sg13g2_tiehi \shift_storage.storage[757]$_SDFFE_PN0P__2208  (.L_HI(net2208));
 sg13g2_tiehi \shift_storage.storage[758]$_SDFFE_PN0P__2209  (.L_HI(net2209));
 sg13g2_tiehi \shift_storage.storage[759]$_SDFFE_PN0P__2210  (.L_HI(net2210));
 sg13g2_tiehi \shift_storage.storage[75]$_SDFFE_PN0P__2211  (.L_HI(net2211));
 sg13g2_tiehi \shift_storage.storage[760]$_SDFFE_PN0P__2212  (.L_HI(net2212));
 sg13g2_tiehi \shift_storage.storage[761]$_SDFFE_PN0P__2213  (.L_HI(net2213));
 sg13g2_tiehi \shift_storage.storage[762]$_SDFFE_PN0P__2214  (.L_HI(net2214));
 sg13g2_tiehi \shift_storage.storage[763]$_SDFFE_PN0P__2215  (.L_HI(net2215));
 sg13g2_tiehi \shift_storage.storage[764]$_SDFFE_PN0P__2216  (.L_HI(net2216));
 sg13g2_tiehi \shift_storage.storage[765]$_SDFFE_PN0P__2217  (.L_HI(net2217));
 sg13g2_tiehi \shift_storage.storage[766]$_SDFFE_PN0P__2218  (.L_HI(net2218));
 sg13g2_tiehi \shift_storage.storage[767]$_SDFFE_PN0P__2219  (.L_HI(net2219));
 sg13g2_tiehi \shift_storage.storage[768]$_SDFFE_PN0P__2220  (.L_HI(net2220));
 sg13g2_tiehi \shift_storage.storage[769]$_SDFFE_PN0P__2221  (.L_HI(net2221));
 sg13g2_tiehi \shift_storage.storage[76]$_SDFFE_PN0P__2222  (.L_HI(net2222));
 sg13g2_tiehi \shift_storage.storage[770]$_SDFFE_PN0P__2223  (.L_HI(net2223));
 sg13g2_tiehi \shift_storage.storage[771]$_SDFFE_PN0P__2224  (.L_HI(net2224));
 sg13g2_tiehi \shift_storage.storage[772]$_SDFFE_PN0P__2225  (.L_HI(net2225));
 sg13g2_tiehi \shift_storage.storage[773]$_SDFFE_PN0P__2226  (.L_HI(net2226));
 sg13g2_tiehi \shift_storage.storage[774]$_SDFFE_PN0P__2227  (.L_HI(net2227));
 sg13g2_tiehi \shift_storage.storage[775]$_SDFFE_PN0P__2228  (.L_HI(net2228));
 sg13g2_tiehi \shift_storage.storage[776]$_SDFFE_PN0P__2229  (.L_HI(net2229));
 sg13g2_tiehi \shift_storage.storage[777]$_SDFFE_PN0P__2230  (.L_HI(net2230));
 sg13g2_tiehi \shift_storage.storage[778]$_SDFFE_PN0P__2231  (.L_HI(net2231));
 sg13g2_tiehi \shift_storage.storage[779]$_SDFFE_PN0P__2232  (.L_HI(net2232));
 sg13g2_tiehi \shift_storage.storage[77]$_SDFFE_PN0P__2233  (.L_HI(net2233));
 sg13g2_tiehi \shift_storage.storage[780]$_SDFFE_PN0P__2234  (.L_HI(net2234));
 sg13g2_tiehi \shift_storage.storage[781]$_SDFFE_PN0P__2235  (.L_HI(net2235));
 sg13g2_tiehi \shift_storage.storage[782]$_SDFFE_PN0P__2236  (.L_HI(net2236));
 sg13g2_tiehi \shift_storage.storage[783]$_SDFFE_PN0P__2237  (.L_HI(net2237));
 sg13g2_tiehi \shift_storage.storage[784]$_SDFFE_PN0P__2238  (.L_HI(net2238));
 sg13g2_tiehi \shift_storage.storage[785]$_SDFFE_PN0P__2239  (.L_HI(net2239));
 sg13g2_tiehi \shift_storage.storage[786]$_SDFFE_PN0P__2240  (.L_HI(net2240));
 sg13g2_tiehi \shift_storage.storage[787]$_SDFFE_PN0P__2241  (.L_HI(net2241));
 sg13g2_tiehi \shift_storage.storage[788]$_SDFFE_PN0P__2242  (.L_HI(net2242));
 sg13g2_tiehi \shift_storage.storage[789]$_SDFFE_PN0P__2243  (.L_HI(net2243));
 sg13g2_tiehi \shift_storage.storage[78]$_SDFFE_PN0P__2244  (.L_HI(net2244));
 sg13g2_tiehi \shift_storage.storage[790]$_SDFFE_PN0P__2245  (.L_HI(net2245));
 sg13g2_tiehi \shift_storage.storage[791]$_SDFFE_PN0P__2246  (.L_HI(net2246));
 sg13g2_tiehi \shift_storage.storage[792]$_SDFFE_PN0P__2247  (.L_HI(net2247));
 sg13g2_tiehi \shift_storage.storage[793]$_SDFFE_PN0P__2248  (.L_HI(net2248));
 sg13g2_tiehi \shift_storage.storage[794]$_SDFFE_PN0P__2249  (.L_HI(net2249));
 sg13g2_tiehi \shift_storage.storage[795]$_SDFFE_PN0P__2250  (.L_HI(net2250));
 sg13g2_tiehi \shift_storage.storage[796]$_SDFFE_PN0P__2251  (.L_HI(net2251));
 sg13g2_tiehi \shift_storage.storage[797]$_SDFFE_PN0P__2252  (.L_HI(net2252));
 sg13g2_tiehi \shift_storage.storage[798]$_SDFFE_PN0P__2253  (.L_HI(net2253));
 sg13g2_tiehi \shift_storage.storage[799]$_SDFFE_PN0P__2254  (.L_HI(net2254));
 sg13g2_tiehi \shift_storage.storage[79]$_SDFFE_PN0P__2255  (.L_HI(net2255));
 sg13g2_tiehi \shift_storage.storage[7]$_SDFFE_PN0P__2256  (.L_HI(net2256));
 sg13g2_tiehi \shift_storage.storage[800]$_SDFFE_PN0P__2257  (.L_HI(net2257));
 sg13g2_tiehi \shift_storage.storage[801]$_SDFFE_PN0P__2258  (.L_HI(net2258));
 sg13g2_tiehi \shift_storage.storage[802]$_SDFFE_PN0P__2259  (.L_HI(net2259));
 sg13g2_tiehi \shift_storage.storage[803]$_SDFFE_PN0P__2260  (.L_HI(net2260));
 sg13g2_tiehi \shift_storage.storage[804]$_SDFFE_PN0P__2261  (.L_HI(net2261));
 sg13g2_tiehi \shift_storage.storage[805]$_SDFFE_PN0P__2262  (.L_HI(net2262));
 sg13g2_tiehi \shift_storage.storage[806]$_SDFFE_PN0P__2263  (.L_HI(net2263));
 sg13g2_tiehi \shift_storage.storage[807]$_SDFFE_PN0P__2264  (.L_HI(net2264));
 sg13g2_tiehi \shift_storage.storage[808]$_SDFFE_PN0P__2265  (.L_HI(net2265));
 sg13g2_tiehi \shift_storage.storage[809]$_SDFFE_PN0P__2266  (.L_HI(net2266));
 sg13g2_tiehi \shift_storage.storage[80]$_SDFFE_PN0P__2267  (.L_HI(net2267));
 sg13g2_tiehi \shift_storage.storage[810]$_SDFFE_PN0P__2268  (.L_HI(net2268));
 sg13g2_tiehi \shift_storage.storage[811]$_SDFFE_PN0P__2269  (.L_HI(net2269));
 sg13g2_tiehi \shift_storage.storage[812]$_SDFFE_PN0P__2270  (.L_HI(net2270));
 sg13g2_tiehi \shift_storage.storage[813]$_SDFFE_PN0P__2271  (.L_HI(net2271));
 sg13g2_tiehi \shift_storage.storage[814]$_SDFFE_PN0P__2272  (.L_HI(net2272));
 sg13g2_tiehi \shift_storage.storage[815]$_SDFFE_PN0P__2273  (.L_HI(net2273));
 sg13g2_tiehi \shift_storage.storage[816]$_SDFFE_PN0P__2274  (.L_HI(net2274));
 sg13g2_tiehi \shift_storage.storage[817]$_SDFFE_PN0P__2275  (.L_HI(net2275));
 sg13g2_tiehi \shift_storage.storage[818]$_SDFFE_PN0P__2276  (.L_HI(net2276));
 sg13g2_tiehi \shift_storage.storage[819]$_SDFFE_PN0P__2277  (.L_HI(net2277));
 sg13g2_tiehi \shift_storage.storage[81]$_SDFFE_PN0P__2278  (.L_HI(net2278));
 sg13g2_tiehi \shift_storage.storage[820]$_SDFFE_PN0P__2279  (.L_HI(net2279));
 sg13g2_tiehi \shift_storage.storage[821]$_SDFFE_PN0P__2280  (.L_HI(net2280));
 sg13g2_tiehi \shift_storage.storage[822]$_SDFFE_PN0P__2281  (.L_HI(net2281));
 sg13g2_tiehi \shift_storage.storage[823]$_SDFFE_PN0P__2282  (.L_HI(net2282));
 sg13g2_tiehi \shift_storage.storage[824]$_SDFFE_PN0P__2283  (.L_HI(net2283));
 sg13g2_tiehi \shift_storage.storage[825]$_SDFFE_PN0P__2284  (.L_HI(net2284));
 sg13g2_tiehi \shift_storage.storage[826]$_SDFFE_PN0P__2285  (.L_HI(net2285));
 sg13g2_tiehi \shift_storage.storage[827]$_SDFFE_PN0P__2286  (.L_HI(net2286));
 sg13g2_tiehi \shift_storage.storage[828]$_SDFFE_PN0P__2287  (.L_HI(net2287));
 sg13g2_tiehi \shift_storage.storage[829]$_SDFFE_PN0P__2288  (.L_HI(net2288));
 sg13g2_tiehi \shift_storage.storage[82]$_SDFFE_PN0P__2289  (.L_HI(net2289));
 sg13g2_tiehi \shift_storage.storage[830]$_SDFFE_PN0P__2290  (.L_HI(net2290));
 sg13g2_tiehi \shift_storage.storage[831]$_SDFFE_PN0P__2291  (.L_HI(net2291));
 sg13g2_tiehi \shift_storage.storage[832]$_SDFFE_PN0P__2292  (.L_HI(net2292));
 sg13g2_tiehi \shift_storage.storage[833]$_SDFFE_PN0P__2293  (.L_HI(net2293));
 sg13g2_tiehi \shift_storage.storage[834]$_SDFFE_PN0P__2294  (.L_HI(net2294));
 sg13g2_tiehi \shift_storage.storage[835]$_SDFFE_PN0P__2295  (.L_HI(net2295));
 sg13g2_tiehi \shift_storage.storage[836]$_SDFFE_PN0P__2296  (.L_HI(net2296));
 sg13g2_tiehi \shift_storage.storage[837]$_SDFFE_PN0P__2297  (.L_HI(net2297));
 sg13g2_tiehi \shift_storage.storage[838]$_SDFFE_PN0P__2298  (.L_HI(net2298));
 sg13g2_tiehi \shift_storage.storage[839]$_SDFFE_PN0P__2299  (.L_HI(net2299));
 sg13g2_tiehi \shift_storage.storage[83]$_SDFFE_PN0P__2300  (.L_HI(net2300));
 sg13g2_tiehi \shift_storage.storage[840]$_SDFFE_PN0P__2301  (.L_HI(net2301));
 sg13g2_tiehi \shift_storage.storage[841]$_SDFFE_PN0P__2302  (.L_HI(net2302));
 sg13g2_tiehi \shift_storage.storage[842]$_SDFFE_PN0P__2303  (.L_HI(net2303));
 sg13g2_tiehi \shift_storage.storage[843]$_SDFFE_PN0P__2304  (.L_HI(net2304));
 sg13g2_tiehi \shift_storage.storage[844]$_SDFFE_PN0P__2305  (.L_HI(net2305));
 sg13g2_tiehi \shift_storage.storage[845]$_SDFFE_PN0P__2306  (.L_HI(net2306));
 sg13g2_tiehi \shift_storage.storage[846]$_SDFFE_PN0P__2307  (.L_HI(net2307));
 sg13g2_tiehi \shift_storage.storage[847]$_SDFFE_PN0P__2308  (.L_HI(net2308));
 sg13g2_tiehi \shift_storage.storage[848]$_SDFFE_PN0P__2309  (.L_HI(net2309));
 sg13g2_tiehi \shift_storage.storage[849]$_SDFFE_PN0P__2310  (.L_HI(net2310));
 sg13g2_tiehi \shift_storage.storage[84]$_SDFFE_PN0P__2311  (.L_HI(net2311));
 sg13g2_tiehi \shift_storage.storage[850]$_SDFFE_PN0P__2312  (.L_HI(net2312));
 sg13g2_tiehi \shift_storage.storage[851]$_SDFFE_PN0P__2313  (.L_HI(net2313));
 sg13g2_tiehi \shift_storage.storage[852]$_SDFFE_PN0P__2314  (.L_HI(net2314));
 sg13g2_tiehi \shift_storage.storage[853]$_SDFFE_PN0P__2315  (.L_HI(net2315));
 sg13g2_tiehi \shift_storage.storage[854]$_SDFFE_PN0P__2316  (.L_HI(net2316));
 sg13g2_tiehi \shift_storage.storage[855]$_SDFFE_PN0P__2317  (.L_HI(net2317));
 sg13g2_tiehi \shift_storage.storage[856]$_SDFFE_PN0P__2318  (.L_HI(net2318));
 sg13g2_tiehi \shift_storage.storage[857]$_SDFFE_PN0P__2319  (.L_HI(net2319));
 sg13g2_tiehi \shift_storage.storage[858]$_SDFFE_PN0P__2320  (.L_HI(net2320));
 sg13g2_tiehi \shift_storage.storage[859]$_SDFFE_PN0P__2321  (.L_HI(net2321));
 sg13g2_tiehi \shift_storage.storage[85]$_SDFFE_PN0P__2322  (.L_HI(net2322));
 sg13g2_tiehi \shift_storage.storage[860]$_SDFFE_PN0P__2323  (.L_HI(net2323));
 sg13g2_tiehi \shift_storage.storage[861]$_SDFFE_PN0P__2324  (.L_HI(net2324));
 sg13g2_tiehi \shift_storage.storage[862]$_SDFFE_PN0P__2325  (.L_HI(net2325));
 sg13g2_tiehi \shift_storage.storage[863]$_SDFFE_PN0P__2326  (.L_HI(net2326));
 sg13g2_tiehi \shift_storage.storage[864]$_SDFFE_PN0P__2327  (.L_HI(net2327));
 sg13g2_tiehi \shift_storage.storage[865]$_SDFFE_PN0P__2328  (.L_HI(net2328));
 sg13g2_tiehi \shift_storage.storage[866]$_SDFFE_PN0P__2329  (.L_HI(net2329));
 sg13g2_tiehi \shift_storage.storage[867]$_SDFFE_PN0P__2330  (.L_HI(net2330));
 sg13g2_tiehi \shift_storage.storage[868]$_SDFFE_PN0P__2331  (.L_HI(net2331));
 sg13g2_tiehi \shift_storage.storage[869]$_SDFFE_PN0P__2332  (.L_HI(net2332));
 sg13g2_tiehi \shift_storage.storage[86]$_SDFFE_PN0P__2333  (.L_HI(net2333));
 sg13g2_tiehi \shift_storage.storage[870]$_SDFFE_PN0P__2334  (.L_HI(net2334));
 sg13g2_tiehi \shift_storage.storage[871]$_SDFFE_PN0P__2335  (.L_HI(net2335));
 sg13g2_tiehi \shift_storage.storage[872]$_SDFFE_PN0P__2336  (.L_HI(net2336));
 sg13g2_tiehi \shift_storage.storage[873]$_SDFFE_PN0P__2337  (.L_HI(net2337));
 sg13g2_tiehi \shift_storage.storage[874]$_SDFFE_PN0P__2338  (.L_HI(net2338));
 sg13g2_tiehi \shift_storage.storage[875]$_SDFFE_PN0P__2339  (.L_HI(net2339));
 sg13g2_tiehi \shift_storage.storage[876]$_SDFFE_PN0P__2340  (.L_HI(net2340));
 sg13g2_tiehi \shift_storage.storage[877]$_SDFFE_PN0P__2341  (.L_HI(net2341));
 sg13g2_tiehi \shift_storage.storage[878]$_SDFFE_PN0P__2342  (.L_HI(net2342));
 sg13g2_tiehi \shift_storage.storage[879]$_SDFFE_PN0P__2343  (.L_HI(net2343));
 sg13g2_tiehi \shift_storage.storage[87]$_SDFFE_PN0P__2344  (.L_HI(net2344));
 sg13g2_tiehi \shift_storage.storage[880]$_SDFFE_PN0P__2345  (.L_HI(net2345));
 sg13g2_tiehi \shift_storage.storage[881]$_SDFFE_PN0P__2346  (.L_HI(net2346));
 sg13g2_tiehi \shift_storage.storage[882]$_SDFFE_PN0P__2347  (.L_HI(net2347));
 sg13g2_tiehi \shift_storage.storage[883]$_SDFFE_PN0P__2348  (.L_HI(net2348));
 sg13g2_tiehi \shift_storage.storage[884]$_SDFFE_PN0P__2349  (.L_HI(net2349));
 sg13g2_tiehi \shift_storage.storage[885]$_SDFFE_PN0P__2350  (.L_HI(net2350));
 sg13g2_tiehi \shift_storage.storage[886]$_SDFFE_PN0P__2351  (.L_HI(net2351));
 sg13g2_tiehi \shift_storage.storage[887]$_SDFFE_PN0P__2352  (.L_HI(net2352));
 sg13g2_tiehi \shift_storage.storage[888]$_SDFFE_PN0P__2353  (.L_HI(net2353));
 sg13g2_tiehi \shift_storage.storage[889]$_SDFFE_PN0P__2354  (.L_HI(net2354));
 sg13g2_tiehi \shift_storage.storage[88]$_SDFFE_PN0P__2355  (.L_HI(net2355));
 sg13g2_tiehi \shift_storage.storage[890]$_SDFFE_PN0P__2356  (.L_HI(net2356));
 sg13g2_tiehi \shift_storage.storage[891]$_SDFFE_PN0P__2357  (.L_HI(net2357));
 sg13g2_tiehi \shift_storage.storage[892]$_SDFFE_PN0P__2358  (.L_HI(net2358));
 sg13g2_tiehi \shift_storage.storage[893]$_SDFFE_PN0P__2359  (.L_HI(net2359));
 sg13g2_tiehi \shift_storage.storage[894]$_SDFFE_PN0P__2360  (.L_HI(net2360));
 sg13g2_tiehi \shift_storage.storage[895]$_SDFFE_PN0P__2361  (.L_HI(net2361));
 sg13g2_tiehi \shift_storage.storage[896]$_SDFFE_PN0P__2362  (.L_HI(net2362));
 sg13g2_tiehi \shift_storage.storage[897]$_SDFFE_PN0P__2363  (.L_HI(net2363));
 sg13g2_tiehi \shift_storage.storage[898]$_SDFFE_PN0P__2364  (.L_HI(net2364));
 sg13g2_tiehi \shift_storage.storage[899]$_SDFFE_PN0P__2365  (.L_HI(net2365));
 sg13g2_tiehi \shift_storage.storage[89]$_SDFFE_PN0P__2366  (.L_HI(net2366));
 sg13g2_tiehi \shift_storage.storage[8]$_SDFFE_PN0P__2367  (.L_HI(net2367));
 sg13g2_tiehi \shift_storage.storage[900]$_SDFFE_PN0P__2368  (.L_HI(net2368));
 sg13g2_tiehi \shift_storage.storage[901]$_SDFFE_PN0P__2369  (.L_HI(net2369));
 sg13g2_tiehi \shift_storage.storage[902]$_SDFFE_PN0P__2370  (.L_HI(net2370));
 sg13g2_tiehi \shift_storage.storage[903]$_SDFFE_PN0P__2371  (.L_HI(net2371));
 sg13g2_tiehi \shift_storage.storage[904]$_SDFFE_PN0P__2372  (.L_HI(net2372));
 sg13g2_tiehi \shift_storage.storage[905]$_SDFFE_PN0P__2373  (.L_HI(net2373));
 sg13g2_tiehi \shift_storage.storage[906]$_SDFFE_PN0P__2374  (.L_HI(net2374));
 sg13g2_tiehi \shift_storage.storage[907]$_SDFFE_PN0P__2375  (.L_HI(net2375));
 sg13g2_tiehi \shift_storage.storage[908]$_SDFFE_PN0P__2376  (.L_HI(net2376));
 sg13g2_tiehi \shift_storage.storage[909]$_SDFFE_PN0P__2377  (.L_HI(net2377));
 sg13g2_tiehi \shift_storage.storage[90]$_SDFFE_PN0P__2378  (.L_HI(net2378));
 sg13g2_tiehi \shift_storage.storage[910]$_SDFFE_PN0P__2379  (.L_HI(net2379));
 sg13g2_tiehi \shift_storage.storage[911]$_SDFFE_PN0P__2380  (.L_HI(net2380));
 sg13g2_tiehi \shift_storage.storage[912]$_SDFFE_PN0P__2381  (.L_HI(net2381));
 sg13g2_tiehi \shift_storage.storage[913]$_SDFFE_PN0P__2382  (.L_HI(net2382));
 sg13g2_tiehi \shift_storage.storage[914]$_SDFFE_PN0P__2383  (.L_HI(net2383));
 sg13g2_tiehi \shift_storage.storage[915]$_SDFFE_PN0P__2384  (.L_HI(net2384));
 sg13g2_tiehi \shift_storage.storage[916]$_SDFFE_PN0P__2385  (.L_HI(net2385));
 sg13g2_tiehi \shift_storage.storage[917]$_SDFFE_PN0P__2386  (.L_HI(net2386));
 sg13g2_tiehi \shift_storage.storage[918]$_SDFFE_PN0P__2387  (.L_HI(net2387));
 sg13g2_tiehi \shift_storage.storage[919]$_SDFFE_PN0P__2388  (.L_HI(net2388));
 sg13g2_tiehi \shift_storage.storage[91]$_SDFFE_PN0P__2389  (.L_HI(net2389));
 sg13g2_tiehi \shift_storage.storage[920]$_SDFFE_PN0P__2390  (.L_HI(net2390));
 sg13g2_tiehi \shift_storage.storage[921]$_SDFFE_PN0P__2391  (.L_HI(net2391));
 sg13g2_tiehi \shift_storage.storage[922]$_SDFFE_PN0P__2392  (.L_HI(net2392));
 sg13g2_tiehi \shift_storage.storage[923]$_SDFFE_PN0P__2393  (.L_HI(net2393));
 sg13g2_tiehi \shift_storage.storage[924]$_SDFFE_PN0P__2394  (.L_HI(net2394));
 sg13g2_tiehi \shift_storage.storage[925]$_SDFFE_PN0P__2395  (.L_HI(net2395));
 sg13g2_tiehi \shift_storage.storage[926]$_SDFFE_PN0P__2396  (.L_HI(net2396));
 sg13g2_tiehi \shift_storage.storage[927]$_SDFFE_PN0P__2397  (.L_HI(net2397));
 sg13g2_tiehi \shift_storage.storage[928]$_SDFFE_PN0P__2398  (.L_HI(net2398));
 sg13g2_tiehi \shift_storage.storage[929]$_SDFFE_PN0P__2399  (.L_HI(net2399));
 sg13g2_tiehi \shift_storage.storage[92]$_SDFFE_PN0P__2400  (.L_HI(net2400));
 sg13g2_tiehi \shift_storage.storage[930]$_SDFFE_PN0P__2401  (.L_HI(net2401));
 sg13g2_tiehi \shift_storage.storage[931]$_SDFFE_PN0P__2402  (.L_HI(net2402));
 sg13g2_tiehi \shift_storage.storage[932]$_SDFFE_PN0P__2403  (.L_HI(net2403));
 sg13g2_tiehi \shift_storage.storage[933]$_SDFFE_PN0P__2404  (.L_HI(net2404));
 sg13g2_tiehi \shift_storage.storage[934]$_SDFFE_PN0P__2405  (.L_HI(net2405));
 sg13g2_tiehi \shift_storage.storage[935]$_SDFFE_PN0P__2406  (.L_HI(net2406));
 sg13g2_tiehi \shift_storage.storage[936]$_SDFFE_PN0P__2407  (.L_HI(net2407));
 sg13g2_tiehi \shift_storage.storage[937]$_SDFFE_PN0P__2408  (.L_HI(net2408));
 sg13g2_tiehi \shift_storage.storage[938]$_SDFFE_PN0P__2409  (.L_HI(net2409));
 sg13g2_tiehi \shift_storage.storage[939]$_SDFFE_PN0P__2410  (.L_HI(net2410));
 sg13g2_tiehi \shift_storage.storage[93]$_SDFFE_PN0P__2411  (.L_HI(net2411));
 sg13g2_tiehi \shift_storage.storage[940]$_SDFFE_PN0P__2412  (.L_HI(net2412));
 sg13g2_tiehi \shift_storage.storage[941]$_SDFFE_PN0P__2413  (.L_HI(net2413));
 sg13g2_tiehi \shift_storage.storage[942]$_SDFFE_PN0P__2414  (.L_HI(net2414));
 sg13g2_tiehi \shift_storage.storage[943]$_SDFFE_PN0P__2415  (.L_HI(net2415));
 sg13g2_tiehi \shift_storage.storage[944]$_SDFFE_PN0P__2416  (.L_HI(net2416));
 sg13g2_tiehi \shift_storage.storage[945]$_SDFFE_PN0P__2417  (.L_HI(net2417));
 sg13g2_tiehi \shift_storage.storage[946]$_SDFFE_PN0P__2418  (.L_HI(net2418));
 sg13g2_tiehi \shift_storage.storage[947]$_SDFFE_PN0P__2419  (.L_HI(net2419));
 sg13g2_tiehi \shift_storage.storage[948]$_SDFFE_PN0P__2420  (.L_HI(net2420));
 sg13g2_tiehi \shift_storage.storage[949]$_SDFFE_PN0P__2421  (.L_HI(net2421));
 sg13g2_tiehi \shift_storage.storage[94]$_SDFFE_PN0P__2422  (.L_HI(net2422));
 sg13g2_tiehi \shift_storage.storage[950]$_SDFFE_PN0P__2423  (.L_HI(net2423));
 sg13g2_tiehi \shift_storage.storage[951]$_SDFFE_PN0P__2424  (.L_HI(net2424));
 sg13g2_tiehi \shift_storage.storage[952]$_SDFFE_PN0P__2425  (.L_HI(net2425));
 sg13g2_tiehi \shift_storage.storage[953]$_SDFFE_PN0P__2426  (.L_HI(net2426));
 sg13g2_tiehi \shift_storage.storage[954]$_SDFFE_PN0P__2427  (.L_HI(net2427));
 sg13g2_tiehi \shift_storage.storage[955]$_SDFFE_PN0P__2428  (.L_HI(net2428));
 sg13g2_tiehi \shift_storage.storage[956]$_SDFFE_PN0P__2429  (.L_HI(net2429));
 sg13g2_tiehi \shift_storage.storage[957]$_SDFFE_PN0P__2430  (.L_HI(net2430));
 sg13g2_tiehi \shift_storage.storage[958]$_SDFFE_PN0P__2431  (.L_HI(net2431));
 sg13g2_tiehi \shift_storage.storage[959]$_SDFFE_PN0P__2432  (.L_HI(net2432));
 sg13g2_tiehi \shift_storage.storage[95]$_SDFFE_PN0P__2433  (.L_HI(net2433));
 sg13g2_tiehi \shift_storage.storage[960]$_SDFFE_PN0P__2434  (.L_HI(net2434));
 sg13g2_tiehi \shift_storage.storage[961]$_SDFFE_PN0P__2435  (.L_HI(net2435));
 sg13g2_tiehi \shift_storage.storage[962]$_SDFFE_PN0P__2436  (.L_HI(net2436));
 sg13g2_tiehi \shift_storage.storage[963]$_SDFFE_PN0P__2437  (.L_HI(net2437));
 sg13g2_tiehi \shift_storage.storage[964]$_SDFFE_PN0P__2438  (.L_HI(net2438));
 sg13g2_tiehi \shift_storage.storage[965]$_SDFFE_PN0P__2439  (.L_HI(net2439));
 sg13g2_tiehi \shift_storage.storage[966]$_SDFFE_PN0P__2440  (.L_HI(net2440));
 sg13g2_tiehi \shift_storage.storage[967]$_SDFFE_PN0P__2441  (.L_HI(net2441));
 sg13g2_tiehi \shift_storage.storage[968]$_SDFFE_PN0P__2442  (.L_HI(net2442));
 sg13g2_tiehi \shift_storage.storage[969]$_SDFFE_PN0P__2443  (.L_HI(net2443));
 sg13g2_tiehi \shift_storage.storage[96]$_SDFFE_PN0P__2444  (.L_HI(net2444));
 sg13g2_tiehi \shift_storage.storage[970]$_SDFFE_PN0P__2445  (.L_HI(net2445));
 sg13g2_tiehi \shift_storage.storage[971]$_SDFFE_PN0P__2446  (.L_HI(net2446));
 sg13g2_tiehi \shift_storage.storage[972]$_SDFFE_PN0P__2447  (.L_HI(net2447));
 sg13g2_tiehi \shift_storage.storage[973]$_SDFFE_PN0P__2448  (.L_HI(net2448));
 sg13g2_tiehi \shift_storage.storage[974]$_SDFFE_PN0P__2449  (.L_HI(net2449));
 sg13g2_tiehi \shift_storage.storage[975]$_SDFFE_PN0P__2450  (.L_HI(net2450));
 sg13g2_tiehi \shift_storage.storage[976]$_SDFFE_PN0P__2451  (.L_HI(net2451));
 sg13g2_tiehi \shift_storage.storage[977]$_SDFFE_PN0P__2452  (.L_HI(net2452));
 sg13g2_tiehi \shift_storage.storage[978]$_SDFFE_PN0P__2453  (.L_HI(net2453));
 sg13g2_tiehi \shift_storage.storage[979]$_SDFFE_PN0P__2454  (.L_HI(net2454));
 sg13g2_tiehi \shift_storage.storage[97]$_SDFFE_PN0P__2455  (.L_HI(net2455));
 sg13g2_tiehi \shift_storage.storage[980]$_SDFFE_PN0P__2456  (.L_HI(net2456));
 sg13g2_tiehi \shift_storage.storage[981]$_SDFFE_PN0P__2457  (.L_HI(net2457));
 sg13g2_tiehi \shift_storage.storage[982]$_SDFFE_PN0P__2458  (.L_HI(net2458));
 sg13g2_tiehi \shift_storage.storage[983]$_SDFFE_PN0P__2459  (.L_HI(net2459));
 sg13g2_tiehi \shift_storage.storage[984]$_SDFFE_PN0P__2460  (.L_HI(net2460));
 sg13g2_tiehi \shift_storage.storage[985]$_SDFFE_PN0P__2461  (.L_HI(net2461));
 sg13g2_tiehi \shift_storage.storage[986]$_SDFFE_PN0P__2462  (.L_HI(net2462));
 sg13g2_tiehi \shift_storage.storage[987]$_SDFFE_PN0P__2463  (.L_HI(net2463));
 sg13g2_tiehi \shift_storage.storage[988]$_SDFFE_PN0P__2464  (.L_HI(net2464));
 sg13g2_tiehi \shift_storage.storage[989]$_SDFFE_PN0P__2465  (.L_HI(net2465));
 sg13g2_tiehi \shift_storage.storage[98]$_SDFFE_PN0P__2466  (.L_HI(net2466));
 sg13g2_tiehi \shift_storage.storage[990]$_SDFFE_PN0P__2467  (.L_HI(net2467));
 sg13g2_tiehi \shift_storage.storage[991]$_SDFFE_PN0P__2468  (.L_HI(net2468));
 sg13g2_tiehi \shift_storage.storage[992]$_SDFFE_PN0P__2469  (.L_HI(net2469));
 sg13g2_tiehi \shift_storage.storage[993]$_SDFFE_PN0P__2470  (.L_HI(net2470));
 sg13g2_tiehi \shift_storage.storage[994]$_SDFFE_PN0P__2471  (.L_HI(net2471));
 sg13g2_tiehi \shift_storage.storage[995]$_SDFFE_PN0P__2472  (.L_HI(net2472));
 sg13g2_tiehi \shift_storage.storage[996]$_SDFFE_PN0P__2473  (.L_HI(net2473));
 sg13g2_tiehi \shift_storage.storage[997]$_SDFFE_PN0P__2474  (.L_HI(net2474));
 sg13g2_tiehi \shift_storage.storage[998]$_SDFFE_PN0P__2475  (.L_HI(net2475));
 sg13g2_tiehi \shift_storage.storage[999]$_SDFFE_PN0P__2476  (.L_HI(net2476));
 sg13g2_tiehi \shift_storage.storage[99]$_SDFFE_PN0P__2477  (.L_HI(net2477));
 sg13g2_tiehi \shift_storage.storage[9]$_SDFFE_PN0P__2478  (.L_HI(net2478));
 sg13g2_buf_4 clkbuf_leaf_1_clk_p2c (.X(clknet_leaf_1_clk_p2c),
    .A(clknet_5_0__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_2_clk_p2c (.X(clknet_leaf_2_clk_p2c),
    .A(clknet_5_0__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_3_clk_p2c (.X(clknet_leaf_3_clk_p2c),
    .A(clknet_5_1__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_4_clk_p2c (.X(clknet_leaf_4_clk_p2c),
    .A(clknet_5_1__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_5_clk_p2c (.X(clknet_leaf_5_clk_p2c),
    .A(clknet_5_3__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_6_clk_p2c (.X(clknet_leaf_6_clk_p2c),
    .A(clknet_5_2__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_7_clk_p2c (.X(clknet_leaf_7_clk_p2c),
    .A(clknet_5_2__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_8_clk_p2c (.X(clknet_leaf_8_clk_p2c),
    .A(clknet_5_2__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_9_clk_p2c (.X(clknet_leaf_9_clk_p2c),
    .A(clknet_5_2__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_10_clk_p2c (.X(clknet_leaf_10_clk_p2c),
    .A(clknet_5_2__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_11_clk_p2c (.X(clknet_leaf_11_clk_p2c),
    .A(clknet_5_2__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_12_clk_p2c (.X(clknet_leaf_12_clk_p2c),
    .A(clknet_5_2__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_13_clk_p2c (.X(clknet_leaf_13_clk_p2c),
    .A(clknet_5_2__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_14_clk_p2c (.X(clknet_leaf_14_clk_p2c),
    .A(clknet_5_8__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_15_clk_p2c (.X(clknet_leaf_15_clk_p2c),
    .A(clknet_5_8__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_16_clk_p2c (.X(clknet_leaf_16_clk_p2c),
    .A(clknet_5_8__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_17_clk_p2c (.X(clknet_leaf_17_clk_p2c),
    .A(clknet_5_2__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_18_clk_p2c (.X(clknet_leaf_18_clk_p2c),
    .A(clknet_5_3__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_19_clk_p2c (.X(clknet_leaf_19_clk_p2c),
    .A(clknet_5_9__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_20_clk_p2c (.X(clknet_leaf_20_clk_p2c),
    .A(clknet_5_9__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_21_clk_p2c (.X(clknet_leaf_21_clk_p2c),
    .A(clknet_5_3__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_22_clk_p2c (.X(clknet_leaf_22_clk_p2c),
    .A(clknet_5_3__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_23_clk_p2c (.X(clknet_leaf_23_clk_p2c),
    .A(clknet_5_3__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_24_clk_p2c (.X(clknet_leaf_24_clk_p2c),
    .A(clknet_5_3__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_25_clk_p2c (.X(clknet_leaf_25_clk_p2c),
    .A(clknet_5_3__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_26_clk_p2c (.X(clknet_leaf_26_clk_p2c),
    .A(clknet_5_6__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_27_clk_p2c (.X(clknet_leaf_27_clk_p2c),
    .A(clknet_5_6__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_28_clk_p2c (.X(clknet_leaf_28_clk_p2c),
    .A(clknet_5_6__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_29_clk_p2c (.X(clknet_leaf_29_clk_p2c),
    .A(clknet_5_6__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_30_clk_p2c (.X(clknet_leaf_30_clk_p2c),
    .A(clknet_5_3__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_31_clk_p2c (.X(clknet_leaf_31_clk_p2c),
    .A(clknet_5_12__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_32_clk_p2c (.X(clknet_leaf_32_clk_p2c),
    .A(clknet_5_6__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_33_clk_p2c (.X(clknet_leaf_33_clk_p2c),
    .A(clknet_5_7__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_34_clk_p2c (.X(clknet_leaf_34_clk_p2c),
    .A(clknet_5_13__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_35_clk_p2c (.X(clknet_leaf_35_clk_p2c),
    .A(clknet_5_13__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_36_clk_p2c (.X(clknet_leaf_36_clk_p2c),
    .A(clknet_5_13__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_37_clk_p2c (.X(clknet_leaf_37_clk_p2c),
    .A(clknet_5_13__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_38_clk_p2c (.X(clknet_leaf_38_clk_p2c),
    .A(clknet_5_13__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_39_clk_p2c (.X(clknet_leaf_39_clk_p2c),
    .A(clknet_5_12__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_40_clk_p2c (.X(clknet_leaf_40_clk_p2c),
    .A(clknet_5_12__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_41_clk_p2c (.X(clknet_leaf_41_clk_p2c),
    .A(clknet_5_12__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_42_clk_p2c (.X(clknet_leaf_42_clk_p2c),
    .A(clknet_5_12__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_43_clk_p2c (.X(clknet_leaf_43_clk_p2c),
    .A(clknet_5_12__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_44_clk_p2c (.X(clknet_leaf_44_clk_p2c),
    .A(clknet_5_12__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_45_clk_p2c (.X(clknet_leaf_45_clk_p2c),
    .A(clknet_5_12__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_46_clk_p2c (.X(clknet_leaf_46_clk_p2c),
    .A(clknet_5_12__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_47_clk_p2c (.X(clknet_leaf_47_clk_p2c),
    .A(clknet_5_12__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_48_clk_p2c (.X(clknet_leaf_48_clk_p2c),
    .A(clknet_5_11__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_49_clk_p2c (.X(clknet_leaf_49_clk_p2c),
    .A(clknet_5_9__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_50_clk_p2c (.X(clknet_leaf_50_clk_p2c),
    .A(clknet_5_9__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_51_clk_p2c (.X(clknet_leaf_51_clk_p2c),
    .A(clknet_5_9__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_52_clk_p2c (.X(clknet_leaf_52_clk_p2c),
    .A(clknet_5_9__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_53_clk_p2c (.X(clknet_leaf_53_clk_p2c),
    .A(clknet_5_9__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_54_clk_p2c (.X(clknet_leaf_54_clk_p2c),
    .A(clknet_5_9__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_55_clk_p2c (.X(clknet_leaf_55_clk_p2c),
    .A(clknet_5_9__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_56_clk_p2c (.X(clknet_leaf_56_clk_p2c),
    .A(clknet_5_8__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_57_clk_p2c (.X(clknet_leaf_57_clk_p2c),
    .A(clknet_5_8__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_58_clk_p2c (.X(clknet_leaf_58_clk_p2c),
    .A(clknet_5_8__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_59_clk_p2c (.X(clknet_leaf_59_clk_p2c),
    .A(clknet_5_8__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_60_clk_p2c (.X(clknet_leaf_60_clk_p2c),
    .A(clknet_5_8__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_61_clk_p2c (.X(clknet_leaf_61_clk_p2c),
    .A(clknet_5_8__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_62_clk_p2c (.X(clknet_leaf_62_clk_p2c),
    .A(clknet_5_8__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_63_clk_p2c (.X(clknet_leaf_63_clk_p2c),
    .A(clknet_5_10__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_64_clk_p2c (.X(clknet_leaf_64_clk_p2c),
    .A(clknet_5_10__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_65_clk_p2c (.X(clknet_leaf_65_clk_p2c),
    .A(clknet_5_8__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_66_clk_p2c (.X(clknet_leaf_66_clk_p2c),
    .A(clknet_5_11__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_67_clk_p2c (.X(clknet_leaf_67_clk_p2c),
    .A(clknet_5_11__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_68_clk_p2c (.X(clknet_leaf_68_clk_p2c),
    .A(clknet_5_11__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_69_clk_p2c (.X(clknet_leaf_69_clk_p2c),
    .A(clknet_5_11__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_70_clk_p2c (.X(clknet_leaf_70_clk_p2c),
    .A(clknet_5_10__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_71_clk_p2c (.X(clknet_leaf_71_clk_p2c),
    .A(clknet_5_11__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_72_clk_p2c (.X(clknet_leaf_72_clk_p2c),
    .A(clknet_5_10__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_73_clk_p2c (.X(clknet_leaf_73_clk_p2c),
    .A(clknet_5_10__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_74_clk_p2c (.X(clknet_leaf_74_clk_p2c),
    .A(clknet_5_10__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_75_clk_p2c (.X(clknet_leaf_75_clk_p2c),
    .A(clknet_5_10__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_76_clk_p2c (.X(clknet_leaf_76_clk_p2c),
    .A(clknet_5_10__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_77_clk_p2c (.X(clknet_leaf_77_clk_p2c),
    .A(clknet_5_10__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_78_clk_p2c (.X(clknet_leaf_78_clk_p2c),
    .A(clknet_5_10__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_79_clk_p2c (.X(clknet_leaf_79_clk_p2c),
    .A(clknet_5_10__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_80_clk_p2c (.X(clknet_leaf_80_clk_p2c),
    .A(clknet_5_10__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_81_clk_p2c (.X(clknet_leaf_81_clk_p2c),
    .A(clknet_5_11__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_82_clk_p2c (.X(clknet_leaf_82_clk_p2c),
    .A(clknet_5_11__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_83_clk_p2c (.X(clknet_leaf_83_clk_p2c),
    .A(clknet_5_14__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_84_clk_p2c (.X(clknet_leaf_84_clk_p2c),
    .A(clknet_5_14__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_85_clk_p2c (.X(clknet_leaf_85_clk_p2c),
    .A(clknet_5_14__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_86_clk_p2c (.X(clknet_leaf_86_clk_p2c),
    .A(clknet_5_14__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_87_clk_p2c (.X(clknet_leaf_87_clk_p2c),
    .A(clknet_5_15__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_88_clk_p2c (.X(clknet_leaf_88_clk_p2c),
    .A(clknet_5_15__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_89_clk_p2c (.X(clknet_leaf_89_clk_p2c),
    .A(clknet_5_15__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_90_clk_p2c (.X(clknet_leaf_90_clk_p2c),
    .A(clknet_5_15__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_91_clk_p2c (.X(clknet_leaf_91_clk_p2c),
    .A(clknet_5_15__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_92_clk_p2c (.X(clknet_leaf_92_clk_p2c),
    .A(clknet_5_15__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_93_clk_p2c (.X(clknet_leaf_93_clk_p2c),
    .A(clknet_5_14__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_94_clk_p2c (.X(clknet_leaf_94_clk_p2c),
    .A(clknet_5_14__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_95_clk_p2c (.X(clknet_leaf_95_clk_p2c),
    .A(clknet_5_14__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_96_clk_p2c (.X(clknet_leaf_96_clk_p2c),
    .A(clknet_5_14__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_97_clk_p2c (.X(clknet_leaf_97_clk_p2c),
    .A(clknet_5_14__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_98_clk_p2c (.X(clknet_leaf_98_clk_p2c),
    .A(clknet_5_13__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_99_clk_p2c (.X(clknet_leaf_99_clk_p2c),
    .A(clknet_5_15__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_100_clk_p2c (.X(clknet_leaf_100_clk_p2c),
    .A(clknet_5_15__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_101_clk_p2c (.X(clknet_leaf_101_clk_p2c),
    .A(clknet_5_15__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_102_clk_p2c (.X(clknet_leaf_102_clk_p2c),
    .A(clknet_5_15__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_103_clk_p2c (.X(clknet_leaf_103_clk_p2c),
    .A(clknet_5_24__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_104_clk_p2c (.X(clknet_leaf_104_clk_p2c),
    .A(clknet_5_13__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_105_clk_p2c (.X(clknet_leaf_105_clk_p2c),
    .A(clknet_5_13__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_106_clk_p2c (.X(clknet_leaf_106_clk_p2c),
    .A(clknet_5_13__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_107_clk_p2c (.X(clknet_leaf_107_clk_p2c),
    .A(clknet_5_13__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_108_clk_p2c (.X(clknet_leaf_108_clk_p2c),
    .A(clknet_5_24__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_109_clk_p2c (.X(clknet_leaf_109_clk_p2c),
    .A(clknet_5_24__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_110_clk_p2c (.X(clknet_leaf_110_clk_p2c),
    .A(clknet_5_24__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_111_clk_p2c (.X(clknet_leaf_111_clk_p2c),
    .A(clknet_5_24__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_112_clk_p2c (.X(clknet_leaf_112_clk_p2c),
    .A(clknet_5_24__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_113_clk_p2c (.X(clknet_leaf_113_clk_p2c),
    .A(clknet_5_26__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_114_clk_p2c (.X(clknet_leaf_114_clk_p2c),
    .A(clknet_5_26__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_115_clk_p2c (.X(clknet_leaf_115_clk_p2c),
    .A(clknet_5_25__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_116_clk_p2c (.X(clknet_leaf_116_clk_p2c),
    .A(clknet_5_25__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_117_clk_p2c (.X(clknet_leaf_117_clk_p2c),
    .A(clknet_5_27__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_118_clk_p2c (.X(clknet_leaf_118_clk_p2c),
    .A(clknet_5_27__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_119_clk_p2c (.X(clknet_leaf_119_clk_p2c),
    .A(clknet_5_27__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_120_clk_p2c (.X(clknet_leaf_120_clk_p2c),
    .A(clknet_5_26__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_121_clk_p2c (.X(clknet_leaf_121_clk_p2c),
    .A(clknet_5_26__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_122_clk_p2c (.X(clknet_leaf_122_clk_p2c),
    .A(clknet_5_26__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_123_clk_p2c (.X(clknet_leaf_123_clk_p2c),
    .A(clknet_5_26__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_124_clk_p2c (.X(clknet_leaf_124_clk_p2c),
    .A(clknet_5_27__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_125_clk_p2c (.X(clknet_leaf_125_clk_p2c),
    .A(clknet_5_26__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_126_clk_p2c (.X(clknet_leaf_126_clk_p2c),
    .A(clknet_5_26__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_127_clk_p2c (.X(clknet_leaf_127_clk_p2c),
    .A(clknet_5_27__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_128_clk_p2c (.X(clknet_leaf_128_clk_p2c),
    .A(clknet_5_27__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_129_clk_p2c (.X(clknet_leaf_129_clk_p2c),
    .A(clknet_5_27__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_130_clk_p2c (.X(clknet_leaf_130_clk_p2c),
    .A(clknet_5_27__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_131_clk_p2c (.X(clknet_leaf_131_clk_p2c),
    .A(clknet_5_30__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_132_clk_p2c (.X(clknet_leaf_132_clk_p2c),
    .A(clknet_5_30__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_133_clk_p2c (.X(clknet_leaf_133_clk_p2c),
    .A(clknet_5_27__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_134_clk_p2c (.X(clknet_leaf_134_clk_p2c),
    .A(clknet_5_30__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_135_clk_p2c (.X(clknet_leaf_135_clk_p2c),
    .A(clknet_5_30__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_136_clk_p2c (.X(clknet_leaf_136_clk_p2c),
    .A(clknet_5_31__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_137_clk_p2c (.X(clknet_leaf_137_clk_p2c),
    .A(clknet_5_31__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_138_clk_p2c (.X(clknet_leaf_138_clk_p2c),
    .A(clknet_5_31__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_139_clk_p2c (.X(clknet_leaf_139_clk_p2c),
    .A(clknet_5_31__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_140_clk_p2c (.X(clknet_leaf_140_clk_p2c),
    .A(clknet_5_31__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_141_clk_p2c (.X(clknet_leaf_141_clk_p2c),
    .A(clknet_5_31__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_142_clk_p2c (.X(clknet_leaf_142_clk_p2c),
    .A(clknet_5_31__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_143_clk_p2c (.X(clknet_leaf_143_clk_p2c),
    .A(clknet_5_30__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_144_clk_p2c (.X(clknet_leaf_144_clk_p2c),
    .A(clknet_5_29__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_145_clk_p2c (.X(clknet_leaf_145_clk_p2c),
    .A(clknet_5_29__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_146_clk_p2c (.X(clknet_leaf_146_clk_p2c),
    .A(clknet_5_29__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_147_clk_p2c (.X(clknet_leaf_147_clk_p2c),
    .A(clknet_5_29__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_148_clk_p2c (.X(clknet_leaf_148_clk_p2c),
    .A(clknet_5_29__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_149_clk_p2c (.X(clknet_leaf_149_clk_p2c),
    .A(clknet_5_29__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_150_clk_p2c (.X(clknet_leaf_150_clk_p2c),
    .A(clknet_5_29__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_151_clk_p2c (.X(clknet_leaf_151_clk_p2c),
    .A(clknet_5_28__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_152_clk_p2c (.X(clknet_leaf_152_clk_p2c),
    .A(clknet_5_28__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_153_clk_p2c (.X(clknet_leaf_153_clk_p2c),
    .A(clknet_5_28__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_154_clk_p2c (.X(clknet_leaf_154_clk_p2c),
    .A(clknet_5_29__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_155_clk_p2c (.X(clknet_leaf_155_clk_p2c),
    .A(clknet_5_29__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_156_clk_p2c (.X(clknet_leaf_156_clk_p2c),
    .A(clknet_5_28__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_157_clk_p2c (.X(clknet_leaf_157_clk_p2c),
    .A(clknet_5_28__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_158_clk_p2c (.X(clknet_leaf_158_clk_p2c),
    .A(clknet_5_28__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_159_clk_p2c (.X(clknet_leaf_159_clk_p2c),
    .A(clknet_5_25__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_160_clk_p2c (.X(clknet_leaf_160_clk_p2c),
    .A(clknet_5_25__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_161_clk_p2c (.X(clknet_leaf_161_clk_p2c),
    .A(clknet_5_28__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_162_clk_p2c (.X(clknet_leaf_162_clk_p2c),
    .A(clknet_5_28__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_163_clk_p2c (.X(clknet_leaf_163_clk_p2c),
    .A(clknet_5_25__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_164_clk_p2c (.X(clknet_leaf_164_clk_p2c),
    .A(clknet_5_25__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_165_clk_p2c (.X(clknet_leaf_165_clk_p2c),
    .A(clknet_5_25__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_166_clk_p2c (.X(clknet_leaf_166_clk_p2c),
    .A(clknet_5_25__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_167_clk_p2c (.X(clknet_leaf_167_clk_p2c),
    .A(clknet_5_24__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_168_clk_p2c (.X(clknet_leaf_168_clk_p2c),
    .A(clknet_5_24__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_169_clk_p2c (.X(clknet_leaf_169_clk_p2c),
    .A(clknet_5_24__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_170_clk_p2c (.X(clknet_leaf_170_clk_p2c),
    .A(clknet_5_19__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_171_clk_p2c (.X(clknet_leaf_171_clk_p2c),
    .A(clknet_5_19__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_172_clk_p2c (.X(clknet_leaf_172_clk_p2c),
    .A(clknet_5_25__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_173_clk_p2c (.X(clknet_leaf_173_clk_p2c),
    .A(clknet_5_19__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_174_clk_p2c (.X(clknet_leaf_174_clk_p2c),
    .A(clknet_5_22__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_175_clk_p2c (.X(clknet_leaf_175_clk_p2c),
    .A(clknet_5_19__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_176_clk_p2c (.X(clknet_leaf_176_clk_p2c),
    .A(clknet_5_19__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_177_clk_p2c (.X(clknet_leaf_177_clk_p2c),
    .A(clknet_5_19__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_178_clk_p2c (.X(clknet_leaf_178_clk_p2c),
    .A(clknet_5_22__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_179_clk_p2c (.X(clknet_leaf_179_clk_p2c),
    .A(clknet_5_22__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_180_clk_p2c (.X(clknet_leaf_180_clk_p2c),
    .A(clknet_5_22__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_181_clk_p2c (.X(clknet_leaf_181_clk_p2c),
    .A(clknet_5_22__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_182_clk_p2c (.X(clknet_leaf_182_clk_p2c),
    .A(clknet_5_23__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_183_clk_p2c (.X(clknet_leaf_183_clk_p2c),
    .A(clknet_5_23__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_184_clk_p2c (.X(clknet_leaf_184_clk_p2c),
    .A(clknet_5_22__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_185_clk_p2c (.X(clknet_leaf_185_clk_p2c),
    .A(clknet_5_22__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_186_clk_p2c (.X(clknet_leaf_186_clk_p2c),
    .A(clknet_5_23__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_187_clk_p2c (.X(clknet_leaf_187_clk_p2c),
    .A(clknet_5_23__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_188_clk_p2c (.X(clknet_leaf_188_clk_p2c),
    .A(clknet_5_23__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_189_clk_p2c (.X(clknet_leaf_189_clk_p2c),
    .A(clknet_5_21__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_190_clk_p2c (.X(clknet_leaf_190_clk_p2c),
    .A(clknet_5_21__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_191_clk_p2c (.X(clknet_leaf_191_clk_p2c),
    .A(clknet_5_23__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_192_clk_p2c (.X(clknet_leaf_192_clk_p2c),
    .A(clknet_5_23__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_193_clk_p2c (.X(clknet_leaf_193_clk_p2c),
    .A(clknet_5_22__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_194_clk_p2c (.X(clknet_leaf_194_clk_p2c),
    .A(clknet_5_23__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_195_clk_p2c (.X(clknet_leaf_195_clk_p2c),
    .A(clknet_5_20__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_196_clk_p2c (.X(clknet_leaf_196_clk_p2c),
    .A(clknet_5_21__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_197_clk_p2c (.X(clknet_leaf_197_clk_p2c),
    .A(clknet_5_21__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_198_clk_p2c (.X(clknet_leaf_198_clk_p2c),
    .A(clknet_5_21__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_199_clk_p2c (.X(clknet_leaf_199_clk_p2c),
    .A(clknet_5_21__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_200_clk_p2c (.X(clknet_leaf_200_clk_p2c),
    .A(clknet_5_21__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_201_clk_p2c (.X(clknet_leaf_201_clk_p2c),
    .A(clknet_5_21__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_202_clk_p2c (.X(clknet_leaf_202_clk_p2c),
    .A(clknet_5_21__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_203_clk_p2c (.X(clknet_leaf_203_clk_p2c),
    .A(clknet_5_21__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_204_clk_p2c (.X(clknet_leaf_204_clk_p2c),
    .A(clknet_5_21__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_205_clk_p2c (.X(clknet_leaf_205_clk_p2c),
    .A(clknet_5_21__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_206_clk_p2c (.X(clknet_leaf_206_clk_p2c),
    .A(clknet_5_21__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_207_clk_p2c (.X(clknet_leaf_207_clk_p2c),
    .A(clknet_5_20__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_208_clk_p2c (.X(clknet_leaf_208_clk_p2c),
    .A(clknet_5_20__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_209_clk_p2c (.X(clknet_leaf_209_clk_p2c),
    .A(clknet_5_20__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_210_clk_p2c (.X(clknet_leaf_210_clk_p2c),
    .A(clknet_5_20__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_211_clk_p2c (.X(clknet_leaf_211_clk_p2c),
    .A(clknet_5_20__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_212_clk_p2c (.X(clknet_leaf_212_clk_p2c),
    .A(clknet_5_20__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_213_clk_p2c (.X(clknet_leaf_213_clk_p2c),
    .A(clknet_5_20__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_214_clk_p2c (.X(clknet_leaf_214_clk_p2c),
    .A(clknet_5_17__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_215_clk_p2c (.X(clknet_leaf_215_clk_p2c),
    .A(clknet_5_17__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_216_clk_p2c (.X(clknet_leaf_216_clk_p2c),
    .A(clknet_5_17__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_217_clk_p2c (.X(clknet_leaf_217_clk_p2c),
    .A(clknet_5_20__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_218_clk_p2c (.X(clknet_leaf_218_clk_p2c),
    .A(clknet_5_17__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_219_clk_p2c (.X(clknet_leaf_219_clk_p2c),
    .A(clknet_5_17__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_220_clk_p2c (.X(clknet_leaf_220_clk_p2c),
    .A(clknet_5_16__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_221_clk_p2c (.X(clknet_leaf_221_clk_p2c),
    .A(clknet_5_16__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_222_clk_p2c (.X(clknet_leaf_222_clk_p2c),
    .A(clknet_5_16__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_223_clk_p2c (.X(clknet_leaf_223_clk_p2c),
    .A(clknet_5_16__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_224_clk_p2c (.X(clknet_leaf_224_clk_p2c),
    .A(clknet_5_16__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_225_clk_p2c (.X(clknet_leaf_225_clk_p2c),
    .A(clknet_5_16__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_226_clk_p2c (.X(clknet_leaf_226_clk_p2c),
    .A(clknet_5_16__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_227_clk_p2c (.X(clknet_leaf_227_clk_p2c),
    .A(clknet_5_16__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_228_clk_p2c (.X(clknet_leaf_228_clk_p2c),
    .A(clknet_5_16__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_229_clk_p2c (.X(clknet_leaf_229_clk_p2c),
    .A(clknet_5_17__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_230_clk_p2c (.X(clknet_leaf_230_clk_p2c),
    .A(clknet_5_17__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_231_clk_p2c (.X(clknet_leaf_231_clk_p2c),
    .A(clknet_5_17__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_232_clk_p2c (.X(clknet_leaf_232_clk_p2c),
    .A(clknet_5_19__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_233_clk_p2c (.X(clknet_leaf_233_clk_p2c),
    .A(clknet_5_19__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_234_clk_p2c (.X(clknet_leaf_234_clk_p2c),
    .A(clknet_5_19__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_235_clk_p2c (.X(clknet_leaf_235_clk_p2c),
    .A(clknet_5_18__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_236_clk_p2c (.X(clknet_leaf_236_clk_p2c),
    .A(clknet_5_18__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_237_clk_p2c (.X(clknet_leaf_237_clk_p2c),
    .A(clknet_5_18__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_238_clk_p2c (.X(clknet_leaf_238_clk_p2c),
    .A(clknet_5_18__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_239_clk_p2c (.X(clknet_leaf_239_clk_p2c),
    .A(clknet_5_18__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_240_clk_p2c (.X(clknet_leaf_240_clk_p2c),
    .A(clknet_5_18__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_241_clk_p2c (.X(clknet_leaf_241_clk_p2c),
    .A(clknet_5_18__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_242_clk_p2c (.X(clknet_leaf_242_clk_p2c),
    .A(clknet_5_18__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_243_clk_p2c (.X(clknet_leaf_243_clk_p2c),
    .A(clknet_5_18__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_244_clk_p2c (.X(clknet_leaf_244_clk_p2c),
    .A(clknet_5_7__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_245_clk_p2c (.X(clknet_leaf_245_clk_p2c),
    .A(clknet_5_7__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_246_clk_p2c (.X(clknet_leaf_246_clk_p2c),
    .A(clknet_5_7__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_247_clk_p2c (.X(clknet_leaf_247_clk_p2c),
    .A(clknet_5_7__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_248_clk_p2c (.X(clknet_leaf_248_clk_p2c),
    .A(clknet_5_7__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_249_clk_p2c (.X(clknet_leaf_249_clk_p2c),
    .A(clknet_5_7__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_250_clk_p2c (.X(clknet_leaf_250_clk_p2c),
    .A(clknet_5_7__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_251_clk_p2c (.X(clknet_leaf_251_clk_p2c),
    .A(clknet_5_7__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_252_clk_p2c (.X(clknet_leaf_252_clk_p2c),
    .A(clknet_5_6__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_253_clk_p2c (.X(clknet_leaf_253_clk_p2c),
    .A(clknet_5_6__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_254_clk_p2c (.X(clknet_leaf_254_clk_p2c),
    .A(clknet_5_6__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_255_clk_p2c (.X(clknet_leaf_255_clk_p2c),
    .A(clknet_5_4__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_256_clk_p2c (.X(clknet_leaf_256_clk_p2c),
    .A(clknet_5_4__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_257_clk_p2c (.X(clknet_leaf_257_clk_p2c),
    .A(clknet_5_4__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_258_clk_p2c (.X(clknet_leaf_258_clk_p2c),
    .A(clknet_5_5__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_259_clk_p2c (.X(clknet_leaf_259_clk_p2c),
    .A(clknet_5_5__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_260_clk_p2c (.X(clknet_leaf_260_clk_p2c),
    .A(clknet_5_5__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_261_clk_p2c (.X(clknet_leaf_261_clk_p2c),
    .A(clknet_5_5__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_262_clk_p2c (.X(clknet_leaf_262_clk_p2c),
    .A(clknet_5_5__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_263_clk_p2c (.X(clknet_leaf_263_clk_p2c),
    .A(clknet_5_5__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_264_clk_p2c (.X(clknet_leaf_264_clk_p2c),
    .A(clknet_5_5__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_265_clk_p2c (.X(clknet_leaf_265_clk_p2c),
    .A(clknet_5_5__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_266_clk_p2c (.X(clknet_leaf_266_clk_p2c),
    .A(clknet_5_5__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_267_clk_p2c (.X(clknet_leaf_267_clk_p2c),
    .A(clknet_5_5__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_268_clk_p2c (.X(clknet_leaf_268_clk_p2c),
    .A(clknet_5_5__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_269_clk_p2c (.X(clknet_leaf_269_clk_p2c),
    .A(clknet_5_4__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_270_clk_p2c (.X(clknet_leaf_270_clk_p2c),
    .A(clknet_5_4__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_271_clk_p2c (.X(clknet_leaf_271_clk_p2c),
    .A(clknet_5_4__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_272_clk_p2c (.X(clknet_leaf_272_clk_p2c),
    .A(clknet_5_4__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_273_clk_p2c (.X(clknet_leaf_273_clk_p2c),
    .A(clknet_5_1__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_274_clk_p2c (.X(clknet_leaf_274_clk_p2c),
    .A(clknet_5_4__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_275_clk_p2c (.X(clknet_leaf_275_clk_p2c),
    .A(clknet_5_4__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_276_clk_p2c (.X(clknet_leaf_276_clk_p2c),
    .A(clknet_5_4__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_277_clk_p2c (.X(clknet_leaf_277_clk_p2c),
    .A(clknet_5_4__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_278_clk_p2c (.X(clknet_leaf_278_clk_p2c),
    .A(clknet_5_1__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_279_clk_p2c (.X(clknet_leaf_279_clk_p2c),
    .A(clknet_5_1__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_280_clk_p2c (.X(clknet_leaf_280_clk_p2c),
    .A(clknet_5_1__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_281_clk_p2c (.X(clknet_leaf_281_clk_p2c),
    .A(clknet_5_1__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_282_clk_p2c (.X(clknet_leaf_282_clk_p2c),
    .A(clknet_5_1__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_283_clk_p2c (.X(clknet_leaf_283_clk_p2c),
    .A(clknet_5_1__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_284_clk_p2c (.X(clknet_leaf_284_clk_p2c),
    .A(clknet_5_1__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_285_clk_p2c (.X(clknet_leaf_285_clk_p2c),
    .A(clknet_5_1__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_286_clk_p2c (.X(clknet_leaf_286_clk_p2c),
    .A(clknet_5_0__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_287_clk_p2c (.X(clknet_leaf_287_clk_p2c),
    .A(clknet_5_0__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_288_clk_p2c (.X(clknet_leaf_288_clk_p2c),
    .A(clknet_5_0__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_289_clk_p2c (.X(clknet_leaf_289_clk_p2c),
    .A(clknet_5_0__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_290_clk_p2c (.X(clknet_leaf_290_clk_p2c),
    .A(clknet_5_0__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_291_clk_p2c (.X(clknet_leaf_291_clk_p2c),
    .A(clknet_5_0__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_292_clk_p2c (.X(clknet_leaf_292_clk_p2c),
    .A(clknet_5_0__leaf_clk_p2c));
 sg13g2_buf_4 clkbuf_leaf_293_clk_p2c (.X(clknet_leaf_293_clk_p2c),
    .A(clknet_5_0__leaf_clk_p2c));
 sg13g2_buf_2 clkbuf_0_clk_p2c (.A(clk_p2c),
    .X(clknet_0_clk_p2c));
 sg13g2_buf_4 clkbuf_4_0_0_clk_p2c (.X(clknet_4_0_0_clk_p2c),
    .A(clknet_0_clk_p2c));
 sg13g2_buf_4 clkbuf_4_1_0_clk_p2c (.X(clknet_4_1_0_clk_p2c),
    .A(clknet_0_clk_p2c));
 sg13g2_buf_4 clkbuf_4_2_0_clk_p2c (.X(clknet_4_2_0_clk_p2c),
    .A(clknet_0_clk_p2c));
 sg13g2_buf_4 clkbuf_4_3_0_clk_p2c (.X(clknet_4_3_0_clk_p2c),
    .A(clknet_0_clk_p2c));
 sg13g2_buf_4 clkbuf_4_4_0_clk_p2c (.X(clknet_4_4_0_clk_p2c),
    .A(clknet_0_clk_p2c));
 sg13g2_buf_4 clkbuf_4_5_0_clk_p2c (.X(clknet_4_5_0_clk_p2c),
    .A(clknet_0_clk_p2c));
 sg13g2_buf_4 clkbuf_4_6_0_clk_p2c (.X(clknet_4_6_0_clk_p2c),
    .A(clknet_0_clk_p2c));
 sg13g2_buf_4 clkbuf_4_7_0_clk_p2c (.X(clknet_4_7_0_clk_p2c),
    .A(clknet_0_clk_p2c));
 sg13g2_buf_4 clkbuf_4_8_0_clk_p2c (.X(clknet_4_8_0_clk_p2c),
    .A(clknet_0_clk_p2c));
 sg13g2_buf_4 clkbuf_4_9_0_clk_p2c (.X(clknet_4_9_0_clk_p2c),
    .A(clknet_0_clk_p2c));
 sg13g2_buf_4 clkbuf_4_10_0_clk_p2c (.X(clknet_4_10_0_clk_p2c),
    .A(clknet_0_clk_p2c));
 sg13g2_buf_4 clkbuf_4_11_0_clk_p2c (.X(clknet_4_11_0_clk_p2c),
    .A(clknet_0_clk_p2c));
 sg13g2_buf_4 clkbuf_4_12_0_clk_p2c (.X(clknet_4_12_0_clk_p2c),
    .A(clknet_0_clk_p2c));
 sg13g2_buf_4 clkbuf_4_13_0_clk_p2c (.X(clknet_4_13_0_clk_p2c),
    .A(clknet_0_clk_p2c));
 sg13g2_buf_4 clkbuf_4_14_0_clk_p2c (.X(clknet_4_14_0_clk_p2c),
    .A(clknet_0_clk_p2c));
 sg13g2_buf_4 clkbuf_4_15_0_clk_p2c (.X(clknet_4_15_0_clk_p2c),
    .A(clknet_0_clk_p2c));
 sg13g2_buf_2 clkbuf_5_0__f_clk_p2c (.A(clknet_4_0_0_clk_p2c),
    .X(clknet_5_0__leaf_clk_p2c));
 sg13g2_buf_2 clkbuf_5_1__f_clk_p2c (.A(clknet_4_0_0_clk_p2c),
    .X(clknet_5_1__leaf_clk_p2c));
 sg13g2_buf_2 clkbuf_5_2__f_clk_p2c (.A(clknet_4_1_0_clk_p2c),
    .X(clknet_5_2__leaf_clk_p2c));
 sg13g2_buf_2 clkbuf_5_3__f_clk_p2c (.A(clknet_4_1_0_clk_p2c),
    .X(clknet_5_3__leaf_clk_p2c));
 sg13g2_buf_2 clkbuf_5_4__f_clk_p2c (.A(clknet_4_2_0_clk_p2c),
    .X(clknet_5_4__leaf_clk_p2c));
 sg13g2_buf_2 clkbuf_5_5__f_clk_p2c (.A(clknet_4_2_0_clk_p2c),
    .X(clknet_5_5__leaf_clk_p2c));
 sg13g2_buf_2 clkbuf_5_6__f_clk_p2c (.A(clknet_4_3_0_clk_p2c),
    .X(clknet_5_6__leaf_clk_p2c));
 sg13g2_buf_2 clkbuf_5_7__f_clk_p2c (.A(clknet_4_3_0_clk_p2c),
    .X(clknet_5_7__leaf_clk_p2c));
 sg13g2_buf_2 clkbuf_5_8__f_clk_p2c (.A(clknet_4_4_0_clk_p2c),
    .X(clknet_5_8__leaf_clk_p2c));
 sg13g2_buf_2 clkbuf_5_9__f_clk_p2c (.A(clknet_4_4_0_clk_p2c),
    .X(clknet_5_9__leaf_clk_p2c));
 sg13g2_buf_2 clkbuf_5_10__f_clk_p2c (.A(clknet_4_5_0_clk_p2c),
    .X(clknet_5_10__leaf_clk_p2c));
 sg13g2_buf_2 clkbuf_5_11__f_clk_p2c (.A(clknet_4_5_0_clk_p2c),
    .X(clknet_5_11__leaf_clk_p2c));
 sg13g2_buf_2 clkbuf_5_12__f_clk_p2c (.A(clknet_4_6_0_clk_p2c),
    .X(clknet_5_12__leaf_clk_p2c));
 sg13g2_buf_2 clkbuf_5_13__f_clk_p2c (.A(clknet_4_6_0_clk_p2c),
    .X(clknet_5_13__leaf_clk_p2c));
 sg13g2_buf_2 clkbuf_5_14__f_clk_p2c (.A(clknet_4_7_0_clk_p2c),
    .X(clknet_5_14__leaf_clk_p2c));
 sg13g2_buf_2 clkbuf_5_15__f_clk_p2c (.A(clknet_4_7_0_clk_p2c),
    .X(clknet_5_15__leaf_clk_p2c));
 sg13g2_buf_2 clkbuf_5_16__f_clk_p2c (.A(clknet_4_8_0_clk_p2c),
    .X(clknet_5_16__leaf_clk_p2c));
 sg13g2_buf_2 clkbuf_5_17__f_clk_p2c (.A(clknet_4_8_0_clk_p2c),
    .X(clknet_5_17__leaf_clk_p2c));
 sg13g2_buf_2 clkbuf_5_18__f_clk_p2c (.A(clknet_4_9_0_clk_p2c),
    .X(clknet_5_18__leaf_clk_p2c));
 sg13g2_buf_2 clkbuf_5_19__f_clk_p2c (.A(clknet_4_9_0_clk_p2c),
    .X(clknet_5_19__leaf_clk_p2c));
 sg13g2_buf_2 clkbuf_5_20__f_clk_p2c (.A(clknet_4_10_0_clk_p2c),
    .X(clknet_5_20__leaf_clk_p2c));
 sg13g2_buf_2 clkbuf_5_21__f_clk_p2c (.A(clknet_4_10_0_clk_p2c),
    .X(clknet_5_21__leaf_clk_p2c));
 sg13g2_buf_2 clkbuf_5_22__f_clk_p2c (.A(clknet_4_11_0_clk_p2c),
    .X(clknet_5_22__leaf_clk_p2c));
 sg13g2_buf_2 clkbuf_5_23__f_clk_p2c (.A(clknet_4_11_0_clk_p2c),
    .X(clknet_5_23__leaf_clk_p2c));
 sg13g2_buf_2 clkbuf_5_24__f_clk_p2c (.A(clknet_4_12_0_clk_p2c),
    .X(clknet_5_24__leaf_clk_p2c));
 sg13g2_buf_2 clkbuf_5_25__f_clk_p2c (.A(clknet_4_12_0_clk_p2c),
    .X(clknet_5_25__leaf_clk_p2c));
 sg13g2_buf_2 clkbuf_5_26__f_clk_p2c (.A(clknet_4_13_0_clk_p2c),
    .X(clknet_5_26__leaf_clk_p2c));
 sg13g2_buf_2 clkbuf_5_27__f_clk_p2c (.A(clknet_4_13_0_clk_p2c),
    .X(clknet_5_27__leaf_clk_p2c));
 sg13g2_buf_2 clkbuf_5_28__f_clk_p2c (.A(clknet_4_14_0_clk_p2c),
    .X(clknet_5_28__leaf_clk_p2c));
 sg13g2_buf_2 clkbuf_5_29__f_clk_p2c (.A(clknet_4_14_0_clk_p2c),
    .X(clknet_5_29__leaf_clk_p2c));
 sg13g2_buf_2 clkbuf_5_30__f_clk_p2c (.A(clknet_4_15_0_clk_p2c),
    .X(clknet_5_30__leaf_clk_p2c));
 sg13g2_buf_2 clkbuf_5_31__f_clk_p2c (.A(clknet_4_15_0_clk_p2c),
    .X(clknet_5_31__leaf_clk_p2c));
 sg13g2_buf_4 clkload0 (.A(clknet_5_3__leaf_clk_p2c));
 sg13g2_buf_4 clkload1 (.A(clknet_5_6__leaf_clk_p2c));
 sg13g2_buf_8 clkload2 (.A(clknet_5_9__leaf_clk_p2c));
 sg13g2_buf_16 clkload3 (.A(clknet_5_11__leaf_clk_p2c));
 sg13g2_buf_4 clkload4 (.A(clknet_5_14__leaf_clk_p2c));
 sg13g2_buf_4 clkload5 (.A(clknet_5_17__leaf_clk_p2c));
 sg13g2_buf_16 clkload6 (.A(clknet_5_20__leaf_clk_p2c));
 sg13g2_buf_4 clkload7 (.A(clknet_5_26__leaf_clk_p2c));
 sg13g2_buf_4 clkload8 (.A(clknet_5_28__leaf_clk_p2c));
 sg13g2_buf_8 clkload9 (.A(clknet_5_30__leaf_clk_p2c));
 sg13g2_inv_1 clkload10 (.A(clknet_leaf_2_clk_p2c));
 sg13g2_inv_2 clkload11 (.A(clknet_leaf_287_clk_p2c));
 sg13g2_inv_1 clkload12 (.A(clknet_leaf_288_clk_p2c));
 sg13g2_inv_1 clkload13 (.A(clknet_leaf_289_clk_p2c));
 sg13g2_inv_1 clkload14 (.A(clknet_leaf_290_clk_p2c));
 sg13g2_inv_2 clkload15 (.A(clknet_leaf_291_clk_p2c));
 sg13g2_inv_1 clkload16 (.A(clknet_leaf_292_clk_p2c));
 sg13g2_inv_1 clkload17 (.A(clknet_leaf_293_clk_p2c));
 sg13g2_inv_2 clkload18 (.A(clknet_leaf_3_clk_p2c));
 sg13g2_inv_1 clkload19 (.A(clknet_leaf_4_clk_p2c));
 sg13g2_inv_2 clkload20 (.A(clknet_leaf_273_clk_p2c));
 sg13g2_inv_1 clkload21 (.A(clknet_leaf_279_clk_p2c));
 sg13g2_inv_1 clkload22 (.A(clknet_leaf_280_clk_p2c));
 sg13g2_inv_2 clkload23 (.A(clknet_leaf_281_clk_p2c));
 sg13g2_inv_1 clkload24 (.A(clknet_leaf_282_clk_p2c));
 sg13g2_inv_1 clkload25 (.A(clknet_leaf_283_clk_p2c));
 sg13g2_inv_1 clkload26 (.A(clknet_leaf_284_clk_p2c));
 sg13g2_inv_1 clkload27 (.A(clknet_leaf_285_clk_p2c));
 sg13g2_inv_1 clkload28 (.A(clknet_leaf_6_clk_p2c));
 sg13g2_inv_1 clkload29 (.A(clknet_leaf_8_clk_p2c));
 sg13g2_inv_1 clkload30 (.A(clknet_leaf_5_clk_p2c));
 sg13g2_inv_1 clkload31 (.A(clknet_leaf_18_clk_p2c));
 sg13g2_inv_2 clkload32 (.A(clknet_leaf_22_clk_p2c));
 sg13g2_inv_1 clkload33 (.A(clknet_leaf_23_clk_p2c));
 sg13g2_inv_2 clkload34 (.A(clknet_leaf_24_clk_p2c));
 sg13g2_buf_8 clkload35 (.A(clknet_leaf_25_clk_p2c));
 sg13g2_inv_1 clkload36 (.A(clknet_leaf_30_clk_p2c));
 sg13g2_inv_1 clkload37 (.A(clknet_leaf_255_clk_p2c));
 sg13g2_inv_1 clkload38 (.A(clknet_leaf_256_clk_p2c));
 sg13g2_inv_1 clkload39 (.A(clknet_leaf_257_clk_p2c));
 sg13g2_inv_2 clkload40 (.A(clknet_leaf_270_clk_p2c));
 sg13g2_inv_1 clkload41 (.A(clknet_leaf_271_clk_p2c));
 sg13g2_inv_1 clkload42 (.A(clknet_leaf_272_clk_p2c));
 sg13g2_inv_1 clkload43 (.A(clknet_leaf_274_clk_p2c));
 sg13g2_inv_1 clkload44 (.A(clknet_leaf_275_clk_p2c));
 sg13g2_inv_1 clkload45 (.A(clknet_leaf_276_clk_p2c));
 sg13g2_inv_1 clkload46 (.A(clknet_leaf_259_clk_p2c));
 sg13g2_inv_1 clkload47 (.A(clknet_leaf_260_clk_p2c));
 sg13g2_inv_1 clkload48 (.A(clknet_leaf_262_clk_p2c));
 sg13g2_inv_1 clkload49 (.A(clknet_leaf_263_clk_p2c));
 sg13g2_inv_1 clkload50 (.A(clknet_leaf_266_clk_p2c));
 sg13g2_inv_1 clkload51 (.A(clknet_leaf_268_clk_p2c));
 sg13g2_inv_1 clkload52 (.A(clknet_leaf_26_clk_p2c));
 sg13g2_inv_1 clkload53 (.A(clknet_leaf_27_clk_p2c));
 sg13g2_inv_1 clkload54 (.A(clknet_leaf_28_clk_p2c));
 sg13g2_inv_1 clkload55 (.A(clknet_leaf_29_clk_p2c));
 sg13g2_inv_1 clkload56 (.A(clknet_leaf_253_clk_p2c));
 sg13g2_inv_1 clkload57 (.A(clknet_leaf_254_clk_p2c));
 sg13g2_inv_1 clkload58 (.A(clknet_leaf_33_clk_p2c));
 sg13g2_inv_2 clkload59 (.A(clknet_leaf_244_clk_p2c));
 sg13g2_inv_1 clkload60 (.A(clknet_leaf_245_clk_p2c));
 sg13g2_inv_2 clkload61 (.A(clknet_leaf_246_clk_p2c));
 sg13g2_inv_1 clkload62 (.A(clknet_leaf_247_clk_p2c));
 sg13g2_inv_1 clkload63 (.A(clknet_leaf_248_clk_p2c));
 sg13g2_inv_1 clkload64 (.A(clknet_leaf_251_clk_p2c));
 sg13g2_inv_1 clkload65 (.A(clknet_leaf_16_clk_p2c));
 sg13g2_inv_1 clkload66 (.A(clknet_leaf_57_clk_p2c));
 sg13g2_inv_1 clkload67 (.A(clknet_leaf_59_clk_p2c));
 sg13g2_inv_1 clkload68 (.A(clknet_leaf_19_clk_p2c));
 sg13g2_inv_1 clkload69 (.A(clknet_leaf_20_clk_p2c));
 sg13g2_inv_1 clkload70 (.A(clknet_leaf_49_clk_p2c));
 sg13g2_inv_1 clkload71 (.A(clknet_leaf_50_clk_p2c));
 sg13g2_inv_1 clkload72 (.A(clknet_leaf_51_clk_p2c));
 sg13g2_inv_2 clkload73 (.A(clknet_leaf_54_clk_p2c));
 sg13g2_inv_2 clkload74 (.A(clknet_leaf_63_clk_p2c));
 sg13g2_inv_2 clkload75 (.A(clknet_leaf_64_clk_p2c));
 sg13g2_inv_1 clkload76 (.A(clknet_leaf_70_clk_p2c));
 sg13g2_buf_8 clkload77 (.A(clknet_leaf_72_clk_p2c));
 sg13g2_inv_1 clkload78 (.A(clknet_leaf_73_clk_p2c));
 sg13g2_inv_1 clkload79 (.A(clknet_leaf_74_clk_p2c));
 sg13g2_inv_1 clkload80 (.A(clknet_leaf_75_clk_p2c));
 sg13g2_inv_1 clkload81 (.A(clknet_leaf_76_clk_p2c));
 sg13g2_inv_1 clkload82 (.A(clknet_leaf_77_clk_p2c));
 sg13g2_inv_1 clkload83 (.A(clknet_leaf_79_clk_p2c));
 sg13g2_inv_1 clkload84 (.A(clknet_leaf_80_clk_p2c));
 sg13g2_inv_1 clkload85 (.A(clknet_leaf_48_clk_p2c));
 sg13g2_inv_1 clkload86 (.A(clknet_leaf_66_clk_p2c));
 sg13g2_inv_1 clkload87 (.A(clknet_leaf_67_clk_p2c));
 sg13g2_inv_1 clkload88 (.A(clknet_leaf_69_clk_p2c));
 sg13g2_inv_1 clkload89 (.A(clknet_leaf_71_clk_p2c));
 sg13g2_inv_1 clkload90 (.A(clknet_leaf_81_clk_p2c));
 sg13g2_buf_8 clkload91 (.A(clknet_leaf_82_clk_p2c));
 sg13g2_inv_1 clkload92 (.A(clknet_leaf_39_clk_p2c));
 sg13g2_inv_2 clkload93 (.A(clknet_leaf_40_clk_p2c));
 sg13g2_inv_1 clkload94 (.A(clknet_leaf_41_clk_p2c));
 sg13g2_inv_1 clkload95 (.A(clknet_leaf_42_clk_p2c));
 sg13g2_inv_2 clkload96 (.A(clknet_leaf_43_clk_p2c));
 sg13g2_inv_1 clkload97 (.A(clknet_leaf_44_clk_p2c));
 sg13g2_inv_2 clkload98 (.A(clknet_leaf_45_clk_p2c));
 sg13g2_inv_1 clkload99 (.A(clknet_leaf_46_clk_p2c));
 sg13g2_inv_2 clkload100 (.A(clknet_leaf_47_clk_p2c));
 sg13g2_inv_1 clkload101 (.A(clknet_leaf_34_clk_p2c));
 sg13g2_inv_1 clkload102 (.A(clknet_leaf_35_clk_p2c));
 sg13g2_inv_1 clkload103 (.A(clknet_leaf_36_clk_p2c));
 sg13g2_inv_1 clkload104 (.A(clknet_leaf_37_clk_p2c));
 sg13g2_inv_1 clkload105 (.A(clknet_leaf_38_clk_p2c));
 sg13g2_inv_1 clkload106 (.A(clknet_leaf_98_clk_p2c));
 sg13g2_inv_1 clkload107 (.A(clknet_leaf_104_clk_p2c));
 sg13g2_inv_2 clkload108 (.A(clknet_leaf_105_clk_p2c));
 sg13g2_inv_2 clkload109 (.A(clknet_leaf_106_clk_p2c));
 sg13g2_inv_1 clkload110 (.A(clknet_leaf_83_clk_p2c));
 sg13g2_inv_2 clkload111 (.A(clknet_leaf_84_clk_p2c));
 sg13g2_inv_1 clkload112 (.A(clknet_leaf_85_clk_p2c));
 sg13g2_buf_8 clkload113 (.A(clknet_leaf_86_clk_p2c));
 sg13g2_inv_1 clkload114 (.A(clknet_leaf_93_clk_p2c));
 sg13g2_inv_2 clkload115 (.A(clknet_leaf_94_clk_p2c));
 sg13g2_inv_1 clkload116 (.A(clknet_leaf_95_clk_p2c));
 sg13g2_inv_1 clkload117 (.A(clknet_leaf_96_clk_p2c));
 sg13g2_inv_1 clkload118 (.A(clknet_leaf_99_clk_p2c));
 sg13g2_inv_1 clkload119 (.A(clknet_leaf_101_clk_p2c));
 sg13g2_inv_2 clkload120 (.A(clknet_leaf_220_clk_p2c));
 sg13g2_inv_1 clkload121 (.A(clknet_leaf_221_clk_p2c));
 sg13g2_inv_2 clkload122 (.A(clknet_leaf_222_clk_p2c));
 sg13g2_inv_1 clkload123 (.A(clknet_leaf_223_clk_p2c));
 sg13g2_inv_1 clkload124 (.A(clknet_leaf_224_clk_p2c));
 sg13g2_inv_2 clkload125 (.A(clknet_leaf_225_clk_p2c));
 sg13g2_inv_2 clkload126 (.A(clknet_leaf_228_clk_p2c));
 sg13g2_inv_1 clkload127 (.A(clknet_leaf_214_clk_p2c));
 sg13g2_inv_1 clkload128 (.A(clknet_leaf_216_clk_p2c));
 sg13g2_inv_2 clkload129 (.A(clknet_leaf_218_clk_p2c));
 sg13g2_inv_1 clkload130 (.A(clknet_leaf_219_clk_p2c));
 sg13g2_inv_1 clkload131 (.A(clknet_leaf_229_clk_p2c));
 sg13g2_inv_1 clkload132 (.A(clknet_leaf_230_clk_p2c));
 sg13g2_inv_1 clkload133 (.A(clknet_leaf_231_clk_p2c));
 sg13g2_inv_1 clkload134 (.A(clknet_leaf_235_clk_p2c));
 sg13g2_inv_2 clkload135 (.A(clknet_leaf_236_clk_p2c));
 sg13g2_inv_1 clkload136 (.A(clknet_leaf_237_clk_p2c));
 sg13g2_inv_1 clkload137 (.A(clknet_leaf_239_clk_p2c));
 sg13g2_inv_1 clkload138 (.A(clknet_leaf_240_clk_p2c));
 sg13g2_inv_1 clkload139 (.A(clknet_leaf_241_clk_p2c));
 sg13g2_inv_1 clkload140 (.A(clknet_leaf_242_clk_p2c));
 sg13g2_inv_1 clkload141 (.A(clknet_leaf_243_clk_p2c));
 sg13g2_inv_1 clkload142 (.A(clknet_leaf_170_clk_p2c));
 sg13g2_inv_1 clkload143 (.A(clknet_leaf_171_clk_p2c));
 sg13g2_inv_1 clkload144 (.A(clknet_leaf_173_clk_p2c));
 sg13g2_inv_2 clkload145 (.A(clknet_leaf_175_clk_p2c));
 sg13g2_inv_1 clkload146 (.A(clknet_leaf_232_clk_p2c));
 sg13g2_inv_1 clkload147 (.A(clknet_leaf_233_clk_p2c));
 sg13g2_buf_8 clkload148 (.A(clknet_leaf_234_clk_p2c));
 sg13g2_inv_1 clkload149 (.A(clknet_leaf_207_clk_p2c));
 sg13g2_inv_2 clkload150 (.A(clknet_leaf_208_clk_p2c));
 sg13g2_inv_1 clkload151 (.A(clknet_leaf_209_clk_p2c));
 sg13g2_inv_2 clkload152 (.A(clknet_leaf_210_clk_p2c));
 sg13g2_inv_1 clkload153 (.A(clknet_leaf_212_clk_p2c));
 sg13g2_inv_1 clkload154 (.A(clknet_leaf_213_clk_p2c));
 sg13g2_inv_2 clkload155 (.A(clknet_leaf_217_clk_p2c));
 sg13g2_inv_1 clkload156 (.A(clknet_leaf_196_clk_p2c));
 sg13g2_inv_1 clkload157 (.A(clknet_leaf_197_clk_p2c));
 sg13g2_inv_1 clkload158 (.A(clknet_leaf_199_clk_p2c));
 sg13g2_inv_2 clkload159 (.A(clknet_leaf_200_clk_p2c));
 sg13g2_inv_1 clkload160 (.A(clknet_leaf_201_clk_p2c));
 sg13g2_inv_1 clkload161 (.A(clknet_leaf_202_clk_p2c));
 sg13g2_inv_2 clkload162 (.A(clknet_leaf_203_clk_p2c));
 sg13g2_inv_1 clkload163 (.A(clknet_leaf_204_clk_p2c));
 sg13g2_inv_1 clkload164 (.A(clknet_leaf_205_clk_p2c));
 sg13g2_inv_1 clkload165 (.A(clknet_leaf_206_clk_p2c));
 sg13g2_inv_1 clkload166 (.A(clknet_leaf_178_clk_p2c));
 sg13g2_inv_1 clkload167 (.A(clknet_leaf_179_clk_p2c));
 sg13g2_inv_1 clkload168 (.A(clknet_leaf_180_clk_p2c));
 sg13g2_inv_2 clkload169 (.A(clknet_leaf_181_clk_p2c));
 sg13g2_inv_1 clkload170 (.A(clknet_leaf_184_clk_p2c));
 sg13g2_inv_2 clkload171 (.A(clknet_leaf_185_clk_p2c));
 sg13g2_inv_1 clkload172 (.A(clknet_leaf_193_clk_p2c));
 sg13g2_inv_2 clkload173 (.A(clknet_leaf_182_clk_p2c));
 sg13g2_inv_1 clkload174 (.A(clknet_leaf_186_clk_p2c));
 sg13g2_inv_1 clkload175 (.A(clknet_leaf_187_clk_p2c));
 sg13g2_buf_8 clkload176 (.A(clknet_leaf_188_clk_p2c));
 sg13g2_inv_1 clkload177 (.A(clknet_leaf_191_clk_p2c));
 sg13g2_inv_1 clkload178 (.A(clknet_leaf_192_clk_p2c));
 sg13g2_inv_2 clkload179 (.A(clknet_leaf_194_clk_p2c));
 sg13g2_inv_1 clkload180 (.A(clknet_leaf_103_clk_p2c));
 sg13g2_inv_1 clkload181 (.A(clknet_leaf_108_clk_p2c));
 sg13g2_inv_1 clkload182 (.A(clknet_leaf_110_clk_p2c));
 sg13g2_inv_1 clkload183 (.A(clknet_leaf_111_clk_p2c));
 sg13g2_inv_1 clkload184 (.A(clknet_leaf_112_clk_p2c));
 sg13g2_inv_1 clkload185 (.A(clknet_leaf_168_clk_p2c));
 sg13g2_inv_1 clkload186 (.A(clknet_leaf_169_clk_p2c));
 sg13g2_inv_1 clkload187 (.A(clknet_leaf_116_clk_p2c));
 sg13g2_inv_1 clkload188 (.A(clknet_leaf_159_clk_p2c));
 sg13g2_inv_1 clkload189 (.A(clknet_leaf_160_clk_p2c));
 sg13g2_inv_1 clkload190 (.A(clknet_leaf_165_clk_p2c));
 sg13g2_inv_1 clkload191 (.A(clknet_leaf_113_clk_p2c));
 sg13g2_inv_1 clkload192 (.A(clknet_leaf_121_clk_p2c));
 sg13g2_buf_8 clkload193 (.A(clknet_leaf_122_clk_p2c));
 sg13g2_inv_1 clkload194 (.A(clknet_leaf_123_clk_p2c));
 sg13g2_inv_1 clkload195 (.A(clknet_leaf_125_clk_p2c));
 sg13g2_inv_1 clkload196 (.A(clknet_leaf_126_clk_p2c));
 sg13g2_inv_1 clkload197 (.A(clknet_leaf_117_clk_p2c));
 sg13g2_inv_2 clkload198 (.A(clknet_leaf_118_clk_p2c));
 sg13g2_inv_2 clkload199 (.A(clknet_leaf_119_clk_p2c));
 sg13g2_inv_1 clkload200 (.A(clknet_leaf_124_clk_p2c));
 sg13g2_inv_1 clkload201 (.A(clknet_leaf_127_clk_p2c));
 sg13g2_inv_1 clkload202 (.A(clknet_leaf_129_clk_p2c));
 sg13g2_inv_2 clkload203 (.A(clknet_leaf_130_clk_p2c));
 sg13g2_buf_16 clkload204 (.A(clknet_leaf_133_clk_p2c));
 sg13g2_inv_1 clkload205 (.A(clknet_leaf_152_clk_p2c));
 sg13g2_inv_1 clkload206 (.A(clknet_leaf_156_clk_p2c));
 sg13g2_inv_1 clkload207 (.A(clknet_leaf_144_clk_p2c));
 sg13g2_inv_1 clkload208 (.A(clknet_leaf_145_clk_p2c));
 sg13g2_buf_8 clkload209 (.A(clknet_leaf_146_clk_p2c));
 sg13g2_inv_1 clkload210 (.A(clknet_leaf_147_clk_p2c));
 sg13g2_inv_1 clkload211 (.A(clknet_leaf_148_clk_p2c));
 sg13g2_inv_2 clkload212 (.A(clknet_leaf_149_clk_p2c));
 sg13g2_inv_1 clkload213 (.A(clknet_leaf_154_clk_p2c));
 sg13g2_inv_2 clkload214 (.A(clknet_leaf_155_clk_p2c));
 sg13g2_inv_2 clkload215 (.A(clknet_leaf_132_clk_p2c));
 sg13g2_inv_2 clkload216 (.A(clknet_leaf_134_clk_p2c));
 sg13g2_inv_1 clkload217 (.A(clknet_leaf_135_clk_p2c));
 sg13g2_inv_2 clkload218 (.A(clknet_leaf_143_clk_p2c));
 sg13g2_inv_1 clkload219 (.A(clknet_leaf_137_clk_p2c));
 sg13g2_inv_1 clkload220 (.A(clknet_leaf_138_clk_p2c));
 sg13g2_inv_1 clkload221 (.A(clknet_leaf_139_clk_p2c));
 sg13g2_inv_2 clkload222 (.A(clknet_leaf_140_clk_p2c));
 sg13g2_inv_2 clkload223 (.A(clknet_leaf_141_clk_p2c));
 sg13g2_buf_8 clkload224 (.A(clknet_leaf_142_clk_p2c));
 sg13g2_antennanp ANTENNA_1 (.A(net356));
 sg13g2_antennanp ANTENNA_2 (.A(net356));
 sg13g2_antennanp ANTENNA_3 (.A(net356));
 sg13g2_antennanp ANTENNA_4 (.A(net356));
 sg13g2_antennanp ANTENNA_5 (.A(net356));
 sg13g2_antennanp ANTENNA_6 (.A(clk_p2c));
 sg13g2_antennanp ANTENNA_7 (.A(clk_p2c));
 sg13g2_antennanp ANTENNA_8 (.A(data_in_p2c_1));
 sg13g2_antennanp ANTENNA_9 (.A(data_in_p2c_1));
 sg13g2_antennanp ANTENNA_10 (.A(data_in_p2c_1));
 sg13g2_antennanp ANTENNA_11 (.A(data_in_p2c_1));
 sg13g2_antennanp ANTENNA_12 (.A(data_in_p2c_1));
 sg13g2_antennanp ANTENNA_13 (.A(data_in_p2c_1));
 sg13g2_antennanp ANTENNA_14 (.A(data_in_p2c_1));
 sg13g2_antennanp ANTENNA_15 (.A(data_in_p2c_1));
 sg13g2_antennanp ANTENNA_16 (.A(data_in_p2c_1));
 sg13g2_antennanp ANTENNA_17 (.A(data_in_p2c_1));
 sg13g2_antennanp ANTENNA_18 (.A(data_in_p2c_2));
 sg13g2_antennanp ANTENNA_19 (.A(data_in_p2c_2));
 sg13g2_antennanp ANTENNA_20 (.A(data_in_p2c_2));
 sg13g2_antennanp ANTENNA_21 (.A(data_in_p2c_3));
 sg13g2_antennanp ANTENNA_22 (.A(data_in_p2c_3));
 sg13g2_antennanp ANTENNA_23 (.A(data_in_p2c_3));
 sg13g2_antennanp ANTENNA_24 (.A(data_in_p2c_3));
 sg13g2_antennanp ANTENNA_25 (.A(data_in_p2c_3));
 sg13g2_antennanp ANTENNA_26 (.A(data_in_p2c_3));
 sg13g2_antennanp ANTENNA_27 (.A(data_in_p2c_3));
 sg13g2_antennanp ANTENNA_28 (.A(data_in_p2c_3));
 sg13g2_antennanp ANTENNA_29 (.A(net356));
 sg13g2_antennanp ANTENNA_30 (.A(net356));
 sg13g2_antennanp ANTENNA_31 (.A(net356));
 sg13g2_antennanp ANTENNA_32 (.A(net356));
 sg13g2_antennanp ANTENNA_33 (.A(net356));
 sg13g2_antennanp ANTENNA_34 (.A(clk_p2c));
 sg13g2_antennanp ANTENNA_35 (.A(clk_p2c));
 sg13g2_antennanp ANTENNA_36 (.A(data_in_p2c_1));
 sg13g2_antennanp ANTENNA_37 (.A(data_in_p2c_1));
 sg13g2_antennanp ANTENNA_38 (.A(data_in_p2c_1));
 sg13g2_antennanp ANTENNA_39 (.A(data_in_p2c_1));
 sg13g2_antennanp ANTENNA_40 (.A(data_in_p2c_1));
 sg13g2_antennanp ANTENNA_41 (.A(data_in_p2c_1));
 sg13g2_antennanp ANTENNA_42 (.A(data_in_p2c_1));
 sg13g2_antennanp ANTENNA_43 (.A(data_in_p2c_1));
 sg13g2_antennanp ANTENNA_44 (.A(data_in_p2c_1));
 sg13g2_antennanp ANTENNA_45 (.A(data_in_p2c_1));
 sg13g2_antennanp ANTENNA_46 (.A(data_in_p2c_2));
 sg13g2_antennanp ANTENNA_47 (.A(data_in_p2c_2));
 sg13g2_antennanp ANTENNA_48 (.A(data_in_p2c_2));
 sg13g2_antennanp ANTENNA_49 (.A(data_in_p2c_3));
 sg13g2_antennanp ANTENNA_50 (.A(data_in_p2c_3));
 sg13g2_antennanp ANTENNA_51 (.A(data_in_p2c_3));
 sg13g2_antennanp ANTENNA_52 (.A(data_in_p2c_3));
 sg13g2_antennanp ANTENNA_53 (.A(data_in_p2c_3));
 sg13g2_antennanp ANTENNA_54 (.A(data_in_p2c_3));
 sg13g2_antennanp ANTENNA_55 (.A(data_in_p2c_3));
 sg13g2_antennanp ANTENNA_56 (.A(data_in_p2c_3));
 sg13g2_antennanp ANTENNA_57 (.A(data_in_p2c_3));
 sg13g2_antennanp ANTENNA_58 (.A(data_in_p2c_3));
 sg13g2_antennanp ANTENNA_59 (.A(data_in_p2c_3));
 sg13g2_antennanp ANTENNA_60 (.A(data_in_p2c_3));
 sg13g2_antennanp ANTENNA_61 (.A(data_in_p2c_3));
 sg13g2_antennanp ANTENNA_62 (.A(data_in_p2c_3));
 sg13g2_antennanp ANTENNA_63 (.A(data_in_p2c_3));
 sg13g2_antennanp ANTENNA_64 (.A(data_in_p2c_3));
 sg13g2_antennanp ANTENNA_65 (.A(data_in_p2c_3));
 sg13g2_antennanp ANTENNA_66 (.A(data_in_p2c_3));
 sg13g2_antennanp ANTENNA_67 (.A(data_in_p2c_3));
 sg13g2_antennanp ANTENNA_68 (.A(data_in_p2c_3));
 sg13g2_antennanp ANTENNA_69 (.A(net356));
 sg13g2_antennanp ANTENNA_70 (.A(net356));
 sg13g2_antennanp ANTENNA_71 (.A(net356));
 sg13g2_antennanp ANTENNA_72 (.A(net356));
 sg13g2_antennanp ANTENNA_73 (.A(net356));
 sg13g2_antennanp ANTENNA_74 (.A(clk_p2c));
 sg13g2_antennanp ANTENNA_75 (.A(clk_p2c));
 sg13g2_antennanp ANTENNA_76 (.A(data_in_p2c_1));
 sg13g2_antennanp ANTENNA_77 (.A(data_in_p2c_1));
 sg13g2_antennanp ANTENNA_78 (.A(data_in_p2c_1));
 sg13g2_antennanp ANTENNA_79 (.A(data_in_p2c_1));
 sg13g2_antennanp ANTENNA_80 (.A(data_in_p2c_1));
 sg13g2_antennanp ANTENNA_81 (.A(data_in_p2c_1));
 sg13g2_antennanp ANTENNA_82 (.A(data_in_p2c_1));
 sg13g2_antennanp ANTENNA_83 (.A(data_in_p2c_1));
 sg13g2_antennanp ANTENNA_84 (.A(data_in_p2c_1));
 sg13g2_antennanp ANTENNA_85 (.A(data_in_p2c_1));
 sg13g2_antennanp ANTENNA_86 (.A(data_in_p2c_2));
 sg13g2_antennanp ANTENNA_87 (.A(data_in_p2c_2));
 sg13g2_antennanp ANTENNA_88 (.A(data_in_p2c_2));
 sg13g2_antennanp ANTENNA_89 (.A(net356));
 sg13g2_antennanp ANTENNA_90 (.A(net356));
 sg13g2_antennanp ANTENNA_91 (.A(net356));
 sg13g2_antennanp ANTENNA_92 (.A(net356));
 sg13g2_antennanp ANTENNA_93 (.A(net356));
 sg13g2_antennanp ANTENNA_94 (.A(clk_p2c));
 sg13g2_antennanp ANTENNA_95 (.A(clk_p2c));
 sg13g2_antennanp ANTENNA_96 (.A(data_in_p2c_2));
 sg13g2_antennanp ANTENNA_97 (.A(data_in_p2c_2));
 sg13g2_antennanp ANTENNA_98 (.A(data_in_p2c_2));
 sg13g2_antennanp ANTENNA_99 (.A(clk_p2c));
 sg13g2_antennanp ANTENNA_100 (.A(clk_p2c));
 sg13g2_antennanp ANTENNA_101 (.A(data_in_p2c_2));
 sg13g2_antennanp ANTENNA_102 (.A(data_in_p2c_2));
 sg13g2_antennanp ANTENNA_103 (.A(data_in_p2c_2));
 sg13g2_decap_8 FILLER_0_0_0 ();
 sg13g2_decap_8 FILLER_0_0_7 ();
 sg13g2_decap_8 FILLER_0_0_14 ();
 sg13g2_decap_8 FILLER_0_0_21 ();
 sg13g2_decap_8 FILLER_0_0_28 ();
 sg13g2_decap_8 FILLER_0_0_35 ();
 sg13g2_decap_8 FILLER_0_0_42 ();
 sg13g2_decap_8 FILLER_0_0_49 ();
 sg13g2_decap_8 FILLER_0_0_56 ();
 sg13g2_decap_8 FILLER_0_0_63 ();
 sg13g2_decap_8 FILLER_0_0_70 ();
 sg13g2_decap_8 FILLER_0_0_77 ();
 sg13g2_decap_8 FILLER_0_0_84 ();
 sg13g2_decap_8 FILLER_0_0_91 ();
 sg13g2_decap_8 FILLER_0_0_98 ();
 sg13g2_decap_8 FILLER_0_0_105 ();
 sg13g2_decap_8 FILLER_0_0_112 ();
 sg13g2_decap_8 FILLER_0_0_119 ();
 sg13g2_decap_8 FILLER_0_0_126 ();
 sg13g2_decap_8 FILLER_0_0_133 ();
 sg13g2_decap_8 FILLER_0_0_140 ();
 sg13g2_decap_8 FILLER_0_0_147 ();
 sg13g2_decap_8 FILLER_0_0_154 ();
 sg13g2_decap_8 FILLER_0_0_161 ();
 sg13g2_decap_8 FILLER_0_0_168 ();
 sg13g2_decap_8 FILLER_0_0_175 ();
 sg13g2_decap_8 FILLER_0_0_182 ();
 sg13g2_decap_8 FILLER_0_0_189 ();
 sg13g2_decap_8 FILLER_0_0_196 ();
 sg13g2_decap_8 FILLER_0_0_203 ();
 sg13g2_decap_8 FILLER_0_0_210 ();
 sg13g2_decap_8 FILLER_0_0_217 ();
 sg13g2_decap_8 FILLER_0_0_224 ();
 sg13g2_decap_8 FILLER_0_0_231 ();
 sg13g2_decap_8 FILLER_0_0_238 ();
 sg13g2_decap_8 FILLER_0_0_245 ();
 sg13g2_decap_8 FILLER_0_0_252 ();
 sg13g2_decap_8 FILLER_0_0_259 ();
 sg13g2_decap_8 FILLER_0_0_266 ();
 sg13g2_decap_8 FILLER_0_0_273 ();
 sg13g2_decap_8 FILLER_0_0_280 ();
 sg13g2_decap_8 FILLER_0_0_287 ();
 sg13g2_decap_8 FILLER_0_0_294 ();
 sg13g2_decap_8 FILLER_0_0_301 ();
 sg13g2_decap_8 FILLER_0_0_308 ();
 sg13g2_decap_8 FILLER_0_0_315 ();
 sg13g2_decap_8 FILLER_0_0_322 ();
 sg13g2_decap_8 FILLER_0_0_329 ();
 sg13g2_decap_8 FILLER_0_0_336 ();
 sg13g2_decap_8 FILLER_0_0_343 ();
 sg13g2_decap_8 FILLER_0_0_350 ();
 sg13g2_decap_8 FILLER_0_0_357 ();
 sg13g2_decap_8 FILLER_0_0_364 ();
 sg13g2_decap_8 FILLER_0_0_371 ();
 sg13g2_decap_8 FILLER_0_0_378 ();
 sg13g2_decap_8 FILLER_0_0_385 ();
 sg13g2_decap_8 FILLER_0_0_392 ();
 sg13g2_decap_8 FILLER_0_0_399 ();
 sg13g2_decap_8 FILLER_0_0_406 ();
 sg13g2_decap_8 FILLER_0_0_413 ();
 sg13g2_decap_8 FILLER_0_0_420 ();
 sg13g2_decap_8 FILLER_0_0_427 ();
 sg13g2_decap_8 FILLER_0_0_434 ();
 sg13g2_decap_8 FILLER_0_0_441 ();
 sg13g2_decap_8 FILLER_0_0_448 ();
 sg13g2_decap_8 FILLER_0_0_455 ();
 sg13g2_decap_8 FILLER_0_0_462 ();
 sg13g2_decap_8 FILLER_0_0_469 ();
 sg13g2_decap_8 FILLER_0_0_476 ();
 sg13g2_decap_8 FILLER_0_0_483 ();
 sg13g2_decap_8 FILLER_0_0_490 ();
 sg13g2_decap_8 FILLER_0_0_497 ();
 sg13g2_decap_8 FILLER_0_0_504 ();
 sg13g2_decap_8 FILLER_0_0_511 ();
 sg13g2_decap_8 FILLER_0_0_518 ();
 sg13g2_decap_8 FILLER_0_0_525 ();
 sg13g2_decap_8 FILLER_0_0_532 ();
 sg13g2_decap_8 FILLER_0_0_539 ();
 sg13g2_decap_8 FILLER_0_0_546 ();
 sg13g2_decap_8 FILLER_0_0_553 ();
 sg13g2_decap_8 FILLER_0_0_560 ();
 sg13g2_decap_8 FILLER_0_0_567 ();
 sg13g2_decap_8 FILLER_0_0_574 ();
 sg13g2_decap_8 FILLER_0_0_581 ();
 sg13g2_decap_8 FILLER_0_0_588 ();
 sg13g2_decap_8 FILLER_0_0_595 ();
 sg13g2_decap_8 FILLER_0_0_602 ();
 sg13g2_decap_8 FILLER_0_0_609 ();
 sg13g2_decap_8 FILLER_0_0_616 ();
 sg13g2_decap_8 FILLER_0_0_623 ();
 sg13g2_decap_8 FILLER_0_0_630 ();
 sg13g2_decap_8 FILLER_0_0_637 ();
 sg13g2_decap_8 FILLER_0_0_644 ();
 sg13g2_decap_8 FILLER_0_0_651 ();
 sg13g2_decap_8 FILLER_0_0_658 ();
 sg13g2_decap_8 FILLER_0_0_665 ();
 sg13g2_decap_8 FILLER_0_0_672 ();
 sg13g2_decap_8 FILLER_0_0_679 ();
 sg13g2_decap_8 FILLER_0_0_686 ();
 sg13g2_decap_8 FILLER_0_0_693 ();
 sg13g2_decap_8 FILLER_0_0_700 ();
 sg13g2_decap_8 FILLER_0_0_707 ();
 sg13g2_decap_8 FILLER_0_0_714 ();
 sg13g2_decap_8 FILLER_0_0_721 ();
 sg13g2_decap_8 FILLER_0_0_728 ();
 sg13g2_decap_8 FILLER_0_0_735 ();
 sg13g2_decap_8 FILLER_0_0_742 ();
 sg13g2_decap_8 FILLER_0_0_749 ();
 sg13g2_decap_8 FILLER_0_0_756 ();
 sg13g2_decap_8 FILLER_0_0_763 ();
 sg13g2_decap_8 FILLER_0_0_770 ();
 sg13g2_decap_8 FILLER_0_0_777 ();
 sg13g2_decap_8 FILLER_0_0_784 ();
 sg13g2_decap_8 FILLER_0_0_791 ();
 sg13g2_decap_8 FILLER_0_0_798 ();
 sg13g2_decap_8 FILLER_0_0_805 ();
 sg13g2_decap_8 FILLER_0_0_812 ();
 sg13g2_decap_8 FILLER_0_0_819 ();
 sg13g2_decap_8 FILLER_0_0_826 ();
 sg13g2_decap_8 FILLER_0_0_833 ();
 sg13g2_decap_8 FILLER_0_0_840 ();
 sg13g2_decap_8 FILLER_0_0_847 ();
 sg13g2_decap_8 FILLER_0_0_854 ();
 sg13g2_decap_8 FILLER_0_0_861 ();
 sg13g2_decap_8 FILLER_0_0_868 ();
 sg13g2_decap_8 FILLER_0_0_875 ();
 sg13g2_decap_8 FILLER_0_0_882 ();
 sg13g2_decap_8 FILLER_0_0_889 ();
 sg13g2_decap_8 FILLER_0_0_896 ();
 sg13g2_decap_8 FILLER_0_0_903 ();
 sg13g2_decap_8 FILLER_0_0_910 ();
 sg13g2_decap_8 FILLER_0_0_917 ();
 sg13g2_decap_8 FILLER_0_0_924 ();
 sg13g2_decap_8 FILLER_0_0_931 ();
 sg13g2_decap_8 FILLER_0_0_938 ();
 sg13g2_decap_8 FILLER_0_0_945 ();
 sg13g2_decap_8 FILLER_0_0_952 ();
 sg13g2_decap_8 FILLER_0_0_959 ();
 sg13g2_decap_8 FILLER_0_0_966 ();
 sg13g2_decap_8 FILLER_0_0_973 ();
 sg13g2_decap_8 FILLER_0_0_980 ();
 sg13g2_decap_8 FILLER_0_0_987 ();
 sg13g2_decap_8 FILLER_0_0_994 ();
 sg13g2_decap_8 FILLER_0_0_1001 ();
 sg13g2_decap_8 FILLER_0_0_1008 ();
 sg13g2_decap_8 FILLER_0_0_1015 ();
 sg13g2_decap_8 FILLER_0_0_1022 ();
 sg13g2_decap_8 FILLER_0_0_1029 ();
 sg13g2_decap_8 FILLER_0_0_1036 ();
 sg13g2_decap_8 FILLER_0_0_1043 ();
 sg13g2_decap_8 FILLER_0_0_1050 ();
 sg13g2_decap_8 FILLER_0_0_1057 ();
 sg13g2_decap_8 FILLER_0_0_1064 ();
 sg13g2_decap_8 FILLER_0_0_1071 ();
 sg13g2_decap_8 FILLER_0_0_1078 ();
 sg13g2_decap_8 FILLER_0_0_1085 ();
 sg13g2_decap_8 FILLER_0_0_1092 ();
 sg13g2_decap_8 FILLER_0_0_1099 ();
 sg13g2_decap_8 FILLER_0_0_1106 ();
 sg13g2_decap_8 FILLER_0_0_1113 ();
 sg13g2_decap_8 FILLER_0_0_1120 ();
 sg13g2_decap_8 FILLER_0_0_1127 ();
 sg13g2_decap_8 FILLER_0_0_1134 ();
 sg13g2_decap_8 FILLER_0_0_1141 ();
 sg13g2_decap_8 FILLER_0_0_1148 ();
 sg13g2_decap_8 FILLER_0_0_1155 ();
 sg13g2_decap_8 FILLER_0_0_1162 ();
 sg13g2_decap_8 FILLER_0_0_1169 ();
 sg13g2_decap_8 FILLER_0_0_1176 ();
 sg13g2_decap_8 FILLER_0_0_1183 ();
 sg13g2_decap_8 FILLER_0_0_1190 ();
 sg13g2_decap_8 FILLER_0_0_1197 ();
 sg13g2_decap_8 FILLER_0_0_1204 ();
 sg13g2_decap_8 FILLER_0_0_1211 ();
 sg13g2_decap_8 FILLER_0_0_1218 ();
 sg13g2_fill_2 FILLER_0_0_1225 ();
 sg13g2_fill_1 FILLER_0_0_1227 ();
 sg13g2_decap_8 FILLER_0_1_0 ();
 sg13g2_decap_8 FILLER_0_1_7 ();
 sg13g2_decap_8 FILLER_0_1_14 ();
 sg13g2_decap_8 FILLER_0_1_21 ();
 sg13g2_decap_8 FILLER_0_1_28 ();
 sg13g2_decap_8 FILLER_0_1_35 ();
 sg13g2_decap_8 FILLER_0_1_42 ();
 sg13g2_decap_8 FILLER_0_1_49 ();
 sg13g2_decap_8 FILLER_0_1_56 ();
 sg13g2_decap_8 FILLER_0_1_63 ();
 sg13g2_decap_8 FILLER_0_1_70 ();
 sg13g2_decap_8 FILLER_0_1_77 ();
 sg13g2_decap_8 FILLER_0_1_84 ();
 sg13g2_decap_8 FILLER_0_1_91 ();
 sg13g2_decap_8 FILLER_0_1_98 ();
 sg13g2_decap_8 FILLER_0_1_105 ();
 sg13g2_decap_8 FILLER_0_1_112 ();
 sg13g2_decap_8 FILLER_0_1_119 ();
 sg13g2_decap_8 FILLER_0_1_126 ();
 sg13g2_decap_8 FILLER_0_1_133 ();
 sg13g2_decap_8 FILLER_0_1_140 ();
 sg13g2_decap_8 FILLER_0_1_147 ();
 sg13g2_decap_8 FILLER_0_1_154 ();
 sg13g2_decap_8 FILLER_0_1_161 ();
 sg13g2_decap_8 FILLER_0_1_168 ();
 sg13g2_decap_8 FILLER_0_1_175 ();
 sg13g2_decap_8 FILLER_0_1_182 ();
 sg13g2_decap_8 FILLER_0_1_189 ();
 sg13g2_decap_8 FILLER_0_1_196 ();
 sg13g2_decap_8 FILLER_0_1_203 ();
 sg13g2_decap_8 FILLER_0_1_210 ();
 sg13g2_decap_8 FILLER_0_1_217 ();
 sg13g2_decap_8 FILLER_0_1_224 ();
 sg13g2_decap_8 FILLER_0_1_231 ();
 sg13g2_decap_8 FILLER_0_1_238 ();
 sg13g2_decap_8 FILLER_0_1_245 ();
 sg13g2_decap_8 FILLER_0_1_252 ();
 sg13g2_decap_8 FILLER_0_1_259 ();
 sg13g2_decap_8 FILLER_0_1_266 ();
 sg13g2_decap_8 FILLER_0_1_273 ();
 sg13g2_decap_8 FILLER_0_1_280 ();
 sg13g2_decap_8 FILLER_0_1_287 ();
 sg13g2_decap_8 FILLER_0_1_294 ();
 sg13g2_decap_8 FILLER_0_1_301 ();
 sg13g2_decap_8 FILLER_0_1_308 ();
 sg13g2_decap_8 FILLER_0_1_315 ();
 sg13g2_decap_8 FILLER_0_1_322 ();
 sg13g2_decap_8 FILLER_0_1_329 ();
 sg13g2_decap_8 FILLER_0_1_336 ();
 sg13g2_decap_8 FILLER_0_1_343 ();
 sg13g2_decap_8 FILLER_0_1_350 ();
 sg13g2_decap_8 FILLER_0_1_357 ();
 sg13g2_decap_8 FILLER_0_1_364 ();
 sg13g2_decap_8 FILLER_0_1_371 ();
 sg13g2_decap_8 FILLER_0_1_378 ();
 sg13g2_decap_8 FILLER_0_1_385 ();
 sg13g2_decap_8 FILLER_0_1_392 ();
 sg13g2_decap_8 FILLER_0_1_399 ();
 sg13g2_decap_8 FILLER_0_1_406 ();
 sg13g2_decap_8 FILLER_0_1_413 ();
 sg13g2_decap_8 FILLER_0_1_420 ();
 sg13g2_decap_8 FILLER_0_1_427 ();
 sg13g2_decap_8 FILLER_0_1_434 ();
 sg13g2_decap_8 FILLER_0_1_441 ();
 sg13g2_decap_8 FILLER_0_1_448 ();
 sg13g2_decap_8 FILLER_0_1_455 ();
 sg13g2_decap_8 FILLER_0_1_462 ();
 sg13g2_decap_8 FILLER_0_1_469 ();
 sg13g2_decap_8 FILLER_0_1_476 ();
 sg13g2_decap_8 FILLER_0_1_483 ();
 sg13g2_decap_8 FILLER_0_1_490 ();
 sg13g2_decap_8 FILLER_0_1_497 ();
 sg13g2_decap_8 FILLER_0_1_504 ();
 sg13g2_decap_8 FILLER_0_1_511 ();
 sg13g2_decap_8 FILLER_0_1_518 ();
 sg13g2_decap_8 FILLER_0_1_525 ();
 sg13g2_decap_8 FILLER_0_1_532 ();
 sg13g2_decap_8 FILLER_0_1_539 ();
 sg13g2_decap_8 FILLER_0_1_546 ();
 sg13g2_decap_8 FILLER_0_1_553 ();
 sg13g2_decap_8 FILLER_0_1_560 ();
 sg13g2_decap_8 FILLER_0_1_567 ();
 sg13g2_decap_8 FILLER_0_1_574 ();
 sg13g2_decap_8 FILLER_0_1_581 ();
 sg13g2_decap_8 FILLER_0_1_588 ();
 sg13g2_decap_8 FILLER_0_1_595 ();
 sg13g2_decap_8 FILLER_0_1_602 ();
 sg13g2_decap_8 FILLER_0_1_609 ();
 sg13g2_decap_8 FILLER_0_1_616 ();
 sg13g2_decap_8 FILLER_0_1_623 ();
 sg13g2_decap_8 FILLER_0_1_630 ();
 sg13g2_decap_8 FILLER_0_1_637 ();
 sg13g2_decap_8 FILLER_0_1_644 ();
 sg13g2_decap_8 FILLER_0_1_651 ();
 sg13g2_decap_8 FILLER_0_1_658 ();
 sg13g2_decap_8 FILLER_0_1_665 ();
 sg13g2_decap_8 FILLER_0_1_672 ();
 sg13g2_decap_8 FILLER_0_1_679 ();
 sg13g2_decap_8 FILLER_0_1_686 ();
 sg13g2_decap_8 FILLER_0_1_693 ();
 sg13g2_decap_8 FILLER_0_1_700 ();
 sg13g2_decap_8 FILLER_0_1_707 ();
 sg13g2_decap_8 FILLER_0_1_714 ();
 sg13g2_decap_8 FILLER_0_1_721 ();
 sg13g2_decap_8 FILLER_0_1_728 ();
 sg13g2_decap_8 FILLER_0_1_735 ();
 sg13g2_decap_8 FILLER_0_1_742 ();
 sg13g2_decap_8 FILLER_0_1_749 ();
 sg13g2_decap_8 FILLER_0_1_756 ();
 sg13g2_decap_8 FILLER_0_1_763 ();
 sg13g2_decap_8 FILLER_0_1_770 ();
 sg13g2_decap_8 FILLER_0_1_777 ();
 sg13g2_decap_8 FILLER_0_1_784 ();
 sg13g2_decap_8 FILLER_0_1_791 ();
 sg13g2_decap_8 FILLER_0_1_798 ();
 sg13g2_decap_8 FILLER_0_1_805 ();
 sg13g2_decap_8 FILLER_0_1_812 ();
 sg13g2_decap_8 FILLER_0_1_819 ();
 sg13g2_decap_8 FILLER_0_1_826 ();
 sg13g2_decap_8 FILLER_0_1_833 ();
 sg13g2_decap_8 FILLER_0_1_840 ();
 sg13g2_decap_8 FILLER_0_1_847 ();
 sg13g2_decap_8 FILLER_0_1_854 ();
 sg13g2_decap_8 FILLER_0_1_861 ();
 sg13g2_decap_8 FILLER_0_1_868 ();
 sg13g2_decap_8 FILLER_0_1_875 ();
 sg13g2_decap_8 FILLER_0_1_882 ();
 sg13g2_decap_8 FILLER_0_1_889 ();
 sg13g2_decap_8 FILLER_0_1_896 ();
 sg13g2_decap_8 FILLER_0_1_903 ();
 sg13g2_decap_8 FILLER_0_1_910 ();
 sg13g2_decap_8 FILLER_0_1_917 ();
 sg13g2_decap_8 FILLER_0_1_924 ();
 sg13g2_decap_8 FILLER_0_1_931 ();
 sg13g2_decap_8 FILLER_0_1_938 ();
 sg13g2_decap_8 FILLER_0_1_945 ();
 sg13g2_decap_8 FILLER_0_1_952 ();
 sg13g2_decap_8 FILLER_0_1_959 ();
 sg13g2_decap_8 FILLER_0_1_966 ();
 sg13g2_decap_8 FILLER_0_1_973 ();
 sg13g2_decap_8 FILLER_0_1_980 ();
 sg13g2_decap_8 FILLER_0_1_987 ();
 sg13g2_decap_8 FILLER_0_1_994 ();
 sg13g2_decap_8 FILLER_0_1_1001 ();
 sg13g2_decap_8 FILLER_0_1_1008 ();
 sg13g2_decap_8 FILLER_0_1_1015 ();
 sg13g2_decap_8 FILLER_0_1_1022 ();
 sg13g2_decap_8 FILLER_0_1_1029 ();
 sg13g2_decap_8 FILLER_0_1_1036 ();
 sg13g2_decap_8 FILLER_0_1_1043 ();
 sg13g2_decap_8 FILLER_0_1_1050 ();
 sg13g2_decap_8 FILLER_0_1_1057 ();
 sg13g2_decap_8 FILLER_0_1_1064 ();
 sg13g2_decap_8 FILLER_0_1_1071 ();
 sg13g2_decap_8 FILLER_0_1_1078 ();
 sg13g2_decap_8 FILLER_0_1_1085 ();
 sg13g2_decap_8 FILLER_0_1_1092 ();
 sg13g2_decap_8 FILLER_0_1_1099 ();
 sg13g2_decap_8 FILLER_0_1_1106 ();
 sg13g2_decap_8 FILLER_0_1_1113 ();
 sg13g2_decap_8 FILLER_0_1_1120 ();
 sg13g2_decap_8 FILLER_0_1_1127 ();
 sg13g2_decap_8 FILLER_0_1_1134 ();
 sg13g2_decap_8 FILLER_0_1_1141 ();
 sg13g2_decap_8 FILLER_0_1_1148 ();
 sg13g2_decap_8 FILLER_0_1_1155 ();
 sg13g2_decap_8 FILLER_0_1_1162 ();
 sg13g2_decap_8 FILLER_0_1_1169 ();
 sg13g2_decap_8 FILLER_0_1_1176 ();
 sg13g2_decap_8 FILLER_0_1_1183 ();
 sg13g2_decap_8 FILLER_0_1_1190 ();
 sg13g2_decap_8 FILLER_0_1_1197 ();
 sg13g2_decap_8 FILLER_0_1_1204 ();
 sg13g2_decap_8 FILLER_0_1_1211 ();
 sg13g2_decap_8 FILLER_0_1_1218 ();
 sg13g2_fill_2 FILLER_0_1_1225 ();
 sg13g2_fill_1 FILLER_0_1_1227 ();
 sg13g2_decap_8 FILLER_0_2_0 ();
 sg13g2_decap_8 FILLER_0_2_7 ();
 sg13g2_decap_8 FILLER_0_2_14 ();
 sg13g2_decap_8 FILLER_0_2_21 ();
 sg13g2_decap_8 FILLER_0_2_28 ();
 sg13g2_decap_8 FILLER_0_2_35 ();
 sg13g2_decap_8 FILLER_0_2_42 ();
 sg13g2_decap_8 FILLER_0_2_49 ();
 sg13g2_decap_8 FILLER_0_2_56 ();
 sg13g2_decap_8 FILLER_0_2_63 ();
 sg13g2_decap_8 FILLER_0_2_70 ();
 sg13g2_decap_8 FILLER_0_2_77 ();
 sg13g2_decap_8 FILLER_0_2_84 ();
 sg13g2_decap_8 FILLER_0_2_91 ();
 sg13g2_decap_8 FILLER_0_2_98 ();
 sg13g2_decap_8 FILLER_0_2_105 ();
 sg13g2_decap_8 FILLER_0_2_112 ();
 sg13g2_decap_8 FILLER_0_2_119 ();
 sg13g2_decap_8 FILLER_0_2_126 ();
 sg13g2_decap_8 FILLER_0_2_133 ();
 sg13g2_decap_8 FILLER_0_2_140 ();
 sg13g2_decap_8 FILLER_0_2_147 ();
 sg13g2_decap_8 FILLER_0_2_154 ();
 sg13g2_decap_8 FILLER_0_2_161 ();
 sg13g2_decap_8 FILLER_0_2_168 ();
 sg13g2_decap_8 FILLER_0_2_175 ();
 sg13g2_decap_8 FILLER_0_2_182 ();
 sg13g2_decap_8 FILLER_0_2_189 ();
 sg13g2_decap_8 FILLER_0_2_196 ();
 sg13g2_decap_8 FILLER_0_2_203 ();
 sg13g2_decap_8 FILLER_0_2_210 ();
 sg13g2_decap_8 FILLER_0_2_217 ();
 sg13g2_decap_8 FILLER_0_2_224 ();
 sg13g2_decap_8 FILLER_0_2_231 ();
 sg13g2_decap_8 FILLER_0_2_238 ();
 sg13g2_decap_8 FILLER_0_2_245 ();
 sg13g2_decap_8 FILLER_0_2_252 ();
 sg13g2_decap_8 FILLER_0_2_259 ();
 sg13g2_decap_8 FILLER_0_2_266 ();
 sg13g2_decap_8 FILLER_0_2_273 ();
 sg13g2_decap_8 FILLER_0_2_280 ();
 sg13g2_decap_8 FILLER_0_2_287 ();
 sg13g2_decap_8 FILLER_0_2_294 ();
 sg13g2_decap_8 FILLER_0_2_301 ();
 sg13g2_decap_8 FILLER_0_2_308 ();
 sg13g2_decap_8 FILLER_0_2_315 ();
 sg13g2_decap_8 FILLER_0_2_322 ();
 sg13g2_decap_8 FILLER_0_2_329 ();
 sg13g2_decap_8 FILLER_0_2_336 ();
 sg13g2_decap_8 FILLER_0_2_343 ();
 sg13g2_decap_8 FILLER_0_2_350 ();
 sg13g2_decap_8 FILLER_0_2_357 ();
 sg13g2_decap_8 FILLER_0_2_364 ();
 sg13g2_decap_8 FILLER_0_2_371 ();
 sg13g2_decap_8 FILLER_0_2_378 ();
 sg13g2_decap_8 FILLER_0_2_385 ();
 sg13g2_decap_8 FILLER_0_2_392 ();
 sg13g2_decap_8 FILLER_0_2_399 ();
 sg13g2_decap_8 FILLER_0_2_406 ();
 sg13g2_decap_8 FILLER_0_2_413 ();
 sg13g2_decap_8 FILLER_0_2_420 ();
 sg13g2_decap_8 FILLER_0_2_427 ();
 sg13g2_decap_8 FILLER_0_2_434 ();
 sg13g2_decap_8 FILLER_0_2_441 ();
 sg13g2_decap_8 FILLER_0_2_448 ();
 sg13g2_decap_8 FILLER_0_2_455 ();
 sg13g2_decap_8 FILLER_0_2_462 ();
 sg13g2_decap_8 FILLER_0_2_469 ();
 sg13g2_decap_8 FILLER_0_2_476 ();
 sg13g2_decap_8 FILLER_0_2_483 ();
 sg13g2_decap_8 FILLER_0_2_490 ();
 sg13g2_decap_8 FILLER_0_2_497 ();
 sg13g2_decap_8 FILLER_0_2_504 ();
 sg13g2_decap_8 FILLER_0_2_511 ();
 sg13g2_decap_8 FILLER_0_2_518 ();
 sg13g2_decap_8 FILLER_0_2_525 ();
 sg13g2_decap_8 FILLER_0_2_532 ();
 sg13g2_decap_8 FILLER_0_2_539 ();
 sg13g2_decap_8 FILLER_0_2_546 ();
 sg13g2_decap_8 FILLER_0_2_553 ();
 sg13g2_decap_8 FILLER_0_2_560 ();
 sg13g2_decap_8 FILLER_0_2_567 ();
 sg13g2_decap_8 FILLER_0_2_574 ();
 sg13g2_decap_8 FILLER_0_2_581 ();
 sg13g2_decap_8 FILLER_0_2_588 ();
 sg13g2_decap_8 FILLER_0_2_595 ();
 sg13g2_decap_8 FILLER_0_2_602 ();
 sg13g2_decap_8 FILLER_0_2_609 ();
 sg13g2_decap_8 FILLER_0_2_616 ();
 sg13g2_decap_8 FILLER_0_2_623 ();
 sg13g2_decap_8 FILLER_0_2_630 ();
 sg13g2_decap_8 FILLER_0_2_637 ();
 sg13g2_decap_8 FILLER_0_2_644 ();
 sg13g2_decap_8 FILLER_0_2_651 ();
 sg13g2_decap_8 FILLER_0_2_658 ();
 sg13g2_decap_8 FILLER_0_2_665 ();
 sg13g2_decap_8 FILLER_0_2_672 ();
 sg13g2_decap_8 FILLER_0_2_679 ();
 sg13g2_decap_8 FILLER_0_2_686 ();
 sg13g2_decap_8 FILLER_0_2_693 ();
 sg13g2_decap_8 FILLER_0_2_700 ();
 sg13g2_decap_8 FILLER_0_2_707 ();
 sg13g2_decap_8 FILLER_0_2_714 ();
 sg13g2_decap_8 FILLER_0_2_721 ();
 sg13g2_decap_8 FILLER_0_2_728 ();
 sg13g2_decap_8 FILLER_0_2_735 ();
 sg13g2_decap_8 FILLER_0_2_742 ();
 sg13g2_decap_8 FILLER_0_2_749 ();
 sg13g2_decap_8 FILLER_0_2_756 ();
 sg13g2_decap_8 FILLER_0_2_763 ();
 sg13g2_decap_8 FILLER_0_2_770 ();
 sg13g2_decap_8 FILLER_0_2_777 ();
 sg13g2_decap_8 FILLER_0_2_784 ();
 sg13g2_decap_8 FILLER_0_2_791 ();
 sg13g2_decap_8 FILLER_0_2_798 ();
 sg13g2_decap_8 FILLER_0_2_805 ();
 sg13g2_decap_8 FILLER_0_2_812 ();
 sg13g2_decap_8 FILLER_0_2_819 ();
 sg13g2_decap_8 FILLER_0_2_826 ();
 sg13g2_decap_8 FILLER_0_2_833 ();
 sg13g2_decap_8 FILLER_0_2_840 ();
 sg13g2_decap_8 FILLER_0_2_847 ();
 sg13g2_decap_8 FILLER_0_2_854 ();
 sg13g2_decap_8 FILLER_0_2_861 ();
 sg13g2_decap_8 FILLER_0_2_868 ();
 sg13g2_decap_8 FILLER_0_2_875 ();
 sg13g2_decap_8 FILLER_0_2_882 ();
 sg13g2_decap_8 FILLER_0_2_889 ();
 sg13g2_decap_8 FILLER_0_2_896 ();
 sg13g2_decap_8 FILLER_0_2_903 ();
 sg13g2_decap_8 FILLER_0_2_910 ();
 sg13g2_decap_8 FILLER_0_2_917 ();
 sg13g2_decap_8 FILLER_0_2_924 ();
 sg13g2_decap_8 FILLER_0_2_931 ();
 sg13g2_decap_8 FILLER_0_2_938 ();
 sg13g2_decap_8 FILLER_0_2_945 ();
 sg13g2_decap_8 FILLER_0_2_952 ();
 sg13g2_decap_8 FILLER_0_2_959 ();
 sg13g2_decap_8 FILLER_0_2_966 ();
 sg13g2_decap_8 FILLER_0_2_973 ();
 sg13g2_decap_8 FILLER_0_2_980 ();
 sg13g2_decap_8 FILLER_0_2_987 ();
 sg13g2_decap_8 FILLER_0_2_994 ();
 sg13g2_decap_8 FILLER_0_2_1001 ();
 sg13g2_decap_8 FILLER_0_2_1008 ();
 sg13g2_decap_8 FILLER_0_2_1015 ();
 sg13g2_decap_8 FILLER_0_2_1022 ();
 sg13g2_decap_8 FILLER_0_2_1029 ();
 sg13g2_decap_8 FILLER_0_2_1036 ();
 sg13g2_decap_8 FILLER_0_2_1043 ();
 sg13g2_decap_8 FILLER_0_2_1050 ();
 sg13g2_decap_8 FILLER_0_2_1057 ();
 sg13g2_decap_8 FILLER_0_2_1064 ();
 sg13g2_decap_8 FILLER_0_2_1071 ();
 sg13g2_decap_8 FILLER_0_2_1078 ();
 sg13g2_decap_8 FILLER_0_2_1085 ();
 sg13g2_decap_8 FILLER_0_2_1092 ();
 sg13g2_decap_8 FILLER_0_2_1099 ();
 sg13g2_decap_8 FILLER_0_2_1106 ();
 sg13g2_decap_8 FILLER_0_2_1113 ();
 sg13g2_decap_8 FILLER_0_2_1120 ();
 sg13g2_decap_8 FILLER_0_2_1127 ();
 sg13g2_decap_8 FILLER_0_2_1134 ();
 sg13g2_decap_8 FILLER_0_2_1141 ();
 sg13g2_decap_8 FILLER_0_2_1148 ();
 sg13g2_decap_8 FILLER_0_2_1155 ();
 sg13g2_decap_8 FILLER_0_2_1162 ();
 sg13g2_decap_8 FILLER_0_2_1169 ();
 sg13g2_decap_8 FILLER_0_2_1176 ();
 sg13g2_decap_8 FILLER_0_2_1183 ();
 sg13g2_decap_8 FILLER_0_2_1190 ();
 sg13g2_decap_8 FILLER_0_2_1197 ();
 sg13g2_decap_8 FILLER_0_2_1204 ();
 sg13g2_decap_8 FILLER_0_2_1211 ();
 sg13g2_decap_8 FILLER_0_2_1218 ();
 sg13g2_fill_2 FILLER_0_2_1225 ();
 sg13g2_fill_1 FILLER_0_2_1227 ();
 sg13g2_decap_8 FILLER_0_3_0 ();
 sg13g2_decap_8 FILLER_0_3_7 ();
 sg13g2_decap_8 FILLER_0_3_14 ();
 sg13g2_decap_8 FILLER_0_3_21 ();
 sg13g2_decap_8 FILLER_0_3_28 ();
 sg13g2_decap_8 FILLER_0_3_35 ();
 sg13g2_decap_8 FILLER_0_3_42 ();
 sg13g2_decap_8 FILLER_0_3_49 ();
 sg13g2_decap_8 FILLER_0_3_56 ();
 sg13g2_decap_8 FILLER_0_3_63 ();
 sg13g2_decap_8 FILLER_0_3_70 ();
 sg13g2_decap_8 FILLER_0_3_77 ();
 sg13g2_decap_8 FILLER_0_3_84 ();
 sg13g2_decap_8 FILLER_0_3_91 ();
 sg13g2_decap_8 FILLER_0_3_98 ();
 sg13g2_decap_8 FILLER_0_3_105 ();
 sg13g2_decap_8 FILLER_0_3_112 ();
 sg13g2_decap_8 FILLER_0_3_119 ();
 sg13g2_decap_8 FILLER_0_3_126 ();
 sg13g2_decap_8 FILLER_0_3_133 ();
 sg13g2_decap_8 FILLER_0_3_140 ();
 sg13g2_decap_8 FILLER_0_3_147 ();
 sg13g2_decap_8 FILLER_0_3_154 ();
 sg13g2_decap_8 FILLER_0_3_161 ();
 sg13g2_decap_8 FILLER_0_3_168 ();
 sg13g2_decap_8 FILLER_0_3_175 ();
 sg13g2_decap_8 FILLER_0_3_182 ();
 sg13g2_decap_8 FILLER_0_3_189 ();
 sg13g2_decap_8 FILLER_0_3_196 ();
 sg13g2_decap_8 FILLER_0_3_203 ();
 sg13g2_decap_8 FILLER_0_3_210 ();
 sg13g2_decap_8 FILLER_0_3_217 ();
 sg13g2_decap_8 FILLER_0_3_224 ();
 sg13g2_decap_8 FILLER_0_3_231 ();
 sg13g2_decap_8 FILLER_0_3_238 ();
 sg13g2_decap_8 FILLER_0_3_245 ();
 sg13g2_decap_8 FILLER_0_3_252 ();
 sg13g2_decap_8 FILLER_0_3_259 ();
 sg13g2_decap_8 FILLER_0_3_266 ();
 sg13g2_decap_8 FILLER_0_3_273 ();
 sg13g2_decap_8 FILLER_0_3_280 ();
 sg13g2_decap_8 FILLER_0_3_287 ();
 sg13g2_decap_8 FILLER_0_3_294 ();
 sg13g2_decap_8 FILLER_0_3_301 ();
 sg13g2_decap_8 FILLER_0_3_308 ();
 sg13g2_decap_8 FILLER_0_3_315 ();
 sg13g2_decap_8 FILLER_0_3_322 ();
 sg13g2_decap_8 FILLER_0_3_329 ();
 sg13g2_decap_8 FILLER_0_3_336 ();
 sg13g2_decap_8 FILLER_0_3_343 ();
 sg13g2_decap_8 FILLER_0_3_350 ();
 sg13g2_decap_8 FILLER_0_3_357 ();
 sg13g2_decap_8 FILLER_0_3_364 ();
 sg13g2_decap_8 FILLER_0_3_371 ();
 sg13g2_decap_8 FILLER_0_3_378 ();
 sg13g2_decap_8 FILLER_0_3_385 ();
 sg13g2_decap_8 FILLER_0_3_392 ();
 sg13g2_decap_8 FILLER_0_3_399 ();
 sg13g2_decap_8 FILLER_0_3_406 ();
 sg13g2_decap_8 FILLER_0_3_413 ();
 sg13g2_decap_8 FILLER_0_3_420 ();
 sg13g2_decap_8 FILLER_0_3_427 ();
 sg13g2_decap_8 FILLER_0_3_434 ();
 sg13g2_decap_8 FILLER_0_3_441 ();
 sg13g2_decap_8 FILLER_0_3_448 ();
 sg13g2_decap_8 FILLER_0_3_455 ();
 sg13g2_decap_8 FILLER_0_3_462 ();
 sg13g2_decap_8 FILLER_0_3_469 ();
 sg13g2_decap_8 FILLER_0_3_476 ();
 sg13g2_decap_8 FILLER_0_3_483 ();
 sg13g2_decap_8 FILLER_0_3_490 ();
 sg13g2_decap_8 FILLER_0_3_497 ();
 sg13g2_decap_8 FILLER_0_3_504 ();
 sg13g2_decap_8 FILLER_0_3_511 ();
 sg13g2_decap_8 FILLER_0_3_518 ();
 sg13g2_decap_8 FILLER_0_3_525 ();
 sg13g2_decap_8 FILLER_0_3_532 ();
 sg13g2_decap_8 FILLER_0_3_539 ();
 sg13g2_decap_8 FILLER_0_3_546 ();
 sg13g2_decap_8 FILLER_0_3_553 ();
 sg13g2_decap_8 FILLER_0_3_560 ();
 sg13g2_decap_8 FILLER_0_3_567 ();
 sg13g2_decap_8 FILLER_0_3_574 ();
 sg13g2_decap_8 FILLER_0_3_581 ();
 sg13g2_decap_8 FILLER_0_3_588 ();
 sg13g2_decap_8 FILLER_0_3_595 ();
 sg13g2_decap_8 FILLER_0_3_602 ();
 sg13g2_decap_8 FILLER_0_3_609 ();
 sg13g2_decap_8 FILLER_0_3_616 ();
 sg13g2_decap_8 FILLER_0_3_623 ();
 sg13g2_decap_8 FILLER_0_3_630 ();
 sg13g2_decap_8 FILLER_0_3_637 ();
 sg13g2_decap_8 FILLER_0_3_644 ();
 sg13g2_decap_8 FILLER_0_3_651 ();
 sg13g2_decap_8 FILLER_0_3_658 ();
 sg13g2_decap_8 FILLER_0_3_665 ();
 sg13g2_decap_8 FILLER_0_3_672 ();
 sg13g2_decap_8 FILLER_0_3_679 ();
 sg13g2_decap_8 FILLER_0_3_686 ();
 sg13g2_decap_8 FILLER_0_3_693 ();
 sg13g2_decap_8 FILLER_0_3_700 ();
 sg13g2_decap_8 FILLER_0_3_707 ();
 sg13g2_decap_8 FILLER_0_3_714 ();
 sg13g2_decap_8 FILLER_0_3_721 ();
 sg13g2_decap_8 FILLER_0_3_728 ();
 sg13g2_decap_8 FILLER_0_3_735 ();
 sg13g2_decap_8 FILLER_0_3_742 ();
 sg13g2_decap_8 FILLER_0_3_749 ();
 sg13g2_decap_8 FILLER_0_3_756 ();
 sg13g2_decap_8 FILLER_0_3_763 ();
 sg13g2_decap_8 FILLER_0_3_770 ();
 sg13g2_decap_8 FILLER_0_3_777 ();
 sg13g2_decap_8 FILLER_0_3_784 ();
 sg13g2_decap_8 FILLER_0_3_791 ();
 sg13g2_decap_8 FILLER_0_3_798 ();
 sg13g2_decap_8 FILLER_0_3_805 ();
 sg13g2_decap_8 FILLER_0_3_812 ();
 sg13g2_decap_8 FILLER_0_3_819 ();
 sg13g2_decap_8 FILLER_0_3_826 ();
 sg13g2_decap_8 FILLER_0_3_833 ();
 sg13g2_decap_8 FILLER_0_3_840 ();
 sg13g2_decap_8 FILLER_0_3_847 ();
 sg13g2_decap_8 FILLER_0_3_854 ();
 sg13g2_decap_8 FILLER_0_3_861 ();
 sg13g2_decap_8 FILLER_0_3_868 ();
 sg13g2_decap_8 FILLER_0_3_875 ();
 sg13g2_decap_8 FILLER_0_3_882 ();
 sg13g2_decap_8 FILLER_0_3_889 ();
 sg13g2_decap_8 FILLER_0_3_896 ();
 sg13g2_decap_8 FILLER_0_3_903 ();
 sg13g2_decap_8 FILLER_0_3_910 ();
 sg13g2_decap_8 FILLER_0_3_917 ();
 sg13g2_decap_8 FILLER_0_3_924 ();
 sg13g2_decap_8 FILLER_0_3_931 ();
 sg13g2_decap_8 FILLER_0_3_938 ();
 sg13g2_decap_8 FILLER_0_3_945 ();
 sg13g2_decap_8 FILLER_0_3_952 ();
 sg13g2_decap_8 FILLER_0_3_959 ();
 sg13g2_decap_8 FILLER_0_3_966 ();
 sg13g2_decap_8 FILLER_0_3_973 ();
 sg13g2_decap_8 FILLER_0_3_980 ();
 sg13g2_decap_8 FILLER_0_3_987 ();
 sg13g2_decap_8 FILLER_0_3_994 ();
 sg13g2_decap_8 FILLER_0_3_1001 ();
 sg13g2_decap_8 FILLER_0_3_1008 ();
 sg13g2_decap_8 FILLER_0_3_1015 ();
 sg13g2_decap_8 FILLER_0_3_1022 ();
 sg13g2_decap_8 FILLER_0_3_1029 ();
 sg13g2_decap_8 FILLER_0_3_1036 ();
 sg13g2_decap_8 FILLER_0_3_1043 ();
 sg13g2_decap_8 FILLER_0_3_1050 ();
 sg13g2_decap_8 FILLER_0_3_1057 ();
 sg13g2_decap_8 FILLER_0_3_1064 ();
 sg13g2_decap_8 FILLER_0_3_1071 ();
 sg13g2_decap_8 FILLER_0_3_1078 ();
 sg13g2_decap_8 FILLER_0_3_1085 ();
 sg13g2_decap_8 FILLER_0_3_1092 ();
 sg13g2_decap_8 FILLER_0_3_1099 ();
 sg13g2_decap_8 FILLER_0_3_1106 ();
 sg13g2_decap_8 FILLER_0_3_1113 ();
 sg13g2_decap_8 FILLER_0_3_1120 ();
 sg13g2_decap_8 FILLER_0_3_1127 ();
 sg13g2_decap_8 FILLER_0_3_1134 ();
 sg13g2_decap_8 FILLER_0_3_1141 ();
 sg13g2_decap_8 FILLER_0_3_1148 ();
 sg13g2_decap_8 FILLER_0_3_1155 ();
 sg13g2_decap_8 FILLER_0_3_1162 ();
 sg13g2_decap_8 FILLER_0_3_1169 ();
 sg13g2_decap_8 FILLER_0_3_1176 ();
 sg13g2_decap_8 FILLER_0_3_1183 ();
 sg13g2_decap_8 FILLER_0_3_1190 ();
 sg13g2_decap_8 FILLER_0_3_1197 ();
 sg13g2_decap_8 FILLER_0_3_1204 ();
 sg13g2_decap_8 FILLER_0_3_1211 ();
 sg13g2_decap_8 FILLER_0_3_1218 ();
 sg13g2_fill_2 FILLER_0_3_1225 ();
 sg13g2_fill_1 FILLER_0_3_1227 ();
 sg13g2_decap_8 FILLER_0_4_0 ();
 sg13g2_decap_8 FILLER_0_4_7 ();
 sg13g2_decap_8 FILLER_0_4_14 ();
 sg13g2_decap_8 FILLER_0_4_21 ();
 sg13g2_decap_8 FILLER_0_4_28 ();
 sg13g2_decap_8 FILLER_0_4_35 ();
 sg13g2_decap_8 FILLER_0_4_42 ();
 sg13g2_decap_8 FILLER_0_4_49 ();
 sg13g2_decap_8 FILLER_0_4_56 ();
 sg13g2_decap_8 FILLER_0_4_63 ();
 sg13g2_decap_8 FILLER_0_4_70 ();
 sg13g2_decap_8 FILLER_0_4_77 ();
 sg13g2_decap_8 FILLER_0_4_84 ();
 sg13g2_decap_8 FILLER_0_4_91 ();
 sg13g2_decap_8 FILLER_0_4_98 ();
 sg13g2_decap_8 FILLER_0_4_105 ();
 sg13g2_decap_8 FILLER_0_4_112 ();
 sg13g2_decap_8 FILLER_0_4_119 ();
 sg13g2_decap_8 FILLER_0_4_126 ();
 sg13g2_decap_8 FILLER_0_4_133 ();
 sg13g2_decap_8 FILLER_0_4_140 ();
 sg13g2_decap_8 FILLER_0_4_147 ();
 sg13g2_decap_8 FILLER_0_4_154 ();
 sg13g2_decap_8 FILLER_0_4_161 ();
 sg13g2_decap_8 FILLER_0_4_168 ();
 sg13g2_decap_8 FILLER_0_4_175 ();
 sg13g2_decap_8 FILLER_0_4_182 ();
 sg13g2_decap_8 FILLER_0_4_189 ();
 sg13g2_decap_8 FILLER_0_4_196 ();
 sg13g2_decap_8 FILLER_0_4_203 ();
 sg13g2_decap_8 FILLER_0_4_210 ();
 sg13g2_decap_8 FILLER_0_4_217 ();
 sg13g2_decap_8 FILLER_0_4_224 ();
 sg13g2_decap_8 FILLER_0_4_231 ();
 sg13g2_decap_8 FILLER_0_4_238 ();
 sg13g2_decap_8 FILLER_0_4_245 ();
 sg13g2_decap_8 FILLER_0_4_252 ();
 sg13g2_decap_8 FILLER_0_4_259 ();
 sg13g2_decap_8 FILLER_0_4_266 ();
 sg13g2_decap_8 FILLER_0_4_273 ();
 sg13g2_decap_8 FILLER_0_4_280 ();
 sg13g2_decap_8 FILLER_0_4_287 ();
 sg13g2_decap_8 FILLER_0_4_294 ();
 sg13g2_decap_8 FILLER_0_4_301 ();
 sg13g2_decap_8 FILLER_0_4_308 ();
 sg13g2_decap_8 FILLER_0_4_315 ();
 sg13g2_decap_8 FILLER_0_4_322 ();
 sg13g2_decap_8 FILLER_0_4_329 ();
 sg13g2_decap_8 FILLER_0_4_336 ();
 sg13g2_decap_8 FILLER_0_4_343 ();
 sg13g2_decap_8 FILLER_0_4_350 ();
 sg13g2_decap_8 FILLER_0_4_357 ();
 sg13g2_decap_8 FILLER_0_4_364 ();
 sg13g2_decap_8 FILLER_0_4_371 ();
 sg13g2_decap_8 FILLER_0_4_378 ();
 sg13g2_decap_8 FILLER_0_4_385 ();
 sg13g2_decap_8 FILLER_0_4_392 ();
 sg13g2_decap_8 FILLER_0_4_399 ();
 sg13g2_decap_8 FILLER_0_4_406 ();
 sg13g2_decap_8 FILLER_0_4_413 ();
 sg13g2_decap_8 FILLER_0_4_420 ();
 sg13g2_decap_8 FILLER_0_4_427 ();
 sg13g2_decap_8 FILLER_0_4_434 ();
 sg13g2_decap_8 FILLER_0_4_441 ();
 sg13g2_decap_8 FILLER_0_4_448 ();
 sg13g2_decap_8 FILLER_0_4_455 ();
 sg13g2_decap_8 FILLER_0_4_462 ();
 sg13g2_decap_8 FILLER_0_4_469 ();
 sg13g2_decap_8 FILLER_0_4_476 ();
 sg13g2_decap_8 FILLER_0_4_483 ();
 sg13g2_decap_8 FILLER_0_4_490 ();
 sg13g2_decap_8 FILLER_0_4_497 ();
 sg13g2_decap_8 FILLER_0_4_504 ();
 sg13g2_decap_8 FILLER_0_4_511 ();
 sg13g2_decap_8 FILLER_0_4_518 ();
 sg13g2_decap_8 FILLER_0_4_525 ();
 sg13g2_decap_8 FILLER_0_4_532 ();
 sg13g2_decap_8 FILLER_0_4_539 ();
 sg13g2_decap_8 FILLER_0_4_546 ();
 sg13g2_decap_8 FILLER_0_4_553 ();
 sg13g2_decap_8 FILLER_0_4_560 ();
 sg13g2_decap_8 FILLER_0_4_567 ();
 sg13g2_decap_8 FILLER_0_4_574 ();
 sg13g2_decap_8 FILLER_0_4_581 ();
 sg13g2_decap_8 FILLER_0_4_588 ();
 sg13g2_decap_8 FILLER_0_4_595 ();
 sg13g2_decap_8 FILLER_0_4_602 ();
 sg13g2_decap_8 FILLER_0_4_609 ();
 sg13g2_decap_8 FILLER_0_4_616 ();
 sg13g2_decap_8 FILLER_0_4_623 ();
 sg13g2_decap_8 FILLER_0_4_630 ();
 sg13g2_decap_8 FILLER_0_4_637 ();
 sg13g2_decap_8 FILLER_0_4_644 ();
 sg13g2_decap_8 FILLER_0_4_651 ();
 sg13g2_decap_8 FILLER_0_4_658 ();
 sg13g2_decap_8 FILLER_0_4_665 ();
 sg13g2_decap_8 FILLER_0_4_672 ();
 sg13g2_decap_8 FILLER_0_4_679 ();
 sg13g2_decap_8 FILLER_0_4_686 ();
 sg13g2_decap_8 FILLER_0_4_693 ();
 sg13g2_decap_8 FILLER_0_4_700 ();
 sg13g2_decap_8 FILLER_0_4_707 ();
 sg13g2_decap_8 FILLER_0_4_714 ();
 sg13g2_decap_8 FILLER_0_4_721 ();
 sg13g2_decap_8 FILLER_0_4_728 ();
 sg13g2_decap_8 FILLER_0_4_735 ();
 sg13g2_decap_8 FILLER_0_4_742 ();
 sg13g2_decap_8 FILLER_0_4_749 ();
 sg13g2_decap_8 FILLER_0_4_756 ();
 sg13g2_decap_8 FILLER_0_4_763 ();
 sg13g2_decap_8 FILLER_0_4_770 ();
 sg13g2_decap_8 FILLER_0_4_777 ();
 sg13g2_decap_8 FILLER_0_4_784 ();
 sg13g2_decap_8 FILLER_0_4_791 ();
 sg13g2_decap_8 FILLER_0_4_798 ();
 sg13g2_decap_8 FILLER_0_4_805 ();
 sg13g2_decap_8 FILLER_0_4_812 ();
 sg13g2_decap_8 FILLER_0_4_819 ();
 sg13g2_decap_8 FILLER_0_4_826 ();
 sg13g2_decap_8 FILLER_0_4_833 ();
 sg13g2_decap_8 FILLER_0_4_840 ();
 sg13g2_decap_8 FILLER_0_4_847 ();
 sg13g2_decap_8 FILLER_0_4_854 ();
 sg13g2_decap_8 FILLER_0_4_861 ();
 sg13g2_decap_8 FILLER_0_4_868 ();
 sg13g2_decap_8 FILLER_0_4_875 ();
 sg13g2_decap_8 FILLER_0_4_882 ();
 sg13g2_decap_8 FILLER_0_4_889 ();
 sg13g2_decap_8 FILLER_0_4_896 ();
 sg13g2_decap_8 FILLER_0_4_903 ();
 sg13g2_decap_8 FILLER_0_4_910 ();
 sg13g2_decap_8 FILLER_0_4_917 ();
 sg13g2_decap_8 FILLER_0_4_924 ();
 sg13g2_decap_8 FILLER_0_4_931 ();
 sg13g2_decap_8 FILLER_0_4_938 ();
 sg13g2_decap_8 FILLER_0_4_945 ();
 sg13g2_decap_8 FILLER_0_4_952 ();
 sg13g2_decap_8 FILLER_0_4_959 ();
 sg13g2_decap_8 FILLER_0_4_966 ();
 sg13g2_decap_8 FILLER_0_4_973 ();
 sg13g2_decap_8 FILLER_0_4_980 ();
 sg13g2_decap_8 FILLER_0_4_987 ();
 sg13g2_decap_8 FILLER_0_4_994 ();
 sg13g2_decap_8 FILLER_0_4_1001 ();
 sg13g2_decap_8 FILLER_0_4_1008 ();
 sg13g2_decap_8 FILLER_0_4_1015 ();
 sg13g2_decap_8 FILLER_0_4_1022 ();
 sg13g2_decap_8 FILLER_0_4_1029 ();
 sg13g2_decap_8 FILLER_0_4_1036 ();
 sg13g2_decap_8 FILLER_0_4_1043 ();
 sg13g2_decap_8 FILLER_0_4_1050 ();
 sg13g2_decap_8 FILLER_0_4_1057 ();
 sg13g2_decap_8 FILLER_0_4_1064 ();
 sg13g2_decap_8 FILLER_0_4_1071 ();
 sg13g2_decap_8 FILLER_0_4_1078 ();
 sg13g2_decap_8 FILLER_0_4_1085 ();
 sg13g2_decap_8 FILLER_0_4_1092 ();
 sg13g2_decap_8 FILLER_0_4_1099 ();
 sg13g2_decap_8 FILLER_0_4_1106 ();
 sg13g2_decap_8 FILLER_0_4_1113 ();
 sg13g2_decap_8 FILLER_0_4_1120 ();
 sg13g2_decap_8 FILLER_0_4_1127 ();
 sg13g2_decap_8 FILLER_0_4_1134 ();
 sg13g2_decap_8 FILLER_0_4_1141 ();
 sg13g2_decap_8 FILLER_0_4_1148 ();
 sg13g2_decap_8 FILLER_0_4_1155 ();
 sg13g2_decap_8 FILLER_0_4_1162 ();
 sg13g2_decap_8 FILLER_0_4_1169 ();
 sg13g2_decap_8 FILLER_0_4_1176 ();
 sg13g2_decap_8 FILLER_0_4_1183 ();
 sg13g2_decap_8 FILLER_0_4_1190 ();
 sg13g2_decap_8 FILLER_0_4_1197 ();
 sg13g2_decap_8 FILLER_0_4_1204 ();
 sg13g2_decap_8 FILLER_0_4_1211 ();
 sg13g2_decap_8 FILLER_0_4_1218 ();
 sg13g2_fill_2 FILLER_0_4_1225 ();
 sg13g2_fill_1 FILLER_0_4_1227 ();
 sg13g2_decap_8 FILLER_0_5_0 ();
 sg13g2_decap_8 FILLER_0_5_7 ();
 sg13g2_decap_8 FILLER_0_5_14 ();
 sg13g2_decap_8 FILLER_0_5_21 ();
 sg13g2_decap_8 FILLER_0_5_28 ();
 sg13g2_decap_8 FILLER_0_5_35 ();
 sg13g2_decap_8 FILLER_0_5_42 ();
 sg13g2_decap_8 FILLER_0_5_49 ();
 sg13g2_decap_8 FILLER_0_5_56 ();
 sg13g2_decap_8 FILLER_0_5_63 ();
 sg13g2_decap_8 FILLER_0_5_70 ();
 sg13g2_decap_8 FILLER_0_5_77 ();
 sg13g2_decap_8 FILLER_0_5_84 ();
 sg13g2_decap_8 FILLER_0_5_91 ();
 sg13g2_decap_8 FILLER_0_5_98 ();
 sg13g2_decap_8 FILLER_0_5_105 ();
 sg13g2_decap_8 FILLER_0_5_112 ();
 sg13g2_decap_8 FILLER_0_5_119 ();
 sg13g2_decap_8 FILLER_0_5_126 ();
 sg13g2_decap_8 FILLER_0_5_133 ();
 sg13g2_decap_8 FILLER_0_5_140 ();
 sg13g2_decap_8 FILLER_0_5_147 ();
 sg13g2_decap_8 FILLER_0_5_154 ();
 sg13g2_decap_8 FILLER_0_5_161 ();
 sg13g2_decap_8 FILLER_0_5_168 ();
 sg13g2_decap_8 FILLER_0_5_175 ();
 sg13g2_decap_8 FILLER_0_5_182 ();
 sg13g2_decap_8 FILLER_0_5_189 ();
 sg13g2_decap_8 FILLER_0_5_196 ();
 sg13g2_decap_8 FILLER_0_5_203 ();
 sg13g2_decap_8 FILLER_0_5_210 ();
 sg13g2_decap_8 FILLER_0_5_217 ();
 sg13g2_decap_8 FILLER_0_5_224 ();
 sg13g2_decap_8 FILLER_0_5_231 ();
 sg13g2_decap_8 FILLER_0_5_238 ();
 sg13g2_decap_8 FILLER_0_5_245 ();
 sg13g2_decap_8 FILLER_0_5_252 ();
 sg13g2_decap_8 FILLER_0_5_259 ();
 sg13g2_decap_8 FILLER_0_5_266 ();
 sg13g2_decap_8 FILLER_0_5_273 ();
 sg13g2_decap_8 FILLER_0_5_280 ();
 sg13g2_decap_8 FILLER_0_5_287 ();
 sg13g2_decap_8 FILLER_0_5_294 ();
 sg13g2_decap_8 FILLER_0_5_301 ();
 sg13g2_decap_8 FILLER_0_5_308 ();
 sg13g2_decap_8 FILLER_0_5_315 ();
 sg13g2_decap_8 FILLER_0_5_322 ();
 sg13g2_decap_8 FILLER_0_5_329 ();
 sg13g2_decap_8 FILLER_0_5_336 ();
 sg13g2_decap_8 FILLER_0_5_343 ();
 sg13g2_decap_8 FILLER_0_5_350 ();
 sg13g2_decap_8 FILLER_0_5_357 ();
 sg13g2_decap_8 FILLER_0_5_364 ();
 sg13g2_decap_8 FILLER_0_5_371 ();
 sg13g2_decap_8 FILLER_0_5_378 ();
 sg13g2_decap_8 FILLER_0_5_385 ();
 sg13g2_decap_8 FILLER_0_5_392 ();
 sg13g2_decap_8 FILLER_0_5_399 ();
 sg13g2_decap_8 FILLER_0_5_406 ();
 sg13g2_decap_8 FILLER_0_5_413 ();
 sg13g2_decap_8 FILLER_0_5_420 ();
 sg13g2_decap_8 FILLER_0_5_427 ();
 sg13g2_decap_8 FILLER_0_5_434 ();
 sg13g2_decap_8 FILLER_0_5_441 ();
 sg13g2_decap_8 FILLER_0_5_448 ();
 sg13g2_decap_8 FILLER_0_5_455 ();
 sg13g2_decap_8 FILLER_0_5_462 ();
 sg13g2_decap_8 FILLER_0_5_469 ();
 sg13g2_decap_8 FILLER_0_5_476 ();
 sg13g2_decap_8 FILLER_0_5_483 ();
 sg13g2_decap_8 FILLER_0_5_490 ();
 sg13g2_decap_8 FILLER_0_5_497 ();
 sg13g2_decap_8 FILLER_0_5_504 ();
 sg13g2_decap_8 FILLER_0_5_511 ();
 sg13g2_decap_8 FILLER_0_5_518 ();
 sg13g2_decap_8 FILLER_0_5_525 ();
 sg13g2_decap_8 FILLER_0_5_532 ();
 sg13g2_decap_8 FILLER_0_5_539 ();
 sg13g2_decap_8 FILLER_0_5_546 ();
 sg13g2_decap_8 FILLER_0_5_553 ();
 sg13g2_decap_8 FILLER_0_5_560 ();
 sg13g2_decap_8 FILLER_0_5_567 ();
 sg13g2_decap_8 FILLER_0_5_574 ();
 sg13g2_decap_8 FILLER_0_5_581 ();
 sg13g2_decap_8 FILLER_0_5_588 ();
 sg13g2_decap_8 FILLER_0_5_595 ();
 sg13g2_decap_8 FILLER_0_5_602 ();
 sg13g2_decap_8 FILLER_0_5_609 ();
 sg13g2_decap_8 FILLER_0_5_616 ();
 sg13g2_decap_8 FILLER_0_5_623 ();
 sg13g2_decap_8 FILLER_0_5_630 ();
 sg13g2_decap_8 FILLER_0_5_637 ();
 sg13g2_decap_8 FILLER_0_5_644 ();
 sg13g2_decap_8 FILLER_0_5_651 ();
 sg13g2_decap_8 FILLER_0_5_658 ();
 sg13g2_decap_8 FILLER_0_5_665 ();
 sg13g2_decap_8 FILLER_0_5_672 ();
 sg13g2_decap_8 FILLER_0_5_679 ();
 sg13g2_decap_8 FILLER_0_5_686 ();
 sg13g2_decap_8 FILLER_0_5_693 ();
 sg13g2_decap_8 FILLER_0_5_700 ();
 sg13g2_decap_8 FILLER_0_5_707 ();
 sg13g2_decap_8 FILLER_0_5_714 ();
 sg13g2_decap_8 FILLER_0_5_721 ();
 sg13g2_decap_8 FILLER_0_5_728 ();
 sg13g2_decap_8 FILLER_0_5_735 ();
 sg13g2_decap_8 FILLER_0_5_742 ();
 sg13g2_decap_8 FILLER_0_5_749 ();
 sg13g2_decap_8 FILLER_0_5_756 ();
 sg13g2_decap_8 FILLER_0_5_763 ();
 sg13g2_decap_8 FILLER_0_5_770 ();
 sg13g2_decap_8 FILLER_0_5_777 ();
 sg13g2_decap_8 FILLER_0_5_784 ();
 sg13g2_decap_8 FILLER_0_5_791 ();
 sg13g2_decap_8 FILLER_0_5_798 ();
 sg13g2_decap_8 FILLER_0_5_805 ();
 sg13g2_decap_8 FILLER_0_5_812 ();
 sg13g2_decap_8 FILLER_0_5_819 ();
 sg13g2_decap_8 FILLER_0_5_826 ();
 sg13g2_decap_8 FILLER_0_5_833 ();
 sg13g2_decap_8 FILLER_0_5_840 ();
 sg13g2_decap_8 FILLER_0_5_847 ();
 sg13g2_decap_8 FILLER_0_5_854 ();
 sg13g2_decap_8 FILLER_0_5_861 ();
 sg13g2_decap_8 FILLER_0_5_868 ();
 sg13g2_decap_8 FILLER_0_5_875 ();
 sg13g2_decap_8 FILLER_0_5_882 ();
 sg13g2_decap_8 FILLER_0_5_889 ();
 sg13g2_decap_8 FILLER_0_5_896 ();
 sg13g2_decap_8 FILLER_0_5_903 ();
 sg13g2_decap_8 FILLER_0_5_910 ();
 sg13g2_decap_8 FILLER_0_5_917 ();
 sg13g2_decap_8 FILLER_0_5_924 ();
 sg13g2_decap_8 FILLER_0_5_931 ();
 sg13g2_decap_8 FILLER_0_5_938 ();
 sg13g2_decap_8 FILLER_0_5_945 ();
 sg13g2_decap_8 FILLER_0_5_952 ();
 sg13g2_decap_8 FILLER_0_5_959 ();
 sg13g2_decap_8 FILLER_0_5_966 ();
 sg13g2_decap_8 FILLER_0_5_973 ();
 sg13g2_decap_8 FILLER_0_5_980 ();
 sg13g2_decap_8 FILLER_0_5_987 ();
 sg13g2_decap_8 FILLER_0_5_994 ();
 sg13g2_decap_8 FILLER_0_5_1001 ();
 sg13g2_decap_8 FILLER_0_5_1008 ();
 sg13g2_decap_8 FILLER_0_5_1015 ();
 sg13g2_decap_8 FILLER_0_5_1022 ();
 sg13g2_decap_8 FILLER_0_5_1029 ();
 sg13g2_decap_8 FILLER_0_5_1036 ();
 sg13g2_decap_8 FILLER_0_5_1043 ();
 sg13g2_decap_8 FILLER_0_5_1050 ();
 sg13g2_decap_8 FILLER_0_5_1057 ();
 sg13g2_decap_8 FILLER_0_5_1064 ();
 sg13g2_decap_8 FILLER_0_5_1071 ();
 sg13g2_decap_8 FILLER_0_5_1078 ();
 sg13g2_decap_8 FILLER_0_5_1085 ();
 sg13g2_decap_8 FILLER_0_5_1092 ();
 sg13g2_decap_8 FILLER_0_5_1099 ();
 sg13g2_decap_8 FILLER_0_5_1106 ();
 sg13g2_decap_8 FILLER_0_5_1113 ();
 sg13g2_decap_8 FILLER_0_5_1120 ();
 sg13g2_decap_8 FILLER_0_5_1127 ();
 sg13g2_decap_8 FILLER_0_5_1134 ();
 sg13g2_decap_8 FILLER_0_5_1141 ();
 sg13g2_decap_8 FILLER_0_5_1148 ();
 sg13g2_decap_8 FILLER_0_5_1155 ();
 sg13g2_decap_8 FILLER_0_5_1162 ();
 sg13g2_decap_8 FILLER_0_5_1169 ();
 sg13g2_decap_8 FILLER_0_5_1176 ();
 sg13g2_decap_8 FILLER_0_5_1183 ();
 sg13g2_decap_8 FILLER_0_5_1190 ();
 sg13g2_decap_8 FILLER_0_5_1197 ();
 sg13g2_decap_8 FILLER_0_5_1204 ();
 sg13g2_decap_8 FILLER_0_5_1211 ();
 sg13g2_decap_8 FILLER_0_5_1218 ();
 sg13g2_fill_2 FILLER_0_5_1225 ();
 sg13g2_fill_1 FILLER_0_5_1227 ();
 sg13g2_decap_8 FILLER_0_6_0 ();
 sg13g2_decap_8 FILLER_0_6_7 ();
 sg13g2_decap_8 FILLER_0_6_14 ();
 sg13g2_decap_8 FILLER_0_6_21 ();
 sg13g2_decap_8 FILLER_0_6_28 ();
 sg13g2_decap_8 FILLER_0_6_35 ();
 sg13g2_decap_8 FILLER_0_6_42 ();
 sg13g2_decap_8 FILLER_0_6_49 ();
 sg13g2_decap_8 FILLER_0_6_56 ();
 sg13g2_decap_8 FILLER_0_6_63 ();
 sg13g2_decap_8 FILLER_0_6_70 ();
 sg13g2_decap_8 FILLER_0_6_77 ();
 sg13g2_decap_8 FILLER_0_6_84 ();
 sg13g2_decap_8 FILLER_0_6_91 ();
 sg13g2_decap_8 FILLER_0_6_98 ();
 sg13g2_decap_8 FILLER_0_6_105 ();
 sg13g2_decap_8 FILLER_0_6_112 ();
 sg13g2_decap_8 FILLER_0_6_119 ();
 sg13g2_decap_8 FILLER_0_6_126 ();
 sg13g2_decap_8 FILLER_0_6_133 ();
 sg13g2_decap_8 FILLER_0_6_140 ();
 sg13g2_decap_8 FILLER_0_6_147 ();
 sg13g2_decap_8 FILLER_0_6_154 ();
 sg13g2_decap_8 FILLER_0_6_161 ();
 sg13g2_decap_8 FILLER_0_6_168 ();
 sg13g2_decap_8 FILLER_0_6_175 ();
 sg13g2_decap_8 FILLER_0_6_182 ();
 sg13g2_decap_8 FILLER_0_6_189 ();
 sg13g2_decap_8 FILLER_0_6_196 ();
 sg13g2_decap_8 FILLER_0_6_203 ();
 sg13g2_decap_8 FILLER_0_6_210 ();
 sg13g2_decap_8 FILLER_0_6_217 ();
 sg13g2_decap_8 FILLER_0_6_224 ();
 sg13g2_decap_8 FILLER_0_6_231 ();
 sg13g2_decap_8 FILLER_0_6_238 ();
 sg13g2_decap_8 FILLER_0_6_245 ();
 sg13g2_decap_8 FILLER_0_6_252 ();
 sg13g2_decap_8 FILLER_0_6_259 ();
 sg13g2_decap_8 FILLER_0_6_266 ();
 sg13g2_decap_8 FILLER_0_6_273 ();
 sg13g2_decap_8 FILLER_0_6_280 ();
 sg13g2_decap_8 FILLER_0_6_287 ();
 sg13g2_decap_8 FILLER_0_6_294 ();
 sg13g2_decap_8 FILLER_0_6_301 ();
 sg13g2_decap_8 FILLER_0_6_308 ();
 sg13g2_decap_8 FILLER_0_6_315 ();
 sg13g2_decap_8 FILLER_0_6_322 ();
 sg13g2_decap_8 FILLER_0_6_329 ();
 sg13g2_decap_8 FILLER_0_6_336 ();
 sg13g2_decap_8 FILLER_0_6_343 ();
 sg13g2_decap_8 FILLER_0_6_350 ();
 sg13g2_decap_8 FILLER_0_6_357 ();
 sg13g2_decap_8 FILLER_0_6_364 ();
 sg13g2_decap_8 FILLER_0_6_371 ();
 sg13g2_decap_8 FILLER_0_6_378 ();
 sg13g2_decap_8 FILLER_0_6_385 ();
 sg13g2_decap_8 FILLER_0_6_392 ();
 sg13g2_decap_8 FILLER_0_6_399 ();
 sg13g2_decap_8 FILLER_0_6_406 ();
 sg13g2_decap_8 FILLER_0_6_413 ();
 sg13g2_decap_8 FILLER_0_6_420 ();
 sg13g2_decap_8 FILLER_0_6_427 ();
 sg13g2_decap_8 FILLER_0_6_434 ();
 sg13g2_decap_8 FILLER_0_6_441 ();
 sg13g2_decap_8 FILLER_0_6_448 ();
 sg13g2_decap_8 FILLER_0_6_455 ();
 sg13g2_decap_8 FILLER_0_6_462 ();
 sg13g2_decap_8 FILLER_0_6_469 ();
 sg13g2_decap_8 FILLER_0_6_476 ();
 sg13g2_decap_8 FILLER_0_6_483 ();
 sg13g2_decap_8 FILLER_0_6_490 ();
 sg13g2_decap_8 FILLER_0_6_497 ();
 sg13g2_decap_8 FILLER_0_6_504 ();
 sg13g2_decap_8 FILLER_0_6_511 ();
 sg13g2_decap_8 FILLER_0_6_518 ();
 sg13g2_decap_8 FILLER_0_6_525 ();
 sg13g2_decap_8 FILLER_0_6_532 ();
 sg13g2_decap_8 FILLER_0_6_539 ();
 sg13g2_decap_8 FILLER_0_6_546 ();
 sg13g2_decap_8 FILLER_0_6_553 ();
 sg13g2_decap_8 FILLER_0_6_560 ();
 sg13g2_decap_8 FILLER_0_6_567 ();
 sg13g2_decap_8 FILLER_0_6_574 ();
 sg13g2_decap_8 FILLER_0_6_581 ();
 sg13g2_decap_8 FILLER_0_6_588 ();
 sg13g2_decap_8 FILLER_0_6_595 ();
 sg13g2_decap_8 FILLER_0_6_602 ();
 sg13g2_decap_8 FILLER_0_6_609 ();
 sg13g2_decap_8 FILLER_0_6_616 ();
 sg13g2_decap_8 FILLER_0_6_623 ();
 sg13g2_decap_8 FILLER_0_6_630 ();
 sg13g2_decap_8 FILLER_0_6_637 ();
 sg13g2_decap_8 FILLER_0_6_644 ();
 sg13g2_decap_8 FILLER_0_6_651 ();
 sg13g2_decap_8 FILLER_0_6_658 ();
 sg13g2_decap_8 FILLER_0_6_665 ();
 sg13g2_decap_8 FILLER_0_6_672 ();
 sg13g2_decap_8 FILLER_0_6_679 ();
 sg13g2_decap_8 FILLER_0_6_686 ();
 sg13g2_decap_8 FILLER_0_6_693 ();
 sg13g2_decap_8 FILLER_0_6_700 ();
 sg13g2_decap_8 FILLER_0_6_707 ();
 sg13g2_decap_8 FILLER_0_6_714 ();
 sg13g2_decap_8 FILLER_0_6_721 ();
 sg13g2_decap_8 FILLER_0_6_728 ();
 sg13g2_decap_8 FILLER_0_6_735 ();
 sg13g2_decap_8 FILLER_0_6_742 ();
 sg13g2_decap_8 FILLER_0_6_749 ();
 sg13g2_decap_8 FILLER_0_6_756 ();
 sg13g2_decap_8 FILLER_0_6_763 ();
 sg13g2_decap_8 FILLER_0_6_770 ();
 sg13g2_decap_8 FILLER_0_6_777 ();
 sg13g2_decap_8 FILLER_0_6_784 ();
 sg13g2_decap_8 FILLER_0_6_791 ();
 sg13g2_decap_8 FILLER_0_6_798 ();
 sg13g2_decap_8 FILLER_0_6_805 ();
 sg13g2_decap_8 FILLER_0_6_812 ();
 sg13g2_decap_8 FILLER_0_6_819 ();
 sg13g2_decap_8 FILLER_0_6_826 ();
 sg13g2_decap_8 FILLER_0_6_833 ();
 sg13g2_decap_8 FILLER_0_6_840 ();
 sg13g2_decap_8 FILLER_0_6_847 ();
 sg13g2_decap_8 FILLER_0_6_854 ();
 sg13g2_decap_8 FILLER_0_6_861 ();
 sg13g2_decap_8 FILLER_0_6_868 ();
 sg13g2_decap_8 FILLER_0_6_875 ();
 sg13g2_decap_8 FILLER_0_6_882 ();
 sg13g2_decap_8 FILLER_0_6_889 ();
 sg13g2_decap_8 FILLER_0_6_896 ();
 sg13g2_decap_8 FILLER_0_6_903 ();
 sg13g2_decap_8 FILLER_0_6_910 ();
 sg13g2_decap_8 FILLER_0_6_917 ();
 sg13g2_decap_8 FILLER_0_6_924 ();
 sg13g2_decap_8 FILLER_0_6_931 ();
 sg13g2_decap_8 FILLER_0_6_938 ();
 sg13g2_decap_8 FILLER_0_6_945 ();
 sg13g2_decap_8 FILLER_0_6_952 ();
 sg13g2_decap_8 FILLER_0_6_959 ();
 sg13g2_decap_8 FILLER_0_6_966 ();
 sg13g2_decap_8 FILLER_0_6_973 ();
 sg13g2_decap_8 FILLER_0_6_980 ();
 sg13g2_decap_8 FILLER_0_6_987 ();
 sg13g2_decap_8 FILLER_0_6_994 ();
 sg13g2_decap_8 FILLER_0_6_1001 ();
 sg13g2_decap_8 FILLER_0_6_1008 ();
 sg13g2_decap_8 FILLER_0_6_1015 ();
 sg13g2_decap_8 FILLER_0_6_1022 ();
 sg13g2_decap_8 FILLER_0_6_1029 ();
 sg13g2_decap_8 FILLER_0_6_1036 ();
 sg13g2_decap_8 FILLER_0_6_1043 ();
 sg13g2_decap_8 FILLER_0_6_1050 ();
 sg13g2_decap_8 FILLER_0_6_1057 ();
 sg13g2_decap_8 FILLER_0_6_1064 ();
 sg13g2_decap_8 FILLER_0_6_1071 ();
 sg13g2_decap_8 FILLER_0_6_1078 ();
 sg13g2_decap_8 FILLER_0_6_1085 ();
 sg13g2_decap_8 FILLER_0_6_1092 ();
 sg13g2_decap_8 FILLER_0_6_1099 ();
 sg13g2_decap_8 FILLER_0_6_1106 ();
 sg13g2_decap_8 FILLER_0_6_1113 ();
 sg13g2_decap_8 FILLER_0_6_1120 ();
 sg13g2_decap_8 FILLER_0_6_1127 ();
 sg13g2_decap_8 FILLER_0_6_1134 ();
 sg13g2_decap_8 FILLER_0_6_1141 ();
 sg13g2_decap_8 FILLER_0_6_1148 ();
 sg13g2_decap_8 FILLER_0_6_1155 ();
 sg13g2_decap_8 FILLER_0_6_1162 ();
 sg13g2_decap_8 FILLER_0_6_1169 ();
 sg13g2_decap_8 FILLER_0_6_1176 ();
 sg13g2_decap_8 FILLER_0_6_1183 ();
 sg13g2_decap_8 FILLER_0_6_1190 ();
 sg13g2_decap_8 FILLER_0_6_1197 ();
 sg13g2_decap_8 FILLER_0_6_1204 ();
 sg13g2_decap_8 FILLER_0_6_1211 ();
 sg13g2_decap_8 FILLER_0_6_1218 ();
 sg13g2_fill_2 FILLER_0_6_1225 ();
 sg13g2_fill_1 FILLER_0_6_1227 ();
 sg13g2_decap_8 FILLER_0_7_0 ();
 sg13g2_decap_8 FILLER_0_7_7 ();
 sg13g2_decap_8 FILLER_0_7_14 ();
 sg13g2_decap_8 FILLER_0_7_21 ();
 sg13g2_decap_8 FILLER_0_7_28 ();
 sg13g2_decap_8 FILLER_0_7_35 ();
 sg13g2_decap_8 FILLER_0_7_42 ();
 sg13g2_decap_8 FILLER_0_7_49 ();
 sg13g2_decap_8 FILLER_0_7_56 ();
 sg13g2_decap_8 FILLER_0_7_63 ();
 sg13g2_decap_8 FILLER_0_7_70 ();
 sg13g2_decap_8 FILLER_0_7_77 ();
 sg13g2_decap_8 FILLER_0_7_84 ();
 sg13g2_decap_8 FILLER_0_7_91 ();
 sg13g2_decap_8 FILLER_0_7_98 ();
 sg13g2_decap_8 FILLER_0_7_105 ();
 sg13g2_decap_8 FILLER_0_7_112 ();
 sg13g2_decap_8 FILLER_0_7_119 ();
 sg13g2_decap_8 FILLER_0_7_126 ();
 sg13g2_decap_8 FILLER_0_7_133 ();
 sg13g2_decap_8 FILLER_0_7_140 ();
 sg13g2_decap_8 FILLER_0_7_147 ();
 sg13g2_decap_8 FILLER_0_7_154 ();
 sg13g2_decap_8 FILLER_0_7_161 ();
 sg13g2_decap_8 FILLER_0_7_168 ();
 sg13g2_decap_8 FILLER_0_7_175 ();
 sg13g2_decap_8 FILLER_0_7_182 ();
 sg13g2_decap_8 FILLER_0_7_189 ();
 sg13g2_decap_8 FILLER_0_7_196 ();
 sg13g2_decap_8 FILLER_0_7_203 ();
 sg13g2_decap_8 FILLER_0_7_210 ();
 sg13g2_decap_8 FILLER_0_7_217 ();
 sg13g2_decap_8 FILLER_0_7_224 ();
 sg13g2_decap_8 FILLER_0_7_231 ();
 sg13g2_decap_8 FILLER_0_7_238 ();
 sg13g2_decap_8 FILLER_0_7_245 ();
 sg13g2_decap_8 FILLER_0_7_252 ();
 sg13g2_decap_8 FILLER_0_7_259 ();
 sg13g2_decap_8 FILLER_0_7_266 ();
 sg13g2_decap_8 FILLER_0_7_273 ();
 sg13g2_decap_8 FILLER_0_7_280 ();
 sg13g2_decap_8 FILLER_0_7_287 ();
 sg13g2_decap_8 FILLER_0_7_294 ();
 sg13g2_decap_8 FILLER_0_7_301 ();
 sg13g2_decap_8 FILLER_0_7_308 ();
 sg13g2_decap_8 FILLER_0_7_315 ();
 sg13g2_decap_8 FILLER_0_7_322 ();
 sg13g2_decap_8 FILLER_0_7_329 ();
 sg13g2_decap_8 FILLER_0_7_336 ();
 sg13g2_decap_8 FILLER_0_7_343 ();
 sg13g2_decap_8 FILLER_0_7_350 ();
 sg13g2_decap_8 FILLER_0_7_357 ();
 sg13g2_decap_8 FILLER_0_7_364 ();
 sg13g2_decap_8 FILLER_0_7_371 ();
 sg13g2_decap_8 FILLER_0_7_378 ();
 sg13g2_decap_8 FILLER_0_7_385 ();
 sg13g2_decap_8 FILLER_0_7_392 ();
 sg13g2_decap_8 FILLER_0_7_399 ();
 sg13g2_decap_8 FILLER_0_7_406 ();
 sg13g2_decap_8 FILLER_0_7_413 ();
 sg13g2_decap_8 FILLER_0_7_420 ();
 sg13g2_decap_8 FILLER_0_7_427 ();
 sg13g2_decap_8 FILLER_0_7_434 ();
 sg13g2_decap_8 FILLER_0_7_441 ();
 sg13g2_decap_8 FILLER_0_7_448 ();
 sg13g2_decap_8 FILLER_0_7_455 ();
 sg13g2_decap_8 FILLER_0_7_462 ();
 sg13g2_decap_8 FILLER_0_7_469 ();
 sg13g2_decap_8 FILLER_0_7_476 ();
 sg13g2_decap_8 FILLER_0_7_483 ();
 sg13g2_decap_8 FILLER_0_7_490 ();
 sg13g2_decap_8 FILLER_0_7_497 ();
 sg13g2_decap_8 FILLER_0_7_504 ();
 sg13g2_decap_8 FILLER_0_7_511 ();
 sg13g2_decap_8 FILLER_0_7_518 ();
 sg13g2_decap_8 FILLER_0_7_525 ();
 sg13g2_decap_8 FILLER_0_7_532 ();
 sg13g2_decap_8 FILLER_0_7_539 ();
 sg13g2_decap_8 FILLER_0_7_546 ();
 sg13g2_decap_8 FILLER_0_7_553 ();
 sg13g2_decap_8 FILLER_0_7_560 ();
 sg13g2_decap_8 FILLER_0_7_567 ();
 sg13g2_decap_8 FILLER_0_7_574 ();
 sg13g2_decap_8 FILLER_0_7_581 ();
 sg13g2_decap_8 FILLER_0_7_588 ();
 sg13g2_decap_8 FILLER_0_7_595 ();
 sg13g2_decap_8 FILLER_0_7_602 ();
 sg13g2_decap_8 FILLER_0_7_609 ();
 sg13g2_decap_8 FILLER_0_7_616 ();
 sg13g2_decap_8 FILLER_0_7_623 ();
 sg13g2_decap_8 FILLER_0_7_630 ();
 sg13g2_decap_8 FILLER_0_7_637 ();
 sg13g2_decap_8 FILLER_0_7_644 ();
 sg13g2_decap_8 FILLER_0_7_651 ();
 sg13g2_decap_8 FILLER_0_7_658 ();
 sg13g2_decap_8 FILLER_0_7_665 ();
 sg13g2_decap_8 FILLER_0_7_672 ();
 sg13g2_decap_8 FILLER_0_7_679 ();
 sg13g2_decap_8 FILLER_0_7_686 ();
 sg13g2_decap_8 FILLER_0_7_693 ();
 sg13g2_decap_8 FILLER_0_7_700 ();
 sg13g2_decap_8 FILLER_0_7_707 ();
 sg13g2_decap_8 FILLER_0_7_714 ();
 sg13g2_decap_8 FILLER_0_7_721 ();
 sg13g2_decap_8 FILLER_0_7_728 ();
 sg13g2_decap_8 FILLER_0_7_735 ();
 sg13g2_decap_8 FILLER_0_7_742 ();
 sg13g2_decap_8 FILLER_0_7_749 ();
 sg13g2_decap_8 FILLER_0_7_756 ();
 sg13g2_decap_8 FILLER_0_7_763 ();
 sg13g2_decap_8 FILLER_0_7_770 ();
 sg13g2_decap_8 FILLER_0_7_777 ();
 sg13g2_decap_8 FILLER_0_7_784 ();
 sg13g2_decap_8 FILLER_0_7_791 ();
 sg13g2_decap_8 FILLER_0_7_798 ();
 sg13g2_decap_8 FILLER_0_7_805 ();
 sg13g2_decap_8 FILLER_0_7_812 ();
 sg13g2_decap_8 FILLER_0_7_819 ();
 sg13g2_decap_8 FILLER_0_7_826 ();
 sg13g2_decap_8 FILLER_0_7_833 ();
 sg13g2_decap_8 FILLER_0_7_840 ();
 sg13g2_decap_8 FILLER_0_7_847 ();
 sg13g2_decap_8 FILLER_0_7_854 ();
 sg13g2_decap_8 FILLER_0_7_861 ();
 sg13g2_decap_8 FILLER_0_7_868 ();
 sg13g2_decap_8 FILLER_0_7_875 ();
 sg13g2_decap_8 FILLER_0_7_882 ();
 sg13g2_decap_8 FILLER_0_7_889 ();
 sg13g2_decap_8 FILLER_0_7_896 ();
 sg13g2_decap_8 FILLER_0_7_903 ();
 sg13g2_decap_8 FILLER_0_7_910 ();
 sg13g2_decap_8 FILLER_0_7_917 ();
 sg13g2_decap_8 FILLER_0_7_924 ();
 sg13g2_decap_8 FILLER_0_7_931 ();
 sg13g2_decap_8 FILLER_0_7_938 ();
 sg13g2_decap_8 FILLER_0_7_945 ();
 sg13g2_decap_8 FILLER_0_7_952 ();
 sg13g2_decap_8 FILLER_0_7_959 ();
 sg13g2_decap_8 FILLER_0_7_966 ();
 sg13g2_decap_8 FILLER_0_7_973 ();
 sg13g2_decap_8 FILLER_0_7_980 ();
 sg13g2_decap_8 FILLER_0_7_987 ();
 sg13g2_decap_8 FILLER_0_7_994 ();
 sg13g2_decap_8 FILLER_0_7_1001 ();
 sg13g2_decap_8 FILLER_0_7_1008 ();
 sg13g2_decap_8 FILLER_0_7_1015 ();
 sg13g2_decap_8 FILLER_0_7_1022 ();
 sg13g2_decap_8 FILLER_0_7_1029 ();
 sg13g2_decap_8 FILLER_0_7_1036 ();
 sg13g2_decap_8 FILLER_0_7_1043 ();
 sg13g2_decap_8 FILLER_0_7_1050 ();
 sg13g2_decap_8 FILLER_0_7_1057 ();
 sg13g2_decap_8 FILLER_0_7_1064 ();
 sg13g2_decap_8 FILLER_0_7_1071 ();
 sg13g2_decap_8 FILLER_0_7_1078 ();
 sg13g2_decap_8 FILLER_0_7_1085 ();
 sg13g2_decap_8 FILLER_0_7_1092 ();
 sg13g2_decap_8 FILLER_0_7_1099 ();
 sg13g2_decap_8 FILLER_0_7_1106 ();
 sg13g2_decap_8 FILLER_0_7_1113 ();
 sg13g2_decap_8 FILLER_0_7_1120 ();
 sg13g2_decap_8 FILLER_0_7_1127 ();
 sg13g2_decap_8 FILLER_0_7_1134 ();
 sg13g2_decap_8 FILLER_0_7_1141 ();
 sg13g2_decap_8 FILLER_0_7_1148 ();
 sg13g2_decap_8 FILLER_0_7_1155 ();
 sg13g2_decap_8 FILLER_0_7_1162 ();
 sg13g2_decap_8 FILLER_0_7_1169 ();
 sg13g2_decap_8 FILLER_0_7_1176 ();
 sg13g2_decap_8 FILLER_0_7_1183 ();
 sg13g2_decap_8 FILLER_0_7_1190 ();
 sg13g2_decap_8 FILLER_0_7_1197 ();
 sg13g2_decap_8 FILLER_0_7_1204 ();
 sg13g2_decap_8 FILLER_0_7_1211 ();
 sg13g2_decap_8 FILLER_0_7_1218 ();
 sg13g2_fill_2 FILLER_0_7_1225 ();
 sg13g2_fill_1 FILLER_0_7_1227 ();
 sg13g2_decap_8 FILLER_0_8_0 ();
 sg13g2_decap_8 FILLER_0_8_7 ();
 sg13g2_decap_8 FILLER_0_8_14 ();
 sg13g2_decap_8 FILLER_0_8_21 ();
 sg13g2_decap_8 FILLER_0_8_28 ();
 sg13g2_decap_8 FILLER_0_8_35 ();
 sg13g2_decap_8 FILLER_0_8_42 ();
 sg13g2_decap_8 FILLER_0_8_49 ();
 sg13g2_decap_8 FILLER_0_8_56 ();
 sg13g2_decap_8 FILLER_0_8_63 ();
 sg13g2_decap_8 FILLER_0_8_70 ();
 sg13g2_decap_8 FILLER_0_8_77 ();
 sg13g2_decap_8 FILLER_0_8_84 ();
 sg13g2_decap_8 FILLER_0_8_91 ();
 sg13g2_decap_8 FILLER_0_8_98 ();
 sg13g2_decap_8 FILLER_0_8_105 ();
 sg13g2_decap_8 FILLER_0_8_112 ();
 sg13g2_decap_8 FILLER_0_8_119 ();
 sg13g2_decap_8 FILLER_0_8_126 ();
 sg13g2_decap_8 FILLER_0_8_133 ();
 sg13g2_decap_8 FILLER_0_8_140 ();
 sg13g2_decap_8 FILLER_0_8_147 ();
 sg13g2_decap_8 FILLER_0_8_154 ();
 sg13g2_decap_8 FILLER_0_8_161 ();
 sg13g2_decap_8 FILLER_0_8_168 ();
 sg13g2_decap_8 FILLER_0_8_175 ();
 sg13g2_decap_8 FILLER_0_8_182 ();
 sg13g2_decap_8 FILLER_0_8_189 ();
 sg13g2_decap_8 FILLER_0_8_196 ();
 sg13g2_decap_8 FILLER_0_8_203 ();
 sg13g2_decap_8 FILLER_0_8_210 ();
 sg13g2_decap_8 FILLER_0_8_217 ();
 sg13g2_decap_8 FILLER_0_8_224 ();
 sg13g2_decap_8 FILLER_0_8_231 ();
 sg13g2_decap_8 FILLER_0_8_238 ();
 sg13g2_decap_8 FILLER_0_8_245 ();
 sg13g2_decap_8 FILLER_0_8_252 ();
 sg13g2_decap_8 FILLER_0_8_259 ();
 sg13g2_decap_8 FILLER_0_8_266 ();
 sg13g2_decap_8 FILLER_0_8_273 ();
 sg13g2_decap_8 FILLER_0_8_280 ();
 sg13g2_decap_8 FILLER_0_8_287 ();
 sg13g2_decap_8 FILLER_0_8_294 ();
 sg13g2_decap_8 FILLER_0_8_301 ();
 sg13g2_decap_8 FILLER_0_8_308 ();
 sg13g2_decap_8 FILLER_0_8_315 ();
 sg13g2_decap_8 FILLER_0_8_322 ();
 sg13g2_decap_8 FILLER_0_8_329 ();
 sg13g2_decap_8 FILLER_0_8_336 ();
 sg13g2_decap_8 FILLER_0_8_343 ();
 sg13g2_decap_8 FILLER_0_8_350 ();
 sg13g2_decap_8 FILLER_0_8_357 ();
 sg13g2_decap_8 FILLER_0_8_364 ();
 sg13g2_decap_8 FILLER_0_8_371 ();
 sg13g2_decap_8 FILLER_0_8_378 ();
 sg13g2_decap_8 FILLER_0_8_385 ();
 sg13g2_decap_8 FILLER_0_8_392 ();
 sg13g2_decap_8 FILLER_0_8_399 ();
 sg13g2_decap_8 FILLER_0_8_406 ();
 sg13g2_decap_8 FILLER_0_8_413 ();
 sg13g2_decap_8 FILLER_0_8_420 ();
 sg13g2_decap_8 FILLER_0_8_427 ();
 sg13g2_decap_8 FILLER_0_8_434 ();
 sg13g2_decap_8 FILLER_0_8_441 ();
 sg13g2_decap_8 FILLER_0_8_448 ();
 sg13g2_decap_8 FILLER_0_8_455 ();
 sg13g2_decap_8 FILLER_0_8_462 ();
 sg13g2_decap_8 FILLER_0_8_469 ();
 sg13g2_decap_8 FILLER_0_8_476 ();
 sg13g2_decap_8 FILLER_0_8_483 ();
 sg13g2_decap_8 FILLER_0_8_490 ();
 sg13g2_decap_8 FILLER_0_8_497 ();
 sg13g2_decap_8 FILLER_0_8_504 ();
 sg13g2_decap_8 FILLER_0_8_511 ();
 sg13g2_decap_8 FILLER_0_8_518 ();
 sg13g2_decap_8 FILLER_0_8_525 ();
 sg13g2_decap_8 FILLER_0_8_532 ();
 sg13g2_decap_8 FILLER_0_8_539 ();
 sg13g2_decap_8 FILLER_0_8_546 ();
 sg13g2_decap_8 FILLER_0_8_553 ();
 sg13g2_decap_8 FILLER_0_8_560 ();
 sg13g2_decap_8 FILLER_0_8_567 ();
 sg13g2_decap_8 FILLER_0_8_574 ();
 sg13g2_decap_8 FILLER_0_8_581 ();
 sg13g2_decap_8 FILLER_0_8_588 ();
 sg13g2_decap_8 FILLER_0_8_595 ();
 sg13g2_decap_8 FILLER_0_8_602 ();
 sg13g2_decap_8 FILLER_0_8_609 ();
 sg13g2_decap_8 FILLER_0_8_616 ();
 sg13g2_decap_8 FILLER_0_8_623 ();
 sg13g2_decap_8 FILLER_0_8_630 ();
 sg13g2_decap_8 FILLER_0_8_637 ();
 sg13g2_decap_8 FILLER_0_8_644 ();
 sg13g2_decap_8 FILLER_0_8_651 ();
 sg13g2_decap_8 FILLER_0_8_658 ();
 sg13g2_decap_8 FILLER_0_8_665 ();
 sg13g2_decap_8 FILLER_0_8_672 ();
 sg13g2_decap_8 FILLER_0_8_679 ();
 sg13g2_decap_8 FILLER_0_8_686 ();
 sg13g2_decap_8 FILLER_0_8_693 ();
 sg13g2_decap_8 FILLER_0_8_700 ();
 sg13g2_decap_8 FILLER_0_8_707 ();
 sg13g2_decap_8 FILLER_0_8_714 ();
 sg13g2_decap_8 FILLER_0_8_721 ();
 sg13g2_decap_8 FILLER_0_8_728 ();
 sg13g2_decap_8 FILLER_0_8_735 ();
 sg13g2_decap_8 FILLER_0_8_742 ();
 sg13g2_decap_8 FILLER_0_8_749 ();
 sg13g2_decap_8 FILLER_0_8_756 ();
 sg13g2_decap_8 FILLER_0_8_763 ();
 sg13g2_decap_8 FILLER_0_8_770 ();
 sg13g2_decap_8 FILLER_0_8_777 ();
 sg13g2_decap_8 FILLER_0_8_784 ();
 sg13g2_decap_8 FILLER_0_8_791 ();
 sg13g2_decap_8 FILLER_0_8_798 ();
 sg13g2_decap_8 FILLER_0_8_805 ();
 sg13g2_decap_8 FILLER_0_8_812 ();
 sg13g2_decap_8 FILLER_0_8_819 ();
 sg13g2_decap_8 FILLER_0_8_826 ();
 sg13g2_decap_8 FILLER_0_8_833 ();
 sg13g2_decap_8 FILLER_0_8_840 ();
 sg13g2_decap_8 FILLER_0_8_847 ();
 sg13g2_decap_8 FILLER_0_8_854 ();
 sg13g2_decap_8 FILLER_0_8_861 ();
 sg13g2_decap_8 FILLER_0_8_868 ();
 sg13g2_decap_8 FILLER_0_8_875 ();
 sg13g2_decap_8 FILLER_0_8_882 ();
 sg13g2_decap_8 FILLER_0_8_889 ();
 sg13g2_decap_8 FILLER_0_8_896 ();
 sg13g2_decap_8 FILLER_0_8_903 ();
 sg13g2_decap_8 FILLER_0_8_910 ();
 sg13g2_decap_8 FILLER_0_8_917 ();
 sg13g2_decap_8 FILLER_0_8_924 ();
 sg13g2_decap_8 FILLER_0_8_931 ();
 sg13g2_decap_8 FILLER_0_8_938 ();
 sg13g2_decap_8 FILLER_0_8_945 ();
 sg13g2_decap_8 FILLER_0_8_952 ();
 sg13g2_decap_8 FILLER_0_8_959 ();
 sg13g2_decap_8 FILLER_0_8_966 ();
 sg13g2_decap_8 FILLER_0_8_973 ();
 sg13g2_decap_8 FILLER_0_8_980 ();
 sg13g2_decap_8 FILLER_0_8_987 ();
 sg13g2_decap_8 FILLER_0_8_994 ();
 sg13g2_decap_8 FILLER_0_8_1001 ();
 sg13g2_decap_8 FILLER_0_8_1008 ();
 sg13g2_decap_8 FILLER_0_8_1015 ();
 sg13g2_decap_8 FILLER_0_8_1022 ();
 sg13g2_decap_8 FILLER_0_8_1029 ();
 sg13g2_decap_8 FILLER_0_8_1036 ();
 sg13g2_decap_8 FILLER_0_8_1043 ();
 sg13g2_decap_8 FILLER_0_8_1050 ();
 sg13g2_decap_8 FILLER_0_8_1057 ();
 sg13g2_decap_8 FILLER_0_8_1064 ();
 sg13g2_decap_8 FILLER_0_8_1071 ();
 sg13g2_decap_8 FILLER_0_8_1078 ();
 sg13g2_decap_8 FILLER_0_8_1085 ();
 sg13g2_decap_8 FILLER_0_8_1092 ();
 sg13g2_decap_8 FILLER_0_8_1099 ();
 sg13g2_decap_8 FILLER_0_8_1106 ();
 sg13g2_decap_8 FILLER_0_8_1113 ();
 sg13g2_decap_8 FILLER_0_8_1120 ();
 sg13g2_decap_8 FILLER_0_8_1127 ();
 sg13g2_decap_8 FILLER_0_8_1134 ();
 sg13g2_decap_8 FILLER_0_8_1141 ();
 sg13g2_decap_8 FILLER_0_8_1148 ();
 sg13g2_decap_8 FILLER_0_8_1155 ();
 sg13g2_decap_8 FILLER_0_8_1162 ();
 sg13g2_decap_8 FILLER_0_8_1169 ();
 sg13g2_decap_8 FILLER_0_8_1176 ();
 sg13g2_decap_8 FILLER_0_8_1183 ();
 sg13g2_decap_8 FILLER_0_8_1190 ();
 sg13g2_decap_8 FILLER_0_8_1197 ();
 sg13g2_decap_8 FILLER_0_8_1204 ();
 sg13g2_decap_8 FILLER_0_8_1211 ();
 sg13g2_decap_8 FILLER_0_8_1218 ();
 sg13g2_fill_2 FILLER_0_8_1225 ();
 sg13g2_fill_1 FILLER_0_8_1227 ();
 sg13g2_decap_8 FILLER_0_9_0 ();
 sg13g2_decap_8 FILLER_0_9_7 ();
 sg13g2_decap_8 FILLER_0_9_14 ();
 sg13g2_decap_8 FILLER_0_9_21 ();
 sg13g2_decap_8 FILLER_0_9_28 ();
 sg13g2_decap_8 FILLER_0_9_35 ();
 sg13g2_decap_8 FILLER_0_9_42 ();
 sg13g2_decap_8 FILLER_0_9_49 ();
 sg13g2_decap_8 FILLER_0_9_56 ();
 sg13g2_decap_8 FILLER_0_9_63 ();
 sg13g2_decap_8 FILLER_0_9_70 ();
 sg13g2_decap_8 FILLER_0_9_77 ();
 sg13g2_decap_8 FILLER_0_9_84 ();
 sg13g2_decap_8 FILLER_0_9_91 ();
 sg13g2_decap_8 FILLER_0_9_98 ();
 sg13g2_decap_8 FILLER_0_9_105 ();
 sg13g2_decap_8 FILLER_0_9_112 ();
 sg13g2_decap_8 FILLER_0_9_119 ();
 sg13g2_decap_8 FILLER_0_9_126 ();
 sg13g2_decap_8 FILLER_0_9_133 ();
 sg13g2_decap_8 FILLER_0_9_140 ();
 sg13g2_decap_8 FILLER_0_9_147 ();
 sg13g2_decap_8 FILLER_0_9_154 ();
 sg13g2_decap_8 FILLER_0_9_161 ();
 sg13g2_decap_8 FILLER_0_9_168 ();
 sg13g2_decap_8 FILLER_0_9_175 ();
 sg13g2_decap_8 FILLER_0_9_182 ();
 sg13g2_decap_8 FILLER_0_9_189 ();
 sg13g2_decap_8 FILLER_0_9_196 ();
 sg13g2_decap_8 FILLER_0_9_203 ();
 sg13g2_decap_8 FILLER_0_9_210 ();
 sg13g2_decap_8 FILLER_0_9_217 ();
 sg13g2_decap_8 FILLER_0_9_224 ();
 sg13g2_decap_8 FILLER_0_9_231 ();
 sg13g2_decap_8 FILLER_0_9_238 ();
 sg13g2_decap_8 FILLER_0_9_245 ();
 sg13g2_decap_8 FILLER_0_9_252 ();
 sg13g2_decap_8 FILLER_0_9_259 ();
 sg13g2_decap_8 FILLER_0_9_266 ();
 sg13g2_decap_8 FILLER_0_9_273 ();
 sg13g2_decap_8 FILLER_0_9_280 ();
 sg13g2_decap_8 FILLER_0_9_287 ();
 sg13g2_decap_8 FILLER_0_9_294 ();
 sg13g2_decap_8 FILLER_0_9_301 ();
 sg13g2_decap_8 FILLER_0_9_308 ();
 sg13g2_decap_8 FILLER_0_9_315 ();
 sg13g2_decap_8 FILLER_0_9_322 ();
 sg13g2_decap_8 FILLER_0_9_329 ();
 sg13g2_decap_8 FILLER_0_9_336 ();
 sg13g2_decap_8 FILLER_0_9_343 ();
 sg13g2_decap_8 FILLER_0_9_350 ();
 sg13g2_decap_8 FILLER_0_9_357 ();
 sg13g2_decap_8 FILLER_0_9_364 ();
 sg13g2_decap_8 FILLER_0_9_371 ();
 sg13g2_decap_8 FILLER_0_9_378 ();
 sg13g2_decap_8 FILLER_0_9_385 ();
 sg13g2_decap_8 FILLER_0_9_392 ();
 sg13g2_decap_8 FILLER_0_9_399 ();
 sg13g2_decap_8 FILLER_0_9_406 ();
 sg13g2_decap_8 FILLER_0_9_413 ();
 sg13g2_decap_8 FILLER_0_9_420 ();
 sg13g2_decap_8 FILLER_0_9_427 ();
 sg13g2_decap_8 FILLER_0_9_434 ();
 sg13g2_decap_8 FILLER_0_9_441 ();
 sg13g2_decap_8 FILLER_0_9_448 ();
 sg13g2_decap_8 FILLER_0_9_455 ();
 sg13g2_decap_8 FILLER_0_9_462 ();
 sg13g2_decap_8 FILLER_0_9_469 ();
 sg13g2_decap_8 FILLER_0_9_476 ();
 sg13g2_decap_8 FILLER_0_9_483 ();
 sg13g2_decap_8 FILLER_0_9_490 ();
 sg13g2_decap_8 FILLER_0_9_497 ();
 sg13g2_decap_8 FILLER_0_9_504 ();
 sg13g2_decap_8 FILLER_0_9_511 ();
 sg13g2_decap_8 FILLER_0_9_518 ();
 sg13g2_decap_8 FILLER_0_9_525 ();
 sg13g2_decap_8 FILLER_0_9_532 ();
 sg13g2_decap_8 FILLER_0_9_539 ();
 sg13g2_decap_8 FILLER_0_9_546 ();
 sg13g2_decap_8 FILLER_0_9_553 ();
 sg13g2_decap_8 FILLER_0_9_560 ();
 sg13g2_decap_8 FILLER_0_9_567 ();
 sg13g2_decap_8 FILLER_0_9_574 ();
 sg13g2_decap_8 FILLER_0_9_581 ();
 sg13g2_decap_8 FILLER_0_9_588 ();
 sg13g2_decap_8 FILLER_0_9_595 ();
 sg13g2_decap_8 FILLER_0_9_602 ();
 sg13g2_decap_8 FILLER_0_9_609 ();
 sg13g2_decap_8 FILLER_0_9_616 ();
 sg13g2_decap_8 FILLER_0_9_623 ();
 sg13g2_decap_8 FILLER_0_9_630 ();
 sg13g2_decap_8 FILLER_0_9_637 ();
 sg13g2_decap_8 FILLER_0_9_644 ();
 sg13g2_decap_8 FILLER_0_9_651 ();
 sg13g2_decap_8 FILLER_0_9_658 ();
 sg13g2_decap_8 FILLER_0_9_665 ();
 sg13g2_decap_8 FILLER_0_9_672 ();
 sg13g2_decap_8 FILLER_0_9_679 ();
 sg13g2_decap_8 FILLER_0_9_686 ();
 sg13g2_decap_8 FILLER_0_9_693 ();
 sg13g2_decap_8 FILLER_0_9_700 ();
 sg13g2_decap_8 FILLER_0_9_707 ();
 sg13g2_decap_8 FILLER_0_9_714 ();
 sg13g2_decap_8 FILLER_0_9_721 ();
 sg13g2_decap_8 FILLER_0_9_728 ();
 sg13g2_decap_8 FILLER_0_9_735 ();
 sg13g2_decap_8 FILLER_0_9_742 ();
 sg13g2_decap_8 FILLER_0_9_749 ();
 sg13g2_decap_8 FILLER_0_9_756 ();
 sg13g2_decap_8 FILLER_0_9_763 ();
 sg13g2_decap_8 FILLER_0_9_770 ();
 sg13g2_decap_8 FILLER_0_9_777 ();
 sg13g2_decap_8 FILLER_0_9_784 ();
 sg13g2_decap_8 FILLER_0_9_791 ();
 sg13g2_decap_8 FILLER_0_9_798 ();
 sg13g2_decap_8 FILLER_0_9_805 ();
 sg13g2_decap_8 FILLER_0_9_812 ();
 sg13g2_decap_8 FILLER_0_9_819 ();
 sg13g2_decap_8 FILLER_0_9_826 ();
 sg13g2_decap_8 FILLER_0_9_833 ();
 sg13g2_decap_8 FILLER_0_9_840 ();
 sg13g2_decap_8 FILLER_0_9_847 ();
 sg13g2_decap_8 FILLER_0_9_854 ();
 sg13g2_decap_8 FILLER_0_9_861 ();
 sg13g2_decap_8 FILLER_0_9_868 ();
 sg13g2_decap_8 FILLER_0_9_875 ();
 sg13g2_decap_8 FILLER_0_9_882 ();
 sg13g2_decap_8 FILLER_0_9_889 ();
 sg13g2_decap_8 FILLER_0_9_896 ();
 sg13g2_decap_8 FILLER_0_9_903 ();
 sg13g2_decap_8 FILLER_0_9_910 ();
 sg13g2_decap_8 FILLER_0_9_917 ();
 sg13g2_decap_8 FILLER_0_9_924 ();
 sg13g2_decap_8 FILLER_0_9_931 ();
 sg13g2_decap_8 FILLER_0_9_938 ();
 sg13g2_decap_8 FILLER_0_9_945 ();
 sg13g2_decap_8 FILLER_0_9_952 ();
 sg13g2_decap_8 FILLER_0_9_959 ();
 sg13g2_decap_8 FILLER_0_9_966 ();
 sg13g2_decap_8 FILLER_0_9_973 ();
 sg13g2_decap_8 FILLER_0_9_980 ();
 sg13g2_decap_8 FILLER_0_9_987 ();
 sg13g2_decap_8 FILLER_0_9_994 ();
 sg13g2_decap_8 FILLER_0_9_1001 ();
 sg13g2_decap_8 FILLER_0_9_1008 ();
 sg13g2_decap_8 FILLER_0_9_1015 ();
 sg13g2_decap_8 FILLER_0_9_1022 ();
 sg13g2_decap_8 FILLER_0_9_1029 ();
 sg13g2_decap_8 FILLER_0_9_1036 ();
 sg13g2_decap_8 FILLER_0_9_1043 ();
 sg13g2_decap_8 FILLER_0_9_1050 ();
 sg13g2_decap_8 FILLER_0_9_1057 ();
 sg13g2_decap_8 FILLER_0_9_1064 ();
 sg13g2_decap_8 FILLER_0_9_1071 ();
 sg13g2_decap_8 FILLER_0_9_1078 ();
 sg13g2_decap_8 FILLER_0_9_1085 ();
 sg13g2_decap_8 FILLER_0_9_1092 ();
 sg13g2_decap_8 FILLER_0_9_1099 ();
 sg13g2_decap_8 FILLER_0_9_1106 ();
 sg13g2_decap_8 FILLER_0_9_1113 ();
 sg13g2_decap_8 FILLER_0_9_1120 ();
 sg13g2_decap_8 FILLER_0_9_1127 ();
 sg13g2_decap_8 FILLER_0_9_1134 ();
 sg13g2_decap_8 FILLER_0_9_1141 ();
 sg13g2_decap_8 FILLER_0_9_1148 ();
 sg13g2_decap_8 FILLER_0_9_1155 ();
 sg13g2_decap_8 FILLER_0_9_1162 ();
 sg13g2_decap_8 FILLER_0_9_1169 ();
 sg13g2_decap_8 FILLER_0_9_1176 ();
 sg13g2_decap_8 FILLER_0_9_1183 ();
 sg13g2_decap_8 FILLER_0_9_1190 ();
 sg13g2_decap_8 FILLER_0_9_1197 ();
 sg13g2_decap_8 FILLER_0_9_1204 ();
 sg13g2_decap_8 FILLER_0_9_1211 ();
 sg13g2_decap_8 FILLER_0_9_1218 ();
 sg13g2_fill_2 FILLER_0_9_1225 ();
 sg13g2_fill_1 FILLER_0_9_1227 ();
 sg13g2_decap_8 FILLER_0_10_0 ();
 sg13g2_decap_8 FILLER_0_10_7 ();
 sg13g2_decap_8 FILLER_0_10_14 ();
 sg13g2_decap_8 FILLER_0_10_21 ();
 sg13g2_decap_8 FILLER_0_10_28 ();
 sg13g2_decap_8 FILLER_0_10_35 ();
 sg13g2_decap_8 FILLER_0_10_42 ();
 sg13g2_decap_8 FILLER_0_10_49 ();
 sg13g2_decap_8 FILLER_0_10_56 ();
 sg13g2_decap_8 FILLER_0_10_63 ();
 sg13g2_decap_8 FILLER_0_10_70 ();
 sg13g2_decap_8 FILLER_0_10_77 ();
 sg13g2_decap_8 FILLER_0_10_84 ();
 sg13g2_decap_8 FILLER_0_10_91 ();
 sg13g2_decap_8 FILLER_0_10_98 ();
 sg13g2_decap_8 FILLER_0_10_105 ();
 sg13g2_decap_8 FILLER_0_10_112 ();
 sg13g2_decap_8 FILLER_0_10_119 ();
 sg13g2_decap_8 FILLER_0_10_126 ();
 sg13g2_decap_8 FILLER_0_10_133 ();
 sg13g2_decap_8 FILLER_0_10_140 ();
 sg13g2_decap_8 FILLER_0_10_147 ();
 sg13g2_decap_8 FILLER_0_10_154 ();
 sg13g2_decap_8 FILLER_0_10_161 ();
 sg13g2_decap_8 FILLER_0_10_168 ();
 sg13g2_decap_8 FILLER_0_10_175 ();
 sg13g2_decap_8 FILLER_0_10_182 ();
 sg13g2_decap_8 FILLER_0_10_189 ();
 sg13g2_decap_8 FILLER_0_10_196 ();
 sg13g2_decap_8 FILLER_0_10_203 ();
 sg13g2_decap_8 FILLER_0_10_210 ();
 sg13g2_decap_8 FILLER_0_10_217 ();
 sg13g2_decap_8 FILLER_0_10_224 ();
 sg13g2_decap_8 FILLER_0_10_231 ();
 sg13g2_decap_8 FILLER_0_10_238 ();
 sg13g2_decap_8 FILLER_0_10_245 ();
 sg13g2_decap_8 FILLER_0_10_252 ();
 sg13g2_decap_8 FILLER_0_10_259 ();
 sg13g2_decap_8 FILLER_0_10_266 ();
 sg13g2_decap_8 FILLER_0_10_273 ();
 sg13g2_decap_8 FILLER_0_10_280 ();
 sg13g2_decap_8 FILLER_0_10_287 ();
 sg13g2_decap_8 FILLER_0_10_294 ();
 sg13g2_decap_8 FILLER_0_10_301 ();
 sg13g2_decap_8 FILLER_0_10_308 ();
 sg13g2_decap_8 FILLER_0_10_315 ();
 sg13g2_decap_8 FILLER_0_10_322 ();
 sg13g2_decap_8 FILLER_0_10_329 ();
 sg13g2_decap_8 FILLER_0_10_336 ();
 sg13g2_decap_8 FILLER_0_10_343 ();
 sg13g2_decap_8 FILLER_0_10_350 ();
 sg13g2_decap_8 FILLER_0_10_357 ();
 sg13g2_decap_8 FILLER_0_10_364 ();
 sg13g2_decap_8 FILLER_0_10_371 ();
 sg13g2_decap_8 FILLER_0_10_378 ();
 sg13g2_decap_8 FILLER_0_10_385 ();
 sg13g2_decap_8 FILLER_0_10_392 ();
 sg13g2_decap_8 FILLER_0_10_399 ();
 sg13g2_decap_8 FILLER_0_10_406 ();
 sg13g2_decap_8 FILLER_0_10_413 ();
 sg13g2_decap_8 FILLER_0_10_420 ();
 sg13g2_decap_8 FILLER_0_10_427 ();
 sg13g2_decap_8 FILLER_0_10_434 ();
 sg13g2_decap_8 FILLER_0_10_441 ();
 sg13g2_decap_8 FILLER_0_10_448 ();
 sg13g2_decap_8 FILLER_0_10_455 ();
 sg13g2_decap_8 FILLER_0_10_462 ();
 sg13g2_decap_8 FILLER_0_10_469 ();
 sg13g2_decap_8 FILLER_0_10_476 ();
 sg13g2_decap_8 FILLER_0_10_483 ();
 sg13g2_decap_8 FILLER_0_10_490 ();
 sg13g2_decap_8 FILLER_0_10_497 ();
 sg13g2_decap_8 FILLER_0_10_504 ();
 sg13g2_decap_8 FILLER_0_10_511 ();
 sg13g2_decap_8 FILLER_0_10_518 ();
 sg13g2_decap_8 FILLER_0_10_525 ();
 sg13g2_decap_8 FILLER_0_10_532 ();
 sg13g2_decap_8 FILLER_0_10_539 ();
 sg13g2_decap_8 FILLER_0_10_546 ();
 sg13g2_decap_8 FILLER_0_10_553 ();
 sg13g2_decap_8 FILLER_0_10_560 ();
 sg13g2_decap_8 FILLER_0_10_567 ();
 sg13g2_decap_8 FILLER_0_10_574 ();
 sg13g2_decap_8 FILLER_0_10_581 ();
 sg13g2_decap_8 FILLER_0_10_588 ();
 sg13g2_decap_8 FILLER_0_10_595 ();
 sg13g2_decap_8 FILLER_0_10_602 ();
 sg13g2_decap_8 FILLER_0_10_609 ();
 sg13g2_decap_8 FILLER_0_10_616 ();
 sg13g2_decap_8 FILLER_0_10_623 ();
 sg13g2_decap_8 FILLER_0_10_630 ();
 sg13g2_decap_8 FILLER_0_10_637 ();
 sg13g2_decap_8 FILLER_0_10_644 ();
 sg13g2_decap_8 FILLER_0_10_651 ();
 sg13g2_decap_8 FILLER_0_10_658 ();
 sg13g2_decap_8 FILLER_0_10_665 ();
 sg13g2_decap_8 FILLER_0_10_672 ();
 sg13g2_decap_8 FILLER_0_10_679 ();
 sg13g2_decap_8 FILLER_0_10_686 ();
 sg13g2_decap_8 FILLER_0_10_693 ();
 sg13g2_decap_8 FILLER_0_10_700 ();
 sg13g2_decap_8 FILLER_0_10_707 ();
 sg13g2_decap_8 FILLER_0_10_714 ();
 sg13g2_decap_8 FILLER_0_10_721 ();
 sg13g2_decap_8 FILLER_0_10_728 ();
 sg13g2_decap_8 FILLER_0_10_735 ();
 sg13g2_decap_8 FILLER_0_10_742 ();
 sg13g2_decap_8 FILLER_0_10_749 ();
 sg13g2_decap_8 FILLER_0_10_756 ();
 sg13g2_decap_8 FILLER_0_10_763 ();
 sg13g2_decap_8 FILLER_0_10_770 ();
 sg13g2_decap_8 FILLER_0_10_777 ();
 sg13g2_decap_8 FILLER_0_10_784 ();
 sg13g2_decap_8 FILLER_0_10_791 ();
 sg13g2_decap_8 FILLER_0_10_798 ();
 sg13g2_decap_8 FILLER_0_10_805 ();
 sg13g2_decap_8 FILLER_0_10_812 ();
 sg13g2_decap_8 FILLER_0_10_819 ();
 sg13g2_decap_8 FILLER_0_10_826 ();
 sg13g2_decap_8 FILLER_0_10_833 ();
 sg13g2_decap_8 FILLER_0_10_840 ();
 sg13g2_decap_8 FILLER_0_10_847 ();
 sg13g2_decap_8 FILLER_0_10_854 ();
 sg13g2_decap_8 FILLER_0_10_861 ();
 sg13g2_decap_8 FILLER_0_10_868 ();
 sg13g2_decap_8 FILLER_0_10_875 ();
 sg13g2_decap_8 FILLER_0_10_882 ();
 sg13g2_decap_8 FILLER_0_10_889 ();
 sg13g2_decap_8 FILLER_0_10_896 ();
 sg13g2_decap_8 FILLER_0_10_903 ();
 sg13g2_decap_8 FILLER_0_10_910 ();
 sg13g2_decap_8 FILLER_0_10_917 ();
 sg13g2_decap_8 FILLER_0_10_924 ();
 sg13g2_decap_8 FILLER_0_10_931 ();
 sg13g2_decap_8 FILLER_0_10_938 ();
 sg13g2_decap_8 FILLER_0_10_945 ();
 sg13g2_decap_8 FILLER_0_10_952 ();
 sg13g2_decap_8 FILLER_0_10_959 ();
 sg13g2_decap_8 FILLER_0_10_966 ();
 sg13g2_decap_8 FILLER_0_10_973 ();
 sg13g2_decap_8 FILLER_0_10_980 ();
 sg13g2_decap_8 FILLER_0_10_987 ();
 sg13g2_decap_8 FILLER_0_10_994 ();
 sg13g2_decap_8 FILLER_0_10_1001 ();
 sg13g2_decap_8 FILLER_0_10_1008 ();
 sg13g2_decap_8 FILLER_0_10_1015 ();
 sg13g2_decap_8 FILLER_0_10_1022 ();
 sg13g2_decap_8 FILLER_0_10_1029 ();
 sg13g2_decap_8 FILLER_0_10_1036 ();
 sg13g2_decap_8 FILLER_0_10_1043 ();
 sg13g2_decap_8 FILLER_0_10_1050 ();
 sg13g2_decap_8 FILLER_0_10_1057 ();
 sg13g2_decap_8 FILLER_0_10_1064 ();
 sg13g2_decap_8 FILLER_0_10_1071 ();
 sg13g2_decap_8 FILLER_0_10_1078 ();
 sg13g2_decap_8 FILLER_0_10_1085 ();
 sg13g2_decap_8 FILLER_0_10_1092 ();
 sg13g2_decap_8 FILLER_0_10_1099 ();
 sg13g2_decap_8 FILLER_0_10_1106 ();
 sg13g2_decap_8 FILLER_0_10_1113 ();
 sg13g2_decap_8 FILLER_0_10_1120 ();
 sg13g2_decap_8 FILLER_0_10_1127 ();
 sg13g2_decap_8 FILLER_0_10_1134 ();
 sg13g2_decap_8 FILLER_0_10_1141 ();
 sg13g2_decap_8 FILLER_0_10_1148 ();
 sg13g2_decap_8 FILLER_0_10_1155 ();
 sg13g2_decap_8 FILLER_0_10_1162 ();
 sg13g2_decap_8 FILLER_0_10_1169 ();
 sg13g2_decap_8 FILLER_0_10_1176 ();
 sg13g2_decap_8 FILLER_0_10_1183 ();
 sg13g2_decap_8 FILLER_0_10_1190 ();
 sg13g2_decap_8 FILLER_0_10_1197 ();
 sg13g2_decap_8 FILLER_0_10_1204 ();
 sg13g2_decap_8 FILLER_0_10_1211 ();
 sg13g2_decap_8 FILLER_0_10_1218 ();
 sg13g2_fill_2 FILLER_0_10_1225 ();
 sg13g2_fill_1 FILLER_0_10_1227 ();
 sg13g2_decap_8 FILLER_0_11_0 ();
 sg13g2_decap_8 FILLER_0_11_7 ();
 sg13g2_decap_8 FILLER_0_11_14 ();
 sg13g2_decap_8 FILLER_0_11_21 ();
 sg13g2_decap_8 FILLER_0_11_28 ();
 sg13g2_decap_8 FILLER_0_11_35 ();
 sg13g2_decap_8 FILLER_0_11_42 ();
 sg13g2_decap_8 FILLER_0_11_49 ();
 sg13g2_decap_8 FILLER_0_11_56 ();
 sg13g2_decap_8 FILLER_0_11_63 ();
 sg13g2_decap_8 FILLER_0_11_70 ();
 sg13g2_decap_8 FILLER_0_11_77 ();
 sg13g2_decap_8 FILLER_0_11_84 ();
 sg13g2_decap_8 FILLER_0_11_91 ();
 sg13g2_decap_8 FILLER_0_11_98 ();
 sg13g2_decap_8 FILLER_0_11_105 ();
 sg13g2_decap_8 FILLER_0_11_112 ();
 sg13g2_decap_8 FILLER_0_11_119 ();
 sg13g2_decap_8 FILLER_0_11_126 ();
 sg13g2_decap_8 FILLER_0_11_133 ();
 sg13g2_decap_8 FILLER_0_11_140 ();
 sg13g2_decap_8 FILLER_0_11_147 ();
 sg13g2_decap_8 FILLER_0_11_154 ();
 sg13g2_decap_8 FILLER_0_11_161 ();
 sg13g2_decap_8 FILLER_0_11_168 ();
 sg13g2_decap_8 FILLER_0_11_175 ();
 sg13g2_decap_8 FILLER_0_11_182 ();
 sg13g2_decap_8 FILLER_0_11_189 ();
 sg13g2_decap_8 FILLER_0_11_196 ();
 sg13g2_decap_8 FILLER_0_11_203 ();
 sg13g2_decap_8 FILLER_0_11_210 ();
 sg13g2_decap_8 FILLER_0_11_217 ();
 sg13g2_decap_8 FILLER_0_11_224 ();
 sg13g2_decap_8 FILLER_0_11_231 ();
 sg13g2_decap_8 FILLER_0_11_238 ();
 sg13g2_decap_8 FILLER_0_11_245 ();
 sg13g2_decap_8 FILLER_0_11_252 ();
 sg13g2_decap_8 FILLER_0_11_259 ();
 sg13g2_decap_8 FILLER_0_11_266 ();
 sg13g2_decap_8 FILLER_0_11_273 ();
 sg13g2_decap_8 FILLER_0_11_280 ();
 sg13g2_decap_8 FILLER_0_11_287 ();
 sg13g2_decap_8 FILLER_0_11_294 ();
 sg13g2_decap_8 FILLER_0_11_301 ();
 sg13g2_decap_8 FILLER_0_11_308 ();
 sg13g2_decap_8 FILLER_0_11_315 ();
 sg13g2_decap_8 FILLER_0_11_322 ();
 sg13g2_decap_8 FILLER_0_11_329 ();
 sg13g2_decap_8 FILLER_0_11_336 ();
 sg13g2_decap_8 FILLER_0_11_343 ();
 sg13g2_decap_8 FILLER_0_11_350 ();
 sg13g2_decap_8 FILLER_0_11_357 ();
 sg13g2_decap_8 FILLER_0_11_364 ();
 sg13g2_decap_8 FILLER_0_11_371 ();
 sg13g2_decap_8 FILLER_0_11_378 ();
 sg13g2_decap_8 FILLER_0_11_385 ();
 sg13g2_decap_8 FILLER_0_11_392 ();
 sg13g2_decap_8 FILLER_0_11_399 ();
 sg13g2_decap_8 FILLER_0_11_406 ();
 sg13g2_decap_8 FILLER_0_11_413 ();
 sg13g2_decap_8 FILLER_0_11_420 ();
 sg13g2_decap_8 FILLER_0_11_427 ();
 sg13g2_decap_8 FILLER_0_11_434 ();
 sg13g2_decap_8 FILLER_0_11_441 ();
 sg13g2_decap_8 FILLER_0_11_448 ();
 sg13g2_decap_8 FILLER_0_11_455 ();
 sg13g2_decap_8 FILLER_0_11_462 ();
 sg13g2_decap_8 FILLER_0_11_469 ();
 sg13g2_decap_8 FILLER_0_11_476 ();
 sg13g2_decap_8 FILLER_0_11_483 ();
 sg13g2_decap_8 FILLER_0_11_490 ();
 sg13g2_decap_8 FILLER_0_11_497 ();
 sg13g2_decap_8 FILLER_0_11_504 ();
 sg13g2_decap_8 FILLER_0_11_511 ();
 sg13g2_decap_8 FILLER_0_11_518 ();
 sg13g2_decap_8 FILLER_0_11_525 ();
 sg13g2_decap_8 FILLER_0_11_532 ();
 sg13g2_decap_8 FILLER_0_11_539 ();
 sg13g2_decap_8 FILLER_0_11_546 ();
 sg13g2_decap_8 FILLER_0_11_553 ();
 sg13g2_decap_8 FILLER_0_11_560 ();
 sg13g2_decap_8 FILLER_0_11_567 ();
 sg13g2_decap_8 FILLER_0_11_574 ();
 sg13g2_decap_8 FILLER_0_11_581 ();
 sg13g2_decap_8 FILLER_0_11_588 ();
 sg13g2_decap_8 FILLER_0_11_595 ();
 sg13g2_decap_8 FILLER_0_11_602 ();
 sg13g2_decap_8 FILLER_0_11_609 ();
 sg13g2_decap_8 FILLER_0_11_616 ();
 sg13g2_decap_8 FILLER_0_11_623 ();
 sg13g2_decap_8 FILLER_0_11_630 ();
 sg13g2_decap_8 FILLER_0_11_637 ();
 sg13g2_decap_8 FILLER_0_11_644 ();
 sg13g2_decap_8 FILLER_0_11_651 ();
 sg13g2_decap_8 FILLER_0_11_658 ();
 sg13g2_decap_8 FILLER_0_11_665 ();
 sg13g2_decap_8 FILLER_0_11_672 ();
 sg13g2_decap_8 FILLER_0_11_679 ();
 sg13g2_decap_8 FILLER_0_11_686 ();
 sg13g2_decap_8 FILLER_0_11_693 ();
 sg13g2_decap_8 FILLER_0_11_700 ();
 sg13g2_decap_8 FILLER_0_11_707 ();
 sg13g2_decap_8 FILLER_0_11_714 ();
 sg13g2_decap_8 FILLER_0_11_721 ();
 sg13g2_decap_8 FILLER_0_11_728 ();
 sg13g2_decap_8 FILLER_0_11_735 ();
 sg13g2_decap_8 FILLER_0_11_742 ();
 sg13g2_decap_8 FILLER_0_11_749 ();
 sg13g2_decap_8 FILLER_0_11_756 ();
 sg13g2_decap_8 FILLER_0_11_763 ();
 sg13g2_decap_8 FILLER_0_11_770 ();
 sg13g2_decap_8 FILLER_0_11_777 ();
 sg13g2_decap_8 FILLER_0_11_784 ();
 sg13g2_decap_8 FILLER_0_11_791 ();
 sg13g2_decap_8 FILLER_0_11_798 ();
 sg13g2_decap_8 FILLER_0_11_805 ();
 sg13g2_decap_8 FILLER_0_11_812 ();
 sg13g2_decap_8 FILLER_0_11_819 ();
 sg13g2_decap_8 FILLER_0_11_826 ();
 sg13g2_decap_8 FILLER_0_11_833 ();
 sg13g2_decap_8 FILLER_0_11_840 ();
 sg13g2_decap_8 FILLER_0_11_847 ();
 sg13g2_decap_8 FILLER_0_11_854 ();
 sg13g2_decap_8 FILLER_0_11_861 ();
 sg13g2_decap_8 FILLER_0_11_868 ();
 sg13g2_decap_8 FILLER_0_11_875 ();
 sg13g2_decap_8 FILLER_0_11_882 ();
 sg13g2_decap_8 FILLER_0_11_889 ();
 sg13g2_decap_8 FILLER_0_11_896 ();
 sg13g2_decap_8 FILLER_0_11_903 ();
 sg13g2_decap_8 FILLER_0_11_910 ();
 sg13g2_decap_8 FILLER_0_11_917 ();
 sg13g2_decap_8 FILLER_0_11_924 ();
 sg13g2_decap_8 FILLER_0_11_931 ();
 sg13g2_decap_8 FILLER_0_11_938 ();
 sg13g2_decap_8 FILLER_0_11_945 ();
 sg13g2_decap_8 FILLER_0_11_952 ();
 sg13g2_decap_8 FILLER_0_11_959 ();
 sg13g2_decap_8 FILLER_0_11_966 ();
 sg13g2_decap_8 FILLER_0_11_973 ();
 sg13g2_decap_8 FILLER_0_11_980 ();
 sg13g2_decap_8 FILLER_0_11_987 ();
 sg13g2_decap_8 FILLER_0_11_994 ();
 sg13g2_decap_8 FILLER_0_11_1001 ();
 sg13g2_decap_8 FILLER_0_11_1008 ();
 sg13g2_decap_8 FILLER_0_11_1015 ();
 sg13g2_decap_8 FILLER_0_11_1022 ();
 sg13g2_decap_8 FILLER_0_11_1029 ();
 sg13g2_decap_8 FILLER_0_11_1036 ();
 sg13g2_decap_8 FILLER_0_11_1043 ();
 sg13g2_decap_8 FILLER_0_11_1050 ();
 sg13g2_decap_8 FILLER_0_11_1057 ();
 sg13g2_decap_8 FILLER_0_11_1064 ();
 sg13g2_decap_8 FILLER_0_11_1071 ();
 sg13g2_decap_8 FILLER_0_11_1078 ();
 sg13g2_decap_8 FILLER_0_11_1085 ();
 sg13g2_decap_8 FILLER_0_11_1092 ();
 sg13g2_decap_8 FILLER_0_11_1099 ();
 sg13g2_decap_8 FILLER_0_11_1106 ();
 sg13g2_decap_8 FILLER_0_11_1113 ();
 sg13g2_decap_8 FILLER_0_11_1120 ();
 sg13g2_decap_8 FILLER_0_11_1127 ();
 sg13g2_decap_8 FILLER_0_11_1134 ();
 sg13g2_decap_8 FILLER_0_11_1141 ();
 sg13g2_decap_8 FILLER_0_11_1148 ();
 sg13g2_decap_8 FILLER_0_11_1155 ();
 sg13g2_decap_8 FILLER_0_11_1162 ();
 sg13g2_decap_8 FILLER_0_11_1169 ();
 sg13g2_decap_8 FILLER_0_11_1176 ();
 sg13g2_decap_8 FILLER_0_11_1183 ();
 sg13g2_decap_8 FILLER_0_11_1190 ();
 sg13g2_decap_8 FILLER_0_11_1197 ();
 sg13g2_decap_8 FILLER_0_11_1204 ();
 sg13g2_decap_8 FILLER_0_11_1211 ();
 sg13g2_decap_8 FILLER_0_11_1218 ();
 sg13g2_fill_2 FILLER_0_11_1225 ();
 sg13g2_fill_1 FILLER_0_11_1227 ();
 sg13g2_decap_8 FILLER_0_12_0 ();
 sg13g2_decap_8 FILLER_0_12_7 ();
 sg13g2_decap_8 FILLER_0_12_14 ();
 sg13g2_decap_8 FILLER_0_12_21 ();
 sg13g2_decap_8 FILLER_0_12_28 ();
 sg13g2_decap_8 FILLER_0_12_35 ();
 sg13g2_decap_8 FILLER_0_12_42 ();
 sg13g2_decap_8 FILLER_0_12_49 ();
 sg13g2_decap_8 FILLER_0_12_56 ();
 sg13g2_decap_8 FILLER_0_12_63 ();
 sg13g2_decap_8 FILLER_0_12_70 ();
 sg13g2_decap_8 FILLER_0_12_77 ();
 sg13g2_decap_8 FILLER_0_12_84 ();
 sg13g2_decap_8 FILLER_0_12_91 ();
 sg13g2_decap_8 FILLER_0_12_98 ();
 sg13g2_decap_8 FILLER_0_12_105 ();
 sg13g2_decap_8 FILLER_0_12_112 ();
 sg13g2_decap_8 FILLER_0_12_119 ();
 sg13g2_decap_8 FILLER_0_12_126 ();
 sg13g2_decap_8 FILLER_0_12_133 ();
 sg13g2_decap_8 FILLER_0_12_140 ();
 sg13g2_decap_8 FILLER_0_12_147 ();
 sg13g2_decap_8 FILLER_0_12_154 ();
 sg13g2_decap_8 FILLER_0_12_161 ();
 sg13g2_decap_8 FILLER_0_12_168 ();
 sg13g2_decap_8 FILLER_0_12_175 ();
 sg13g2_decap_8 FILLER_0_12_182 ();
 sg13g2_decap_8 FILLER_0_12_189 ();
 sg13g2_decap_8 FILLER_0_12_196 ();
 sg13g2_decap_8 FILLER_0_12_203 ();
 sg13g2_decap_8 FILLER_0_12_210 ();
 sg13g2_decap_8 FILLER_0_12_217 ();
 sg13g2_decap_8 FILLER_0_12_224 ();
 sg13g2_decap_8 FILLER_0_12_231 ();
 sg13g2_decap_8 FILLER_0_12_238 ();
 sg13g2_decap_8 FILLER_0_12_245 ();
 sg13g2_decap_8 FILLER_0_12_252 ();
 sg13g2_decap_8 FILLER_0_12_259 ();
 sg13g2_decap_8 FILLER_0_12_266 ();
 sg13g2_decap_8 FILLER_0_12_273 ();
 sg13g2_decap_8 FILLER_0_12_280 ();
 sg13g2_decap_8 FILLER_0_12_287 ();
 sg13g2_decap_8 FILLER_0_12_294 ();
 sg13g2_decap_8 FILLER_0_12_301 ();
 sg13g2_decap_8 FILLER_0_12_308 ();
 sg13g2_decap_8 FILLER_0_12_315 ();
 sg13g2_decap_8 FILLER_0_12_322 ();
 sg13g2_decap_8 FILLER_0_12_329 ();
 sg13g2_decap_8 FILLER_0_12_336 ();
 sg13g2_decap_8 FILLER_0_12_343 ();
 sg13g2_decap_8 FILLER_0_12_350 ();
 sg13g2_decap_8 FILLER_0_12_357 ();
 sg13g2_decap_8 FILLER_0_12_364 ();
 sg13g2_decap_8 FILLER_0_12_371 ();
 sg13g2_decap_8 FILLER_0_12_378 ();
 sg13g2_decap_8 FILLER_0_12_385 ();
 sg13g2_decap_8 FILLER_0_12_392 ();
 sg13g2_decap_8 FILLER_0_12_399 ();
 sg13g2_decap_8 FILLER_0_12_406 ();
 sg13g2_decap_8 FILLER_0_12_413 ();
 sg13g2_decap_8 FILLER_0_12_420 ();
 sg13g2_decap_8 FILLER_0_12_427 ();
 sg13g2_decap_8 FILLER_0_12_434 ();
 sg13g2_decap_8 FILLER_0_12_441 ();
 sg13g2_decap_8 FILLER_0_12_448 ();
 sg13g2_decap_8 FILLER_0_12_455 ();
 sg13g2_decap_8 FILLER_0_12_462 ();
 sg13g2_decap_8 FILLER_0_12_469 ();
 sg13g2_decap_8 FILLER_0_12_476 ();
 sg13g2_decap_8 FILLER_0_12_483 ();
 sg13g2_decap_8 FILLER_0_12_490 ();
 sg13g2_decap_8 FILLER_0_12_497 ();
 sg13g2_decap_8 FILLER_0_12_504 ();
 sg13g2_decap_8 FILLER_0_12_511 ();
 sg13g2_decap_8 FILLER_0_12_518 ();
 sg13g2_decap_8 FILLER_0_12_525 ();
 sg13g2_decap_8 FILLER_0_12_532 ();
 sg13g2_decap_8 FILLER_0_12_539 ();
 sg13g2_decap_8 FILLER_0_12_546 ();
 sg13g2_decap_8 FILLER_0_12_553 ();
 sg13g2_decap_8 FILLER_0_12_560 ();
 sg13g2_decap_8 FILLER_0_12_567 ();
 sg13g2_decap_8 FILLER_0_12_574 ();
 sg13g2_decap_8 FILLER_0_12_581 ();
 sg13g2_decap_8 FILLER_0_12_588 ();
 sg13g2_decap_8 FILLER_0_12_595 ();
 sg13g2_decap_8 FILLER_0_12_602 ();
 sg13g2_decap_8 FILLER_0_12_609 ();
 sg13g2_decap_8 FILLER_0_12_616 ();
 sg13g2_decap_8 FILLER_0_12_623 ();
 sg13g2_decap_8 FILLER_0_12_630 ();
 sg13g2_decap_8 FILLER_0_12_637 ();
 sg13g2_decap_8 FILLER_0_12_644 ();
 sg13g2_decap_8 FILLER_0_12_651 ();
 sg13g2_decap_8 FILLER_0_12_658 ();
 sg13g2_decap_8 FILLER_0_12_665 ();
 sg13g2_decap_8 FILLER_0_12_672 ();
 sg13g2_decap_8 FILLER_0_12_679 ();
 sg13g2_decap_8 FILLER_0_12_686 ();
 sg13g2_decap_8 FILLER_0_12_693 ();
 sg13g2_decap_8 FILLER_0_12_700 ();
 sg13g2_decap_8 FILLER_0_12_707 ();
 sg13g2_decap_8 FILLER_0_12_714 ();
 sg13g2_decap_8 FILLER_0_12_721 ();
 sg13g2_decap_8 FILLER_0_12_728 ();
 sg13g2_decap_8 FILLER_0_12_735 ();
 sg13g2_decap_8 FILLER_0_12_742 ();
 sg13g2_decap_8 FILLER_0_12_749 ();
 sg13g2_decap_8 FILLER_0_12_756 ();
 sg13g2_decap_8 FILLER_0_12_763 ();
 sg13g2_decap_8 FILLER_0_12_770 ();
 sg13g2_decap_8 FILLER_0_12_777 ();
 sg13g2_decap_8 FILLER_0_12_784 ();
 sg13g2_decap_8 FILLER_0_12_791 ();
 sg13g2_decap_8 FILLER_0_12_798 ();
 sg13g2_decap_8 FILLER_0_12_805 ();
 sg13g2_decap_8 FILLER_0_12_812 ();
 sg13g2_decap_8 FILLER_0_12_819 ();
 sg13g2_decap_8 FILLER_0_12_826 ();
 sg13g2_decap_8 FILLER_0_12_833 ();
 sg13g2_decap_8 FILLER_0_12_840 ();
 sg13g2_decap_8 FILLER_0_12_847 ();
 sg13g2_decap_8 FILLER_0_12_854 ();
 sg13g2_decap_8 FILLER_0_12_861 ();
 sg13g2_decap_8 FILLER_0_12_868 ();
 sg13g2_decap_8 FILLER_0_12_875 ();
 sg13g2_decap_8 FILLER_0_12_882 ();
 sg13g2_decap_8 FILLER_0_12_889 ();
 sg13g2_decap_8 FILLER_0_12_896 ();
 sg13g2_decap_8 FILLER_0_12_903 ();
 sg13g2_decap_8 FILLER_0_12_910 ();
 sg13g2_decap_8 FILLER_0_12_917 ();
 sg13g2_decap_8 FILLER_0_12_924 ();
 sg13g2_decap_8 FILLER_0_12_931 ();
 sg13g2_decap_8 FILLER_0_12_938 ();
 sg13g2_decap_8 FILLER_0_12_945 ();
 sg13g2_decap_8 FILLER_0_12_952 ();
 sg13g2_decap_8 FILLER_0_12_959 ();
 sg13g2_decap_8 FILLER_0_12_966 ();
 sg13g2_decap_8 FILLER_0_12_973 ();
 sg13g2_decap_8 FILLER_0_12_980 ();
 sg13g2_decap_8 FILLER_0_12_987 ();
 sg13g2_decap_8 FILLER_0_12_994 ();
 sg13g2_decap_8 FILLER_0_12_1001 ();
 sg13g2_decap_8 FILLER_0_12_1008 ();
 sg13g2_decap_8 FILLER_0_12_1015 ();
 sg13g2_decap_8 FILLER_0_12_1022 ();
 sg13g2_decap_8 FILLER_0_12_1029 ();
 sg13g2_decap_8 FILLER_0_12_1036 ();
 sg13g2_decap_8 FILLER_0_12_1043 ();
 sg13g2_decap_8 FILLER_0_12_1050 ();
 sg13g2_decap_8 FILLER_0_12_1057 ();
 sg13g2_decap_8 FILLER_0_12_1064 ();
 sg13g2_decap_8 FILLER_0_12_1071 ();
 sg13g2_decap_8 FILLER_0_12_1078 ();
 sg13g2_decap_8 FILLER_0_12_1085 ();
 sg13g2_decap_8 FILLER_0_12_1092 ();
 sg13g2_decap_8 FILLER_0_12_1099 ();
 sg13g2_decap_8 FILLER_0_12_1106 ();
 sg13g2_decap_8 FILLER_0_12_1113 ();
 sg13g2_decap_8 FILLER_0_12_1120 ();
 sg13g2_decap_8 FILLER_0_12_1127 ();
 sg13g2_decap_8 FILLER_0_12_1134 ();
 sg13g2_decap_8 FILLER_0_12_1141 ();
 sg13g2_decap_8 FILLER_0_12_1148 ();
 sg13g2_decap_8 FILLER_0_12_1155 ();
 sg13g2_decap_8 FILLER_0_12_1162 ();
 sg13g2_decap_8 FILLER_0_12_1169 ();
 sg13g2_decap_8 FILLER_0_12_1176 ();
 sg13g2_decap_8 FILLER_0_12_1183 ();
 sg13g2_decap_8 FILLER_0_12_1190 ();
 sg13g2_decap_8 FILLER_0_12_1197 ();
 sg13g2_decap_8 FILLER_0_12_1204 ();
 sg13g2_decap_8 FILLER_0_12_1211 ();
 sg13g2_decap_8 FILLER_0_12_1218 ();
 sg13g2_fill_2 FILLER_0_12_1225 ();
 sg13g2_fill_1 FILLER_0_12_1227 ();
 sg13g2_decap_8 FILLER_0_13_0 ();
 sg13g2_decap_8 FILLER_0_13_7 ();
 sg13g2_decap_8 FILLER_0_13_14 ();
 sg13g2_decap_8 FILLER_0_13_21 ();
 sg13g2_decap_8 FILLER_0_13_28 ();
 sg13g2_decap_8 FILLER_0_13_35 ();
 sg13g2_decap_8 FILLER_0_13_42 ();
 sg13g2_decap_8 FILLER_0_13_49 ();
 sg13g2_decap_8 FILLER_0_13_56 ();
 sg13g2_decap_8 FILLER_0_13_63 ();
 sg13g2_decap_8 FILLER_0_13_70 ();
 sg13g2_decap_8 FILLER_0_13_77 ();
 sg13g2_decap_8 FILLER_0_13_84 ();
 sg13g2_decap_8 FILLER_0_13_91 ();
 sg13g2_decap_8 FILLER_0_13_98 ();
 sg13g2_decap_8 FILLER_0_13_105 ();
 sg13g2_decap_8 FILLER_0_13_112 ();
 sg13g2_decap_8 FILLER_0_13_119 ();
 sg13g2_decap_8 FILLER_0_13_126 ();
 sg13g2_decap_8 FILLER_0_13_133 ();
 sg13g2_decap_8 FILLER_0_13_140 ();
 sg13g2_decap_8 FILLER_0_13_147 ();
 sg13g2_decap_8 FILLER_0_13_154 ();
 sg13g2_decap_8 FILLER_0_13_161 ();
 sg13g2_decap_8 FILLER_0_13_168 ();
 sg13g2_decap_8 FILLER_0_13_175 ();
 sg13g2_decap_8 FILLER_0_13_182 ();
 sg13g2_decap_8 FILLER_0_13_189 ();
 sg13g2_decap_8 FILLER_0_13_196 ();
 sg13g2_decap_8 FILLER_0_13_203 ();
 sg13g2_decap_8 FILLER_0_13_210 ();
 sg13g2_decap_8 FILLER_0_13_217 ();
 sg13g2_decap_8 FILLER_0_13_224 ();
 sg13g2_decap_8 FILLER_0_13_231 ();
 sg13g2_decap_8 FILLER_0_13_238 ();
 sg13g2_decap_8 FILLER_0_13_245 ();
 sg13g2_decap_8 FILLER_0_13_252 ();
 sg13g2_decap_8 FILLER_0_13_259 ();
 sg13g2_decap_8 FILLER_0_13_266 ();
 sg13g2_decap_8 FILLER_0_13_273 ();
 sg13g2_decap_8 FILLER_0_13_280 ();
 sg13g2_decap_8 FILLER_0_13_287 ();
 sg13g2_decap_8 FILLER_0_13_294 ();
 sg13g2_decap_8 FILLER_0_13_301 ();
 sg13g2_decap_8 FILLER_0_13_308 ();
 sg13g2_decap_8 FILLER_0_13_315 ();
 sg13g2_decap_8 FILLER_0_13_322 ();
 sg13g2_decap_8 FILLER_0_13_329 ();
 sg13g2_decap_8 FILLER_0_13_336 ();
 sg13g2_decap_8 FILLER_0_13_343 ();
 sg13g2_decap_8 FILLER_0_13_350 ();
 sg13g2_decap_8 FILLER_0_13_357 ();
 sg13g2_decap_8 FILLER_0_13_364 ();
 sg13g2_decap_8 FILLER_0_13_371 ();
 sg13g2_decap_8 FILLER_0_13_378 ();
 sg13g2_decap_8 FILLER_0_13_385 ();
 sg13g2_decap_8 FILLER_0_13_392 ();
 sg13g2_decap_8 FILLER_0_13_399 ();
 sg13g2_decap_8 FILLER_0_13_406 ();
 sg13g2_decap_8 FILLER_0_13_413 ();
 sg13g2_decap_8 FILLER_0_13_420 ();
 sg13g2_decap_8 FILLER_0_13_427 ();
 sg13g2_decap_8 FILLER_0_13_434 ();
 sg13g2_decap_8 FILLER_0_13_441 ();
 sg13g2_decap_8 FILLER_0_13_448 ();
 sg13g2_decap_8 FILLER_0_13_455 ();
 sg13g2_decap_8 FILLER_0_13_462 ();
 sg13g2_decap_8 FILLER_0_13_469 ();
 sg13g2_decap_8 FILLER_0_13_476 ();
 sg13g2_decap_8 FILLER_0_13_483 ();
 sg13g2_decap_8 FILLER_0_13_490 ();
 sg13g2_decap_8 FILLER_0_13_497 ();
 sg13g2_decap_8 FILLER_0_13_504 ();
 sg13g2_decap_8 FILLER_0_13_511 ();
 sg13g2_decap_8 FILLER_0_13_518 ();
 sg13g2_decap_8 FILLER_0_13_525 ();
 sg13g2_decap_8 FILLER_0_13_532 ();
 sg13g2_decap_8 FILLER_0_13_539 ();
 sg13g2_decap_8 FILLER_0_13_546 ();
 sg13g2_decap_8 FILLER_0_13_553 ();
 sg13g2_decap_8 FILLER_0_13_560 ();
 sg13g2_decap_8 FILLER_0_13_567 ();
 sg13g2_decap_8 FILLER_0_13_574 ();
 sg13g2_decap_8 FILLER_0_13_581 ();
 sg13g2_decap_8 FILLER_0_13_588 ();
 sg13g2_decap_8 FILLER_0_13_595 ();
 sg13g2_decap_8 FILLER_0_13_602 ();
 sg13g2_decap_8 FILLER_0_13_609 ();
 sg13g2_decap_8 FILLER_0_13_616 ();
 sg13g2_decap_8 FILLER_0_13_623 ();
 sg13g2_decap_8 FILLER_0_13_630 ();
 sg13g2_decap_8 FILLER_0_13_637 ();
 sg13g2_decap_8 FILLER_0_13_644 ();
 sg13g2_decap_8 FILLER_0_13_651 ();
 sg13g2_decap_8 FILLER_0_13_658 ();
 sg13g2_decap_8 FILLER_0_13_665 ();
 sg13g2_decap_8 FILLER_0_13_672 ();
 sg13g2_decap_8 FILLER_0_13_679 ();
 sg13g2_decap_8 FILLER_0_13_686 ();
 sg13g2_decap_8 FILLER_0_13_693 ();
 sg13g2_decap_8 FILLER_0_13_700 ();
 sg13g2_decap_8 FILLER_0_13_707 ();
 sg13g2_decap_8 FILLER_0_13_714 ();
 sg13g2_decap_8 FILLER_0_13_721 ();
 sg13g2_decap_8 FILLER_0_13_728 ();
 sg13g2_decap_8 FILLER_0_13_735 ();
 sg13g2_decap_8 FILLER_0_13_742 ();
 sg13g2_decap_8 FILLER_0_13_749 ();
 sg13g2_decap_8 FILLER_0_13_756 ();
 sg13g2_decap_8 FILLER_0_13_763 ();
 sg13g2_decap_8 FILLER_0_13_770 ();
 sg13g2_decap_8 FILLER_0_13_777 ();
 sg13g2_decap_8 FILLER_0_13_784 ();
 sg13g2_decap_8 FILLER_0_13_791 ();
 sg13g2_decap_8 FILLER_0_13_798 ();
 sg13g2_decap_8 FILLER_0_13_805 ();
 sg13g2_decap_8 FILLER_0_13_812 ();
 sg13g2_decap_8 FILLER_0_13_819 ();
 sg13g2_decap_8 FILLER_0_13_826 ();
 sg13g2_decap_8 FILLER_0_13_833 ();
 sg13g2_decap_8 FILLER_0_13_840 ();
 sg13g2_decap_8 FILLER_0_13_847 ();
 sg13g2_decap_8 FILLER_0_13_854 ();
 sg13g2_decap_8 FILLER_0_13_861 ();
 sg13g2_decap_8 FILLER_0_13_868 ();
 sg13g2_decap_8 FILLER_0_13_875 ();
 sg13g2_decap_8 FILLER_0_13_882 ();
 sg13g2_decap_8 FILLER_0_13_889 ();
 sg13g2_decap_8 FILLER_0_13_896 ();
 sg13g2_decap_8 FILLER_0_13_903 ();
 sg13g2_decap_8 FILLER_0_13_910 ();
 sg13g2_decap_8 FILLER_0_13_917 ();
 sg13g2_decap_8 FILLER_0_13_924 ();
 sg13g2_decap_8 FILLER_0_13_931 ();
 sg13g2_decap_8 FILLER_0_13_938 ();
 sg13g2_decap_8 FILLER_0_13_945 ();
 sg13g2_decap_8 FILLER_0_13_952 ();
 sg13g2_decap_8 FILLER_0_13_959 ();
 sg13g2_decap_8 FILLER_0_13_966 ();
 sg13g2_decap_8 FILLER_0_13_973 ();
 sg13g2_decap_8 FILLER_0_13_980 ();
 sg13g2_decap_8 FILLER_0_13_987 ();
 sg13g2_decap_8 FILLER_0_13_994 ();
 sg13g2_decap_8 FILLER_0_13_1001 ();
 sg13g2_decap_8 FILLER_0_13_1008 ();
 sg13g2_decap_8 FILLER_0_13_1015 ();
 sg13g2_decap_8 FILLER_0_13_1022 ();
 sg13g2_decap_8 FILLER_0_13_1029 ();
 sg13g2_decap_8 FILLER_0_13_1036 ();
 sg13g2_decap_8 FILLER_0_13_1043 ();
 sg13g2_decap_8 FILLER_0_13_1050 ();
 sg13g2_decap_8 FILLER_0_13_1057 ();
 sg13g2_decap_8 FILLER_0_13_1064 ();
 sg13g2_decap_8 FILLER_0_13_1071 ();
 sg13g2_decap_8 FILLER_0_13_1078 ();
 sg13g2_decap_8 FILLER_0_13_1085 ();
 sg13g2_decap_8 FILLER_0_13_1092 ();
 sg13g2_decap_8 FILLER_0_13_1099 ();
 sg13g2_decap_8 FILLER_0_13_1106 ();
 sg13g2_decap_8 FILLER_0_13_1113 ();
 sg13g2_decap_8 FILLER_0_13_1120 ();
 sg13g2_decap_8 FILLER_0_13_1127 ();
 sg13g2_decap_8 FILLER_0_13_1134 ();
 sg13g2_decap_8 FILLER_0_13_1141 ();
 sg13g2_decap_8 FILLER_0_13_1148 ();
 sg13g2_decap_8 FILLER_0_13_1155 ();
 sg13g2_decap_8 FILLER_0_13_1162 ();
 sg13g2_decap_8 FILLER_0_13_1169 ();
 sg13g2_decap_8 FILLER_0_13_1176 ();
 sg13g2_decap_8 FILLER_0_13_1183 ();
 sg13g2_decap_8 FILLER_0_13_1190 ();
 sg13g2_decap_8 FILLER_0_13_1197 ();
 sg13g2_decap_8 FILLER_0_13_1204 ();
 sg13g2_decap_8 FILLER_0_13_1211 ();
 sg13g2_decap_8 FILLER_0_13_1218 ();
 sg13g2_fill_2 FILLER_0_13_1225 ();
 sg13g2_fill_1 FILLER_0_13_1227 ();
 sg13g2_decap_8 FILLER_0_14_0 ();
 sg13g2_decap_8 FILLER_0_14_7 ();
 sg13g2_decap_8 FILLER_0_14_14 ();
 sg13g2_decap_8 FILLER_0_14_21 ();
 sg13g2_decap_8 FILLER_0_14_28 ();
 sg13g2_decap_8 FILLER_0_14_35 ();
 sg13g2_decap_8 FILLER_0_14_42 ();
 sg13g2_decap_8 FILLER_0_14_49 ();
 sg13g2_decap_8 FILLER_0_14_56 ();
 sg13g2_decap_8 FILLER_0_14_63 ();
 sg13g2_decap_8 FILLER_0_14_70 ();
 sg13g2_decap_8 FILLER_0_14_77 ();
 sg13g2_decap_8 FILLER_0_14_84 ();
 sg13g2_decap_8 FILLER_0_14_91 ();
 sg13g2_decap_8 FILLER_0_14_98 ();
 sg13g2_decap_8 FILLER_0_14_105 ();
 sg13g2_decap_8 FILLER_0_14_112 ();
 sg13g2_decap_8 FILLER_0_14_119 ();
 sg13g2_decap_8 FILLER_0_14_126 ();
 sg13g2_decap_8 FILLER_0_14_133 ();
 sg13g2_decap_8 FILLER_0_14_140 ();
 sg13g2_decap_8 FILLER_0_14_147 ();
 sg13g2_decap_8 FILLER_0_14_154 ();
 sg13g2_decap_8 FILLER_0_14_161 ();
 sg13g2_decap_8 FILLER_0_14_168 ();
 sg13g2_decap_8 FILLER_0_14_175 ();
 sg13g2_decap_8 FILLER_0_14_182 ();
 sg13g2_decap_8 FILLER_0_14_189 ();
 sg13g2_decap_8 FILLER_0_14_196 ();
 sg13g2_decap_8 FILLER_0_14_203 ();
 sg13g2_decap_8 FILLER_0_14_210 ();
 sg13g2_decap_8 FILLER_0_14_217 ();
 sg13g2_decap_8 FILLER_0_14_224 ();
 sg13g2_decap_8 FILLER_0_14_231 ();
 sg13g2_decap_8 FILLER_0_14_238 ();
 sg13g2_decap_8 FILLER_0_14_245 ();
 sg13g2_decap_8 FILLER_0_14_252 ();
 sg13g2_decap_8 FILLER_0_14_259 ();
 sg13g2_decap_8 FILLER_0_14_266 ();
 sg13g2_decap_8 FILLER_0_14_273 ();
 sg13g2_decap_8 FILLER_0_14_280 ();
 sg13g2_decap_8 FILLER_0_14_287 ();
 sg13g2_decap_8 FILLER_0_14_294 ();
 sg13g2_decap_8 FILLER_0_14_301 ();
 sg13g2_decap_8 FILLER_0_14_308 ();
 sg13g2_decap_8 FILLER_0_14_315 ();
 sg13g2_decap_8 FILLER_0_14_322 ();
 sg13g2_decap_8 FILLER_0_14_329 ();
 sg13g2_decap_8 FILLER_0_14_336 ();
 sg13g2_decap_8 FILLER_0_14_343 ();
 sg13g2_decap_8 FILLER_0_14_350 ();
 sg13g2_decap_8 FILLER_0_14_357 ();
 sg13g2_decap_8 FILLER_0_14_364 ();
 sg13g2_decap_8 FILLER_0_14_371 ();
 sg13g2_decap_8 FILLER_0_14_378 ();
 sg13g2_decap_8 FILLER_0_14_385 ();
 sg13g2_decap_8 FILLER_0_14_392 ();
 sg13g2_decap_8 FILLER_0_14_399 ();
 sg13g2_decap_8 FILLER_0_14_406 ();
 sg13g2_decap_8 FILLER_0_14_413 ();
 sg13g2_decap_8 FILLER_0_14_420 ();
 sg13g2_decap_8 FILLER_0_14_427 ();
 sg13g2_decap_8 FILLER_0_14_434 ();
 sg13g2_decap_8 FILLER_0_14_441 ();
 sg13g2_decap_8 FILLER_0_14_448 ();
 sg13g2_decap_8 FILLER_0_14_455 ();
 sg13g2_decap_8 FILLER_0_14_462 ();
 sg13g2_decap_8 FILLER_0_14_469 ();
 sg13g2_decap_8 FILLER_0_14_476 ();
 sg13g2_decap_8 FILLER_0_14_483 ();
 sg13g2_decap_8 FILLER_0_14_490 ();
 sg13g2_decap_8 FILLER_0_14_497 ();
 sg13g2_decap_8 FILLER_0_14_504 ();
 sg13g2_decap_8 FILLER_0_14_511 ();
 sg13g2_decap_8 FILLER_0_14_518 ();
 sg13g2_decap_8 FILLER_0_14_525 ();
 sg13g2_decap_8 FILLER_0_14_532 ();
 sg13g2_decap_8 FILLER_0_14_539 ();
 sg13g2_decap_8 FILLER_0_14_546 ();
 sg13g2_decap_8 FILLER_0_14_553 ();
 sg13g2_decap_8 FILLER_0_14_560 ();
 sg13g2_decap_8 FILLER_0_14_567 ();
 sg13g2_decap_8 FILLER_0_14_574 ();
 sg13g2_decap_8 FILLER_0_14_581 ();
 sg13g2_decap_8 FILLER_0_14_588 ();
 sg13g2_decap_8 FILLER_0_14_595 ();
 sg13g2_decap_8 FILLER_0_14_602 ();
 sg13g2_decap_8 FILLER_0_14_609 ();
 sg13g2_decap_8 FILLER_0_14_616 ();
 sg13g2_decap_8 FILLER_0_14_623 ();
 sg13g2_decap_8 FILLER_0_14_630 ();
 sg13g2_decap_8 FILLER_0_14_637 ();
 sg13g2_decap_8 FILLER_0_14_644 ();
 sg13g2_decap_8 FILLER_0_14_651 ();
 sg13g2_decap_8 FILLER_0_14_658 ();
 sg13g2_decap_8 FILLER_0_14_665 ();
 sg13g2_decap_8 FILLER_0_14_672 ();
 sg13g2_decap_8 FILLER_0_14_679 ();
 sg13g2_decap_8 FILLER_0_14_686 ();
 sg13g2_decap_8 FILLER_0_14_693 ();
 sg13g2_decap_8 FILLER_0_14_700 ();
 sg13g2_decap_8 FILLER_0_14_707 ();
 sg13g2_decap_8 FILLER_0_14_714 ();
 sg13g2_decap_8 FILLER_0_14_721 ();
 sg13g2_decap_8 FILLER_0_14_728 ();
 sg13g2_decap_8 FILLER_0_14_735 ();
 sg13g2_decap_8 FILLER_0_14_742 ();
 sg13g2_decap_8 FILLER_0_14_749 ();
 sg13g2_decap_8 FILLER_0_14_756 ();
 sg13g2_decap_8 FILLER_0_14_763 ();
 sg13g2_decap_8 FILLER_0_14_770 ();
 sg13g2_decap_8 FILLER_0_14_777 ();
 sg13g2_decap_8 FILLER_0_14_784 ();
 sg13g2_decap_8 FILLER_0_14_791 ();
 sg13g2_decap_8 FILLER_0_14_798 ();
 sg13g2_decap_8 FILLER_0_14_805 ();
 sg13g2_decap_8 FILLER_0_14_812 ();
 sg13g2_decap_8 FILLER_0_14_819 ();
 sg13g2_decap_8 FILLER_0_14_826 ();
 sg13g2_decap_8 FILLER_0_14_833 ();
 sg13g2_decap_8 FILLER_0_14_840 ();
 sg13g2_decap_8 FILLER_0_14_847 ();
 sg13g2_decap_8 FILLER_0_14_854 ();
 sg13g2_decap_8 FILLER_0_14_861 ();
 sg13g2_decap_8 FILLER_0_14_868 ();
 sg13g2_decap_8 FILLER_0_14_875 ();
 sg13g2_decap_8 FILLER_0_14_882 ();
 sg13g2_decap_8 FILLER_0_14_889 ();
 sg13g2_decap_8 FILLER_0_14_896 ();
 sg13g2_decap_8 FILLER_0_14_903 ();
 sg13g2_decap_8 FILLER_0_14_910 ();
 sg13g2_decap_8 FILLER_0_14_917 ();
 sg13g2_decap_8 FILLER_0_14_924 ();
 sg13g2_decap_8 FILLER_0_14_931 ();
 sg13g2_decap_8 FILLER_0_14_938 ();
 sg13g2_decap_8 FILLER_0_14_945 ();
 sg13g2_decap_8 FILLER_0_14_952 ();
 sg13g2_decap_8 FILLER_0_14_959 ();
 sg13g2_decap_8 FILLER_0_14_966 ();
 sg13g2_decap_8 FILLER_0_14_973 ();
 sg13g2_decap_8 FILLER_0_14_980 ();
 sg13g2_decap_8 FILLER_0_14_987 ();
 sg13g2_decap_8 FILLER_0_14_994 ();
 sg13g2_decap_8 FILLER_0_14_1001 ();
 sg13g2_decap_8 FILLER_0_14_1008 ();
 sg13g2_decap_8 FILLER_0_14_1015 ();
 sg13g2_decap_8 FILLER_0_14_1022 ();
 sg13g2_decap_8 FILLER_0_14_1029 ();
 sg13g2_decap_8 FILLER_0_14_1036 ();
 sg13g2_decap_8 FILLER_0_14_1043 ();
 sg13g2_decap_8 FILLER_0_14_1050 ();
 sg13g2_decap_8 FILLER_0_14_1057 ();
 sg13g2_decap_8 FILLER_0_14_1064 ();
 sg13g2_decap_8 FILLER_0_14_1071 ();
 sg13g2_decap_8 FILLER_0_14_1078 ();
 sg13g2_decap_8 FILLER_0_14_1085 ();
 sg13g2_decap_8 FILLER_0_14_1092 ();
 sg13g2_decap_8 FILLER_0_14_1099 ();
 sg13g2_decap_8 FILLER_0_14_1106 ();
 sg13g2_decap_8 FILLER_0_14_1113 ();
 sg13g2_decap_8 FILLER_0_14_1120 ();
 sg13g2_decap_8 FILLER_0_14_1127 ();
 sg13g2_decap_8 FILLER_0_14_1134 ();
 sg13g2_decap_8 FILLER_0_14_1141 ();
 sg13g2_decap_8 FILLER_0_14_1148 ();
 sg13g2_decap_8 FILLER_0_14_1155 ();
 sg13g2_decap_8 FILLER_0_14_1162 ();
 sg13g2_decap_8 FILLER_0_14_1169 ();
 sg13g2_decap_8 FILLER_0_14_1176 ();
 sg13g2_decap_8 FILLER_0_14_1183 ();
 sg13g2_decap_8 FILLER_0_14_1190 ();
 sg13g2_decap_8 FILLER_0_14_1197 ();
 sg13g2_decap_8 FILLER_0_14_1204 ();
 sg13g2_decap_8 FILLER_0_14_1211 ();
 sg13g2_decap_8 FILLER_0_14_1218 ();
 sg13g2_fill_2 FILLER_0_14_1225 ();
 sg13g2_fill_1 FILLER_0_14_1227 ();
 sg13g2_decap_8 FILLER_0_15_0 ();
 sg13g2_decap_8 FILLER_0_15_7 ();
 sg13g2_decap_8 FILLER_0_15_14 ();
 sg13g2_decap_8 FILLER_0_15_21 ();
 sg13g2_decap_8 FILLER_0_15_28 ();
 sg13g2_decap_8 FILLER_0_15_35 ();
 sg13g2_decap_8 FILLER_0_15_42 ();
 sg13g2_decap_8 FILLER_0_15_49 ();
 sg13g2_decap_8 FILLER_0_15_56 ();
 sg13g2_decap_8 FILLER_0_15_63 ();
 sg13g2_decap_8 FILLER_0_15_70 ();
 sg13g2_decap_8 FILLER_0_15_77 ();
 sg13g2_decap_8 FILLER_0_15_84 ();
 sg13g2_decap_8 FILLER_0_15_91 ();
 sg13g2_decap_8 FILLER_0_15_98 ();
 sg13g2_decap_8 FILLER_0_15_105 ();
 sg13g2_decap_8 FILLER_0_15_112 ();
 sg13g2_decap_8 FILLER_0_15_119 ();
 sg13g2_decap_8 FILLER_0_15_126 ();
 sg13g2_decap_8 FILLER_0_15_133 ();
 sg13g2_decap_8 FILLER_0_15_140 ();
 sg13g2_decap_8 FILLER_0_15_147 ();
 sg13g2_decap_8 FILLER_0_15_154 ();
 sg13g2_decap_8 FILLER_0_15_161 ();
 sg13g2_decap_8 FILLER_0_15_168 ();
 sg13g2_decap_8 FILLER_0_15_175 ();
 sg13g2_decap_8 FILLER_0_15_182 ();
 sg13g2_decap_8 FILLER_0_15_189 ();
 sg13g2_decap_8 FILLER_0_15_196 ();
 sg13g2_decap_8 FILLER_0_15_203 ();
 sg13g2_decap_8 FILLER_0_15_210 ();
 sg13g2_decap_8 FILLER_0_15_217 ();
 sg13g2_decap_8 FILLER_0_15_224 ();
 sg13g2_decap_8 FILLER_0_15_231 ();
 sg13g2_decap_8 FILLER_0_15_238 ();
 sg13g2_decap_8 FILLER_0_15_245 ();
 sg13g2_decap_8 FILLER_0_15_252 ();
 sg13g2_decap_8 FILLER_0_15_259 ();
 sg13g2_decap_8 FILLER_0_15_266 ();
 sg13g2_decap_8 FILLER_0_15_273 ();
 sg13g2_decap_8 FILLER_0_15_280 ();
 sg13g2_decap_8 FILLER_0_15_287 ();
 sg13g2_decap_8 FILLER_0_15_294 ();
 sg13g2_decap_8 FILLER_0_15_301 ();
 sg13g2_decap_8 FILLER_0_15_308 ();
 sg13g2_decap_8 FILLER_0_15_315 ();
 sg13g2_decap_8 FILLER_0_15_322 ();
 sg13g2_decap_8 FILLER_0_15_329 ();
 sg13g2_decap_8 FILLER_0_15_336 ();
 sg13g2_decap_8 FILLER_0_15_343 ();
 sg13g2_decap_8 FILLER_0_15_350 ();
 sg13g2_decap_8 FILLER_0_15_357 ();
 sg13g2_decap_8 FILLER_0_15_364 ();
 sg13g2_decap_8 FILLER_0_15_371 ();
 sg13g2_decap_8 FILLER_0_15_378 ();
 sg13g2_decap_8 FILLER_0_15_385 ();
 sg13g2_decap_8 FILLER_0_15_392 ();
 sg13g2_decap_8 FILLER_0_15_399 ();
 sg13g2_decap_8 FILLER_0_15_406 ();
 sg13g2_decap_8 FILLER_0_15_413 ();
 sg13g2_decap_8 FILLER_0_15_420 ();
 sg13g2_decap_8 FILLER_0_15_427 ();
 sg13g2_decap_8 FILLER_0_15_434 ();
 sg13g2_decap_8 FILLER_0_15_441 ();
 sg13g2_decap_8 FILLER_0_15_448 ();
 sg13g2_decap_8 FILLER_0_15_455 ();
 sg13g2_decap_8 FILLER_0_15_462 ();
 sg13g2_decap_8 FILLER_0_15_469 ();
 sg13g2_decap_8 FILLER_0_15_476 ();
 sg13g2_decap_8 FILLER_0_15_483 ();
 sg13g2_decap_8 FILLER_0_15_490 ();
 sg13g2_decap_8 FILLER_0_15_497 ();
 sg13g2_decap_8 FILLER_0_15_504 ();
 sg13g2_decap_8 FILLER_0_15_511 ();
 sg13g2_decap_8 FILLER_0_15_518 ();
 sg13g2_decap_8 FILLER_0_15_525 ();
 sg13g2_decap_8 FILLER_0_15_532 ();
 sg13g2_decap_8 FILLER_0_15_539 ();
 sg13g2_decap_8 FILLER_0_15_546 ();
 sg13g2_decap_8 FILLER_0_15_553 ();
 sg13g2_decap_8 FILLER_0_15_560 ();
 sg13g2_decap_8 FILLER_0_15_567 ();
 sg13g2_decap_8 FILLER_0_15_574 ();
 sg13g2_decap_8 FILLER_0_15_581 ();
 sg13g2_decap_8 FILLER_0_15_588 ();
 sg13g2_decap_8 FILLER_0_15_595 ();
 sg13g2_decap_8 FILLER_0_15_602 ();
 sg13g2_decap_8 FILLER_0_15_609 ();
 sg13g2_decap_8 FILLER_0_15_616 ();
 sg13g2_decap_8 FILLER_0_15_623 ();
 sg13g2_decap_8 FILLER_0_15_630 ();
 sg13g2_decap_8 FILLER_0_15_637 ();
 sg13g2_decap_8 FILLER_0_15_644 ();
 sg13g2_decap_8 FILLER_0_15_651 ();
 sg13g2_decap_8 FILLER_0_15_658 ();
 sg13g2_decap_8 FILLER_0_15_665 ();
 sg13g2_decap_8 FILLER_0_15_672 ();
 sg13g2_decap_8 FILLER_0_15_679 ();
 sg13g2_decap_8 FILLER_0_15_686 ();
 sg13g2_decap_8 FILLER_0_15_693 ();
 sg13g2_decap_8 FILLER_0_15_700 ();
 sg13g2_decap_8 FILLER_0_15_707 ();
 sg13g2_decap_8 FILLER_0_15_714 ();
 sg13g2_decap_8 FILLER_0_15_721 ();
 sg13g2_decap_8 FILLER_0_15_728 ();
 sg13g2_decap_8 FILLER_0_15_735 ();
 sg13g2_decap_8 FILLER_0_15_742 ();
 sg13g2_decap_8 FILLER_0_15_749 ();
 sg13g2_decap_8 FILLER_0_15_756 ();
 sg13g2_decap_8 FILLER_0_15_763 ();
 sg13g2_decap_8 FILLER_0_15_770 ();
 sg13g2_decap_8 FILLER_0_15_777 ();
 sg13g2_decap_8 FILLER_0_15_784 ();
 sg13g2_decap_8 FILLER_0_15_791 ();
 sg13g2_decap_8 FILLER_0_15_798 ();
 sg13g2_decap_8 FILLER_0_15_805 ();
 sg13g2_decap_8 FILLER_0_15_812 ();
 sg13g2_decap_8 FILLER_0_15_819 ();
 sg13g2_decap_8 FILLER_0_15_826 ();
 sg13g2_decap_8 FILLER_0_15_833 ();
 sg13g2_decap_8 FILLER_0_15_840 ();
 sg13g2_decap_8 FILLER_0_15_847 ();
 sg13g2_decap_8 FILLER_0_15_854 ();
 sg13g2_decap_8 FILLER_0_15_861 ();
 sg13g2_decap_8 FILLER_0_15_868 ();
 sg13g2_decap_8 FILLER_0_15_875 ();
 sg13g2_decap_8 FILLER_0_15_882 ();
 sg13g2_decap_8 FILLER_0_15_889 ();
 sg13g2_decap_8 FILLER_0_15_896 ();
 sg13g2_decap_8 FILLER_0_15_903 ();
 sg13g2_decap_8 FILLER_0_15_910 ();
 sg13g2_decap_8 FILLER_0_15_917 ();
 sg13g2_decap_8 FILLER_0_15_924 ();
 sg13g2_decap_8 FILLER_0_15_931 ();
 sg13g2_decap_8 FILLER_0_15_938 ();
 sg13g2_decap_8 FILLER_0_15_945 ();
 sg13g2_decap_8 FILLER_0_15_952 ();
 sg13g2_decap_8 FILLER_0_15_959 ();
 sg13g2_decap_8 FILLER_0_15_966 ();
 sg13g2_decap_8 FILLER_0_15_973 ();
 sg13g2_decap_8 FILLER_0_15_980 ();
 sg13g2_decap_8 FILLER_0_15_987 ();
 sg13g2_decap_8 FILLER_0_15_994 ();
 sg13g2_decap_8 FILLER_0_15_1001 ();
 sg13g2_decap_8 FILLER_0_15_1008 ();
 sg13g2_decap_8 FILLER_0_15_1015 ();
 sg13g2_decap_8 FILLER_0_15_1022 ();
 sg13g2_decap_8 FILLER_0_15_1029 ();
 sg13g2_decap_8 FILLER_0_15_1036 ();
 sg13g2_decap_8 FILLER_0_15_1043 ();
 sg13g2_decap_8 FILLER_0_15_1050 ();
 sg13g2_decap_8 FILLER_0_15_1057 ();
 sg13g2_decap_8 FILLER_0_15_1064 ();
 sg13g2_decap_8 FILLER_0_15_1071 ();
 sg13g2_decap_8 FILLER_0_15_1078 ();
 sg13g2_decap_8 FILLER_0_15_1085 ();
 sg13g2_decap_8 FILLER_0_15_1092 ();
 sg13g2_decap_8 FILLER_0_15_1099 ();
 sg13g2_decap_8 FILLER_0_15_1106 ();
 sg13g2_decap_8 FILLER_0_15_1113 ();
 sg13g2_decap_8 FILLER_0_15_1120 ();
 sg13g2_decap_8 FILLER_0_15_1127 ();
 sg13g2_decap_8 FILLER_0_15_1134 ();
 sg13g2_decap_8 FILLER_0_15_1141 ();
 sg13g2_decap_8 FILLER_0_15_1148 ();
 sg13g2_decap_8 FILLER_0_15_1155 ();
 sg13g2_decap_8 FILLER_0_15_1162 ();
 sg13g2_decap_8 FILLER_0_15_1169 ();
 sg13g2_decap_8 FILLER_0_15_1176 ();
 sg13g2_decap_8 FILLER_0_15_1183 ();
 sg13g2_decap_8 FILLER_0_15_1190 ();
 sg13g2_decap_8 FILLER_0_15_1197 ();
 sg13g2_decap_8 FILLER_0_15_1204 ();
 sg13g2_decap_8 FILLER_0_15_1211 ();
 sg13g2_decap_8 FILLER_0_15_1218 ();
 sg13g2_fill_2 FILLER_0_15_1225 ();
 sg13g2_fill_1 FILLER_0_15_1227 ();
 sg13g2_decap_8 FILLER_0_16_0 ();
 sg13g2_decap_8 FILLER_0_16_7 ();
 sg13g2_decap_8 FILLER_0_16_14 ();
 sg13g2_decap_8 FILLER_0_16_21 ();
 sg13g2_decap_8 FILLER_0_16_28 ();
 sg13g2_decap_8 FILLER_0_16_35 ();
 sg13g2_decap_8 FILLER_0_16_42 ();
 sg13g2_decap_8 FILLER_0_16_49 ();
 sg13g2_decap_8 FILLER_0_16_56 ();
 sg13g2_decap_8 FILLER_0_16_63 ();
 sg13g2_decap_8 FILLER_0_16_70 ();
 sg13g2_decap_8 FILLER_0_16_77 ();
 sg13g2_decap_8 FILLER_0_16_84 ();
 sg13g2_decap_8 FILLER_0_16_91 ();
 sg13g2_decap_8 FILLER_0_16_98 ();
 sg13g2_decap_8 FILLER_0_16_105 ();
 sg13g2_decap_8 FILLER_0_16_112 ();
 sg13g2_decap_8 FILLER_0_16_119 ();
 sg13g2_decap_8 FILLER_0_16_126 ();
 sg13g2_decap_8 FILLER_0_16_133 ();
 sg13g2_decap_8 FILLER_0_16_140 ();
 sg13g2_decap_8 FILLER_0_16_147 ();
 sg13g2_decap_8 FILLER_0_16_154 ();
 sg13g2_decap_8 FILLER_0_16_161 ();
 sg13g2_decap_8 FILLER_0_16_168 ();
 sg13g2_decap_8 FILLER_0_16_175 ();
 sg13g2_decap_8 FILLER_0_16_182 ();
 sg13g2_decap_8 FILLER_0_16_189 ();
 sg13g2_decap_8 FILLER_0_16_196 ();
 sg13g2_decap_8 FILLER_0_16_203 ();
 sg13g2_decap_8 FILLER_0_16_210 ();
 sg13g2_decap_8 FILLER_0_16_217 ();
 sg13g2_decap_8 FILLER_0_16_224 ();
 sg13g2_decap_8 FILLER_0_16_231 ();
 sg13g2_decap_8 FILLER_0_16_238 ();
 sg13g2_decap_8 FILLER_0_16_245 ();
 sg13g2_decap_8 FILLER_0_16_252 ();
 sg13g2_decap_8 FILLER_0_16_259 ();
 sg13g2_decap_8 FILLER_0_16_266 ();
 sg13g2_decap_8 FILLER_0_16_273 ();
 sg13g2_decap_8 FILLER_0_16_280 ();
 sg13g2_decap_8 FILLER_0_16_287 ();
 sg13g2_decap_8 FILLER_0_16_294 ();
 sg13g2_decap_8 FILLER_0_16_301 ();
 sg13g2_decap_8 FILLER_0_16_308 ();
 sg13g2_decap_8 FILLER_0_16_315 ();
 sg13g2_decap_8 FILLER_0_16_322 ();
 sg13g2_decap_8 FILLER_0_16_329 ();
 sg13g2_decap_8 FILLER_0_16_336 ();
 sg13g2_decap_8 FILLER_0_16_343 ();
 sg13g2_decap_8 FILLER_0_16_350 ();
 sg13g2_decap_8 FILLER_0_16_357 ();
 sg13g2_decap_8 FILLER_0_16_364 ();
 sg13g2_decap_8 FILLER_0_16_371 ();
 sg13g2_decap_8 FILLER_0_16_378 ();
 sg13g2_decap_8 FILLER_0_16_385 ();
 sg13g2_decap_8 FILLER_0_16_392 ();
 sg13g2_decap_8 FILLER_0_16_399 ();
 sg13g2_decap_8 FILLER_0_16_406 ();
 sg13g2_decap_8 FILLER_0_16_413 ();
 sg13g2_decap_8 FILLER_0_16_420 ();
 sg13g2_decap_8 FILLER_0_16_427 ();
 sg13g2_decap_8 FILLER_0_16_434 ();
 sg13g2_decap_8 FILLER_0_16_441 ();
 sg13g2_decap_8 FILLER_0_16_448 ();
 sg13g2_decap_8 FILLER_0_16_455 ();
 sg13g2_decap_8 FILLER_0_16_462 ();
 sg13g2_decap_8 FILLER_0_16_469 ();
 sg13g2_decap_8 FILLER_0_16_476 ();
 sg13g2_decap_8 FILLER_0_16_483 ();
 sg13g2_decap_8 FILLER_0_16_490 ();
 sg13g2_decap_8 FILLER_0_16_497 ();
 sg13g2_decap_8 FILLER_0_16_504 ();
 sg13g2_decap_8 FILLER_0_16_511 ();
 sg13g2_decap_8 FILLER_0_16_518 ();
 sg13g2_decap_8 FILLER_0_16_525 ();
 sg13g2_decap_8 FILLER_0_16_532 ();
 sg13g2_decap_8 FILLER_0_16_539 ();
 sg13g2_decap_8 FILLER_0_16_546 ();
 sg13g2_decap_8 FILLER_0_16_553 ();
 sg13g2_decap_8 FILLER_0_16_560 ();
 sg13g2_decap_8 FILLER_0_16_567 ();
 sg13g2_decap_8 FILLER_0_16_574 ();
 sg13g2_decap_8 FILLER_0_16_581 ();
 sg13g2_decap_8 FILLER_0_16_588 ();
 sg13g2_decap_8 FILLER_0_16_595 ();
 sg13g2_decap_8 FILLER_0_16_602 ();
 sg13g2_decap_8 FILLER_0_16_609 ();
 sg13g2_decap_8 FILLER_0_16_616 ();
 sg13g2_decap_8 FILLER_0_16_623 ();
 sg13g2_decap_8 FILLER_0_16_630 ();
 sg13g2_decap_8 FILLER_0_16_637 ();
 sg13g2_decap_8 FILLER_0_16_644 ();
 sg13g2_decap_8 FILLER_0_16_651 ();
 sg13g2_decap_8 FILLER_0_16_658 ();
 sg13g2_decap_8 FILLER_0_16_665 ();
 sg13g2_decap_8 FILLER_0_16_672 ();
 sg13g2_decap_8 FILLER_0_16_679 ();
 sg13g2_decap_8 FILLER_0_16_686 ();
 sg13g2_decap_8 FILLER_0_16_693 ();
 sg13g2_decap_8 FILLER_0_16_700 ();
 sg13g2_decap_8 FILLER_0_16_707 ();
 sg13g2_decap_8 FILLER_0_16_714 ();
 sg13g2_decap_8 FILLER_0_16_721 ();
 sg13g2_decap_8 FILLER_0_16_728 ();
 sg13g2_decap_8 FILLER_0_16_735 ();
 sg13g2_decap_8 FILLER_0_16_742 ();
 sg13g2_decap_8 FILLER_0_16_749 ();
 sg13g2_decap_8 FILLER_0_16_756 ();
 sg13g2_decap_8 FILLER_0_16_763 ();
 sg13g2_decap_8 FILLER_0_16_770 ();
 sg13g2_decap_8 FILLER_0_16_777 ();
 sg13g2_decap_8 FILLER_0_16_784 ();
 sg13g2_decap_8 FILLER_0_16_791 ();
 sg13g2_decap_8 FILLER_0_16_798 ();
 sg13g2_decap_8 FILLER_0_16_805 ();
 sg13g2_decap_8 FILLER_0_16_812 ();
 sg13g2_decap_8 FILLER_0_16_819 ();
 sg13g2_decap_8 FILLER_0_16_826 ();
 sg13g2_decap_8 FILLER_0_16_833 ();
 sg13g2_decap_8 FILLER_0_16_840 ();
 sg13g2_decap_8 FILLER_0_16_847 ();
 sg13g2_decap_8 FILLER_0_16_854 ();
 sg13g2_decap_8 FILLER_0_16_861 ();
 sg13g2_decap_8 FILLER_0_16_868 ();
 sg13g2_decap_8 FILLER_0_16_875 ();
 sg13g2_decap_8 FILLER_0_16_882 ();
 sg13g2_decap_8 FILLER_0_16_889 ();
 sg13g2_decap_8 FILLER_0_16_896 ();
 sg13g2_decap_8 FILLER_0_16_903 ();
 sg13g2_decap_8 FILLER_0_16_910 ();
 sg13g2_decap_8 FILLER_0_16_917 ();
 sg13g2_decap_8 FILLER_0_16_924 ();
 sg13g2_decap_8 FILLER_0_16_931 ();
 sg13g2_decap_8 FILLER_0_16_938 ();
 sg13g2_decap_8 FILLER_0_16_945 ();
 sg13g2_decap_8 FILLER_0_16_952 ();
 sg13g2_decap_8 FILLER_0_16_959 ();
 sg13g2_decap_8 FILLER_0_16_966 ();
 sg13g2_decap_8 FILLER_0_16_973 ();
 sg13g2_decap_8 FILLER_0_16_980 ();
 sg13g2_decap_8 FILLER_0_16_987 ();
 sg13g2_decap_8 FILLER_0_16_994 ();
 sg13g2_decap_8 FILLER_0_16_1001 ();
 sg13g2_decap_8 FILLER_0_16_1008 ();
 sg13g2_decap_8 FILLER_0_16_1015 ();
 sg13g2_decap_8 FILLER_0_16_1022 ();
 sg13g2_decap_8 FILLER_0_16_1029 ();
 sg13g2_decap_8 FILLER_0_16_1036 ();
 sg13g2_decap_8 FILLER_0_16_1043 ();
 sg13g2_decap_8 FILLER_0_16_1050 ();
 sg13g2_decap_8 FILLER_0_16_1057 ();
 sg13g2_decap_8 FILLER_0_16_1064 ();
 sg13g2_decap_8 FILLER_0_16_1071 ();
 sg13g2_decap_8 FILLER_0_16_1078 ();
 sg13g2_decap_8 FILLER_0_16_1085 ();
 sg13g2_decap_8 FILLER_0_16_1092 ();
 sg13g2_decap_8 FILLER_0_16_1099 ();
 sg13g2_decap_8 FILLER_0_16_1106 ();
 sg13g2_decap_8 FILLER_0_16_1113 ();
 sg13g2_decap_8 FILLER_0_16_1120 ();
 sg13g2_decap_8 FILLER_0_16_1127 ();
 sg13g2_decap_8 FILLER_0_16_1134 ();
 sg13g2_decap_8 FILLER_0_16_1141 ();
 sg13g2_decap_8 FILLER_0_16_1148 ();
 sg13g2_decap_8 FILLER_0_16_1155 ();
 sg13g2_decap_8 FILLER_0_16_1162 ();
 sg13g2_decap_8 FILLER_0_16_1169 ();
 sg13g2_decap_8 FILLER_0_16_1176 ();
 sg13g2_decap_8 FILLER_0_16_1183 ();
 sg13g2_decap_8 FILLER_0_16_1190 ();
 sg13g2_decap_8 FILLER_0_16_1197 ();
 sg13g2_decap_8 FILLER_0_16_1204 ();
 sg13g2_decap_8 FILLER_0_16_1211 ();
 sg13g2_decap_8 FILLER_0_16_1218 ();
 sg13g2_fill_2 FILLER_0_16_1225 ();
 sg13g2_fill_1 FILLER_0_16_1227 ();
 sg13g2_decap_8 FILLER_0_17_0 ();
 sg13g2_decap_8 FILLER_0_17_7 ();
 sg13g2_decap_8 FILLER_0_17_14 ();
 sg13g2_decap_8 FILLER_0_17_21 ();
 sg13g2_decap_8 FILLER_0_17_28 ();
 sg13g2_decap_8 FILLER_0_17_35 ();
 sg13g2_decap_8 FILLER_0_17_42 ();
 sg13g2_decap_8 FILLER_0_17_49 ();
 sg13g2_decap_8 FILLER_0_17_56 ();
 sg13g2_decap_8 FILLER_0_17_63 ();
 sg13g2_decap_8 FILLER_0_17_70 ();
 sg13g2_decap_8 FILLER_0_17_77 ();
 sg13g2_decap_8 FILLER_0_17_84 ();
 sg13g2_decap_8 FILLER_0_17_91 ();
 sg13g2_decap_8 FILLER_0_17_98 ();
 sg13g2_decap_8 FILLER_0_17_105 ();
 sg13g2_decap_8 FILLER_0_17_112 ();
 sg13g2_decap_8 FILLER_0_17_119 ();
 sg13g2_decap_8 FILLER_0_17_126 ();
 sg13g2_decap_8 FILLER_0_17_133 ();
 sg13g2_decap_8 FILLER_0_17_140 ();
 sg13g2_decap_8 FILLER_0_17_147 ();
 sg13g2_decap_8 FILLER_0_17_154 ();
 sg13g2_decap_8 FILLER_0_17_161 ();
 sg13g2_decap_8 FILLER_0_17_168 ();
 sg13g2_decap_8 FILLER_0_17_175 ();
 sg13g2_decap_8 FILLER_0_17_182 ();
 sg13g2_decap_8 FILLER_0_17_189 ();
 sg13g2_decap_8 FILLER_0_17_196 ();
 sg13g2_decap_8 FILLER_0_17_203 ();
 sg13g2_decap_8 FILLER_0_17_210 ();
 sg13g2_decap_8 FILLER_0_17_217 ();
 sg13g2_decap_8 FILLER_0_17_224 ();
 sg13g2_decap_8 FILLER_0_17_231 ();
 sg13g2_decap_8 FILLER_0_17_238 ();
 sg13g2_decap_8 FILLER_0_17_245 ();
 sg13g2_decap_8 FILLER_0_17_252 ();
 sg13g2_decap_8 FILLER_0_17_259 ();
 sg13g2_decap_8 FILLER_0_17_266 ();
 sg13g2_decap_8 FILLER_0_17_273 ();
 sg13g2_decap_8 FILLER_0_17_280 ();
 sg13g2_decap_8 FILLER_0_17_287 ();
 sg13g2_decap_8 FILLER_0_17_294 ();
 sg13g2_decap_8 FILLER_0_17_301 ();
 sg13g2_decap_8 FILLER_0_17_308 ();
 sg13g2_decap_8 FILLER_0_17_315 ();
 sg13g2_decap_8 FILLER_0_17_322 ();
 sg13g2_decap_8 FILLER_0_17_329 ();
 sg13g2_decap_8 FILLER_0_17_336 ();
 sg13g2_decap_8 FILLER_0_17_343 ();
 sg13g2_decap_8 FILLER_0_17_350 ();
 sg13g2_decap_8 FILLER_0_17_357 ();
 sg13g2_decap_8 FILLER_0_17_364 ();
 sg13g2_decap_8 FILLER_0_17_371 ();
 sg13g2_decap_8 FILLER_0_17_378 ();
 sg13g2_decap_8 FILLER_0_17_385 ();
 sg13g2_decap_8 FILLER_0_17_392 ();
 sg13g2_decap_8 FILLER_0_17_399 ();
 sg13g2_decap_8 FILLER_0_17_406 ();
 sg13g2_decap_8 FILLER_0_17_413 ();
 sg13g2_decap_8 FILLER_0_17_420 ();
 sg13g2_decap_8 FILLER_0_17_427 ();
 sg13g2_decap_8 FILLER_0_17_434 ();
 sg13g2_decap_8 FILLER_0_17_441 ();
 sg13g2_decap_8 FILLER_0_17_448 ();
 sg13g2_decap_8 FILLER_0_17_455 ();
 sg13g2_decap_8 FILLER_0_17_462 ();
 sg13g2_decap_8 FILLER_0_17_469 ();
 sg13g2_decap_8 FILLER_0_17_476 ();
 sg13g2_decap_8 FILLER_0_17_483 ();
 sg13g2_decap_8 FILLER_0_17_490 ();
 sg13g2_decap_8 FILLER_0_17_497 ();
 sg13g2_decap_8 FILLER_0_17_504 ();
 sg13g2_decap_8 FILLER_0_17_511 ();
 sg13g2_decap_8 FILLER_0_17_518 ();
 sg13g2_decap_8 FILLER_0_17_525 ();
 sg13g2_decap_8 FILLER_0_17_532 ();
 sg13g2_decap_8 FILLER_0_17_539 ();
 sg13g2_decap_8 FILLER_0_17_546 ();
 sg13g2_decap_8 FILLER_0_17_553 ();
 sg13g2_decap_8 FILLER_0_17_560 ();
 sg13g2_decap_8 FILLER_0_17_567 ();
 sg13g2_decap_8 FILLER_0_17_574 ();
 sg13g2_decap_8 FILLER_0_17_581 ();
 sg13g2_decap_8 FILLER_0_17_588 ();
 sg13g2_decap_8 FILLER_0_17_595 ();
 sg13g2_decap_8 FILLER_0_17_602 ();
 sg13g2_decap_8 FILLER_0_17_609 ();
 sg13g2_decap_8 FILLER_0_17_616 ();
 sg13g2_decap_8 FILLER_0_17_623 ();
 sg13g2_decap_8 FILLER_0_17_630 ();
 sg13g2_decap_8 FILLER_0_17_637 ();
 sg13g2_decap_8 FILLER_0_17_644 ();
 sg13g2_decap_8 FILLER_0_17_651 ();
 sg13g2_decap_8 FILLER_0_17_658 ();
 sg13g2_decap_8 FILLER_0_17_665 ();
 sg13g2_decap_8 FILLER_0_17_672 ();
 sg13g2_decap_8 FILLER_0_17_679 ();
 sg13g2_decap_8 FILLER_0_17_686 ();
 sg13g2_decap_8 FILLER_0_17_693 ();
 sg13g2_decap_8 FILLER_0_17_700 ();
 sg13g2_decap_8 FILLER_0_17_707 ();
 sg13g2_decap_8 FILLER_0_17_714 ();
 sg13g2_decap_8 FILLER_0_17_721 ();
 sg13g2_decap_8 FILLER_0_17_728 ();
 sg13g2_decap_8 FILLER_0_17_735 ();
 sg13g2_decap_8 FILLER_0_17_742 ();
 sg13g2_decap_8 FILLER_0_17_749 ();
 sg13g2_decap_8 FILLER_0_17_756 ();
 sg13g2_decap_8 FILLER_0_17_763 ();
 sg13g2_decap_8 FILLER_0_17_770 ();
 sg13g2_decap_8 FILLER_0_17_777 ();
 sg13g2_decap_8 FILLER_0_17_784 ();
 sg13g2_decap_8 FILLER_0_17_791 ();
 sg13g2_decap_8 FILLER_0_17_798 ();
 sg13g2_decap_8 FILLER_0_17_805 ();
 sg13g2_decap_8 FILLER_0_17_812 ();
 sg13g2_decap_8 FILLER_0_17_819 ();
 sg13g2_decap_8 FILLER_0_17_826 ();
 sg13g2_decap_8 FILLER_0_17_833 ();
 sg13g2_decap_8 FILLER_0_17_840 ();
 sg13g2_decap_8 FILLER_0_17_847 ();
 sg13g2_decap_8 FILLER_0_17_854 ();
 sg13g2_decap_8 FILLER_0_17_861 ();
 sg13g2_decap_8 FILLER_0_17_868 ();
 sg13g2_decap_8 FILLER_0_17_875 ();
 sg13g2_decap_8 FILLER_0_17_882 ();
 sg13g2_decap_8 FILLER_0_17_889 ();
 sg13g2_decap_8 FILLER_0_17_896 ();
 sg13g2_decap_8 FILLER_0_17_903 ();
 sg13g2_decap_8 FILLER_0_17_910 ();
 sg13g2_decap_8 FILLER_0_17_917 ();
 sg13g2_decap_8 FILLER_0_17_924 ();
 sg13g2_decap_8 FILLER_0_17_931 ();
 sg13g2_decap_8 FILLER_0_17_938 ();
 sg13g2_decap_8 FILLER_0_17_945 ();
 sg13g2_decap_8 FILLER_0_17_952 ();
 sg13g2_decap_8 FILLER_0_17_959 ();
 sg13g2_decap_8 FILLER_0_17_966 ();
 sg13g2_decap_8 FILLER_0_17_973 ();
 sg13g2_decap_8 FILLER_0_17_980 ();
 sg13g2_decap_8 FILLER_0_17_987 ();
 sg13g2_decap_8 FILLER_0_17_994 ();
 sg13g2_decap_8 FILLER_0_17_1001 ();
 sg13g2_decap_8 FILLER_0_17_1008 ();
 sg13g2_decap_8 FILLER_0_17_1015 ();
 sg13g2_decap_8 FILLER_0_17_1022 ();
 sg13g2_decap_8 FILLER_0_17_1029 ();
 sg13g2_decap_8 FILLER_0_17_1036 ();
 sg13g2_decap_8 FILLER_0_17_1043 ();
 sg13g2_decap_8 FILLER_0_17_1050 ();
 sg13g2_decap_8 FILLER_0_17_1057 ();
 sg13g2_decap_8 FILLER_0_17_1064 ();
 sg13g2_decap_8 FILLER_0_17_1071 ();
 sg13g2_decap_8 FILLER_0_17_1078 ();
 sg13g2_decap_8 FILLER_0_17_1085 ();
 sg13g2_decap_8 FILLER_0_17_1092 ();
 sg13g2_decap_8 FILLER_0_17_1099 ();
 sg13g2_decap_8 FILLER_0_17_1106 ();
 sg13g2_decap_8 FILLER_0_17_1113 ();
 sg13g2_decap_8 FILLER_0_17_1120 ();
 sg13g2_decap_8 FILLER_0_17_1127 ();
 sg13g2_decap_8 FILLER_0_17_1134 ();
 sg13g2_decap_8 FILLER_0_17_1141 ();
 sg13g2_decap_8 FILLER_0_17_1148 ();
 sg13g2_decap_8 FILLER_0_17_1155 ();
 sg13g2_decap_8 FILLER_0_17_1162 ();
 sg13g2_decap_8 FILLER_0_17_1169 ();
 sg13g2_decap_8 FILLER_0_17_1176 ();
 sg13g2_decap_8 FILLER_0_17_1183 ();
 sg13g2_decap_8 FILLER_0_17_1190 ();
 sg13g2_decap_8 FILLER_0_17_1197 ();
 sg13g2_decap_8 FILLER_0_17_1204 ();
 sg13g2_decap_8 FILLER_0_17_1211 ();
 sg13g2_decap_8 FILLER_0_17_1218 ();
 sg13g2_fill_2 FILLER_0_17_1225 ();
 sg13g2_fill_1 FILLER_0_17_1227 ();
 sg13g2_decap_8 FILLER_0_18_0 ();
 sg13g2_decap_8 FILLER_0_18_7 ();
 sg13g2_decap_8 FILLER_0_18_14 ();
 sg13g2_decap_8 FILLER_0_18_21 ();
 sg13g2_decap_8 FILLER_0_18_28 ();
 sg13g2_decap_8 FILLER_0_18_35 ();
 sg13g2_decap_8 FILLER_0_18_42 ();
 sg13g2_decap_8 FILLER_0_18_49 ();
 sg13g2_decap_8 FILLER_0_18_56 ();
 sg13g2_decap_8 FILLER_0_18_63 ();
 sg13g2_decap_8 FILLER_0_18_70 ();
 sg13g2_decap_8 FILLER_0_18_77 ();
 sg13g2_decap_8 FILLER_0_18_84 ();
 sg13g2_decap_8 FILLER_0_18_91 ();
 sg13g2_decap_8 FILLER_0_18_98 ();
 sg13g2_decap_8 FILLER_0_18_105 ();
 sg13g2_decap_8 FILLER_0_18_112 ();
 sg13g2_decap_8 FILLER_0_18_119 ();
 sg13g2_decap_8 FILLER_0_18_126 ();
 sg13g2_decap_8 FILLER_0_18_133 ();
 sg13g2_decap_8 FILLER_0_18_140 ();
 sg13g2_decap_8 FILLER_0_18_147 ();
 sg13g2_decap_8 FILLER_0_18_154 ();
 sg13g2_decap_8 FILLER_0_18_161 ();
 sg13g2_decap_8 FILLER_0_18_168 ();
 sg13g2_decap_8 FILLER_0_18_175 ();
 sg13g2_decap_8 FILLER_0_18_182 ();
 sg13g2_decap_8 FILLER_0_18_189 ();
 sg13g2_decap_8 FILLER_0_18_196 ();
 sg13g2_decap_8 FILLER_0_18_203 ();
 sg13g2_decap_8 FILLER_0_18_210 ();
 sg13g2_decap_8 FILLER_0_18_217 ();
 sg13g2_decap_8 FILLER_0_18_224 ();
 sg13g2_decap_8 FILLER_0_18_231 ();
 sg13g2_decap_8 FILLER_0_18_238 ();
 sg13g2_decap_8 FILLER_0_18_245 ();
 sg13g2_decap_8 FILLER_0_18_252 ();
 sg13g2_decap_8 FILLER_0_18_259 ();
 sg13g2_decap_8 FILLER_0_18_266 ();
 sg13g2_decap_8 FILLER_0_18_273 ();
 sg13g2_decap_8 FILLER_0_18_280 ();
 sg13g2_decap_8 FILLER_0_18_287 ();
 sg13g2_decap_8 FILLER_0_18_294 ();
 sg13g2_decap_8 FILLER_0_18_301 ();
 sg13g2_decap_8 FILLER_0_18_308 ();
 sg13g2_decap_8 FILLER_0_18_315 ();
 sg13g2_decap_8 FILLER_0_18_322 ();
 sg13g2_decap_8 FILLER_0_18_329 ();
 sg13g2_decap_8 FILLER_0_18_336 ();
 sg13g2_decap_8 FILLER_0_18_343 ();
 sg13g2_decap_8 FILLER_0_18_350 ();
 sg13g2_decap_8 FILLER_0_18_357 ();
 sg13g2_decap_8 FILLER_0_18_364 ();
 sg13g2_decap_8 FILLER_0_18_371 ();
 sg13g2_decap_8 FILLER_0_18_378 ();
 sg13g2_decap_8 FILLER_0_18_385 ();
 sg13g2_decap_8 FILLER_0_18_392 ();
 sg13g2_decap_8 FILLER_0_18_399 ();
 sg13g2_decap_8 FILLER_0_18_406 ();
 sg13g2_decap_8 FILLER_0_18_413 ();
 sg13g2_decap_8 FILLER_0_18_420 ();
 sg13g2_decap_8 FILLER_0_18_427 ();
 sg13g2_decap_8 FILLER_0_18_434 ();
 sg13g2_decap_8 FILLER_0_18_441 ();
 sg13g2_decap_8 FILLER_0_18_448 ();
 sg13g2_decap_8 FILLER_0_18_455 ();
 sg13g2_decap_8 FILLER_0_18_462 ();
 sg13g2_decap_8 FILLER_0_18_469 ();
 sg13g2_decap_8 FILLER_0_18_476 ();
 sg13g2_decap_8 FILLER_0_18_483 ();
 sg13g2_decap_8 FILLER_0_18_490 ();
 sg13g2_decap_8 FILLER_0_18_497 ();
 sg13g2_decap_8 FILLER_0_18_504 ();
 sg13g2_decap_8 FILLER_0_18_511 ();
 sg13g2_decap_8 FILLER_0_18_518 ();
 sg13g2_decap_8 FILLER_0_18_525 ();
 sg13g2_decap_8 FILLER_0_18_532 ();
 sg13g2_decap_8 FILLER_0_18_539 ();
 sg13g2_decap_8 FILLER_0_18_546 ();
 sg13g2_decap_8 FILLER_0_18_553 ();
 sg13g2_decap_8 FILLER_0_18_560 ();
 sg13g2_decap_8 FILLER_0_18_567 ();
 sg13g2_decap_8 FILLER_0_18_574 ();
 sg13g2_decap_8 FILLER_0_18_581 ();
 sg13g2_decap_8 FILLER_0_18_588 ();
 sg13g2_decap_8 FILLER_0_18_595 ();
 sg13g2_decap_8 FILLER_0_18_602 ();
 sg13g2_decap_8 FILLER_0_18_609 ();
 sg13g2_decap_8 FILLER_0_18_616 ();
 sg13g2_decap_8 FILLER_0_18_623 ();
 sg13g2_decap_8 FILLER_0_18_630 ();
 sg13g2_decap_8 FILLER_0_18_637 ();
 sg13g2_decap_8 FILLER_0_18_644 ();
 sg13g2_decap_8 FILLER_0_18_651 ();
 sg13g2_decap_8 FILLER_0_18_658 ();
 sg13g2_decap_8 FILLER_0_18_665 ();
 sg13g2_decap_8 FILLER_0_18_672 ();
 sg13g2_decap_8 FILLER_0_18_679 ();
 sg13g2_decap_8 FILLER_0_18_686 ();
 sg13g2_decap_8 FILLER_0_18_693 ();
 sg13g2_decap_8 FILLER_0_18_700 ();
 sg13g2_decap_8 FILLER_0_18_707 ();
 sg13g2_decap_8 FILLER_0_18_714 ();
 sg13g2_decap_8 FILLER_0_18_721 ();
 sg13g2_decap_8 FILLER_0_18_728 ();
 sg13g2_decap_8 FILLER_0_18_735 ();
 sg13g2_decap_8 FILLER_0_18_742 ();
 sg13g2_decap_8 FILLER_0_18_749 ();
 sg13g2_decap_8 FILLER_0_18_756 ();
 sg13g2_decap_8 FILLER_0_18_763 ();
 sg13g2_decap_8 FILLER_0_18_770 ();
 sg13g2_decap_8 FILLER_0_18_777 ();
 sg13g2_decap_8 FILLER_0_18_784 ();
 sg13g2_decap_8 FILLER_0_18_791 ();
 sg13g2_decap_8 FILLER_0_18_798 ();
 sg13g2_decap_8 FILLER_0_18_805 ();
 sg13g2_decap_8 FILLER_0_18_812 ();
 sg13g2_decap_8 FILLER_0_18_819 ();
 sg13g2_decap_8 FILLER_0_18_826 ();
 sg13g2_decap_8 FILLER_0_18_833 ();
 sg13g2_decap_8 FILLER_0_18_840 ();
 sg13g2_decap_8 FILLER_0_18_847 ();
 sg13g2_decap_8 FILLER_0_18_854 ();
 sg13g2_decap_8 FILLER_0_18_861 ();
 sg13g2_decap_8 FILLER_0_18_868 ();
 sg13g2_decap_8 FILLER_0_18_875 ();
 sg13g2_decap_8 FILLER_0_18_882 ();
 sg13g2_decap_8 FILLER_0_18_889 ();
 sg13g2_decap_8 FILLER_0_18_896 ();
 sg13g2_decap_8 FILLER_0_18_903 ();
 sg13g2_decap_8 FILLER_0_18_910 ();
 sg13g2_decap_8 FILLER_0_18_917 ();
 sg13g2_decap_8 FILLER_0_18_924 ();
 sg13g2_decap_8 FILLER_0_18_931 ();
 sg13g2_decap_8 FILLER_0_18_938 ();
 sg13g2_decap_8 FILLER_0_18_945 ();
 sg13g2_decap_8 FILLER_0_18_952 ();
 sg13g2_decap_8 FILLER_0_18_959 ();
 sg13g2_decap_8 FILLER_0_18_966 ();
 sg13g2_decap_8 FILLER_0_18_973 ();
 sg13g2_decap_8 FILLER_0_18_980 ();
 sg13g2_decap_8 FILLER_0_18_987 ();
 sg13g2_decap_8 FILLER_0_18_994 ();
 sg13g2_decap_8 FILLER_0_18_1001 ();
 sg13g2_decap_8 FILLER_0_18_1008 ();
 sg13g2_decap_8 FILLER_0_18_1015 ();
 sg13g2_decap_8 FILLER_0_18_1022 ();
 sg13g2_decap_8 FILLER_0_18_1029 ();
 sg13g2_decap_8 FILLER_0_18_1036 ();
 sg13g2_decap_8 FILLER_0_18_1043 ();
 sg13g2_decap_8 FILLER_0_18_1050 ();
 sg13g2_decap_8 FILLER_0_18_1057 ();
 sg13g2_decap_8 FILLER_0_18_1064 ();
 sg13g2_decap_8 FILLER_0_18_1071 ();
 sg13g2_decap_8 FILLER_0_18_1078 ();
 sg13g2_decap_8 FILLER_0_18_1085 ();
 sg13g2_decap_8 FILLER_0_18_1092 ();
 sg13g2_decap_8 FILLER_0_18_1099 ();
 sg13g2_decap_8 FILLER_0_18_1106 ();
 sg13g2_decap_8 FILLER_0_18_1113 ();
 sg13g2_decap_8 FILLER_0_18_1120 ();
 sg13g2_decap_8 FILLER_0_18_1127 ();
 sg13g2_decap_8 FILLER_0_18_1134 ();
 sg13g2_decap_8 FILLER_0_18_1141 ();
 sg13g2_decap_8 FILLER_0_18_1148 ();
 sg13g2_decap_8 FILLER_0_18_1155 ();
 sg13g2_decap_8 FILLER_0_18_1162 ();
 sg13g2_decap_8 FILLER_0_18_1169 ();
 sg13g2_decap_8 FILLER_0_18_1176 ();
 sg13g2_decap_8 FILLER_0_18_1183 ();
 sg13g2_decap_8 FILLER_0_18_1190 ();
 sg13g2_decap_8 FILLER_0_18_1197 ();
 sg13g2_decap_8 FILLER_0_18_1204 ();
 sg13g2_decap_8 FILLER_0_18_1211 ();
 sg13g2_decap_8 FILLER_0_18_1218 ();
 sg13g2_fill_2 FILLER_0_18_1225 ();
 sg13g2_fill_1 FILLER_0_18_1227 ();
 sg13g2_decap_8 FILLER_0_19_0 ();
 sg13g2_decap_8 FILLER_0_19_7 ();
 sg13g2_decap_8 FILLER_0_19_14 ();
 sg13g2_decap_8 FILLER_0_19_21 ();
 sg13g2_decap_8 FILLER_0_19_28 ();
 sg13g2_decap_8 FILLER_0_19_35 ();
 sg13g2_decap_8 FILLER_0_19_42 ();
 sg13g2_decap_8 FILLER_0_19_49 ();
 sg13g2_decap_8 FILLER_0_19_56 ();
 sg13g2_decap_8 FILLER_0_19_63 ();
 sg13g2_decap_8 FILLER_0_19_70 ();
 sg13g2_decap_8 FILLER_0_19_77 ();
 sg13g2_decap_8 FILLER_0_19_84 ();
 sg13g2_decap_8 FILLER_0_19_91 ();
 sg13g2_decap_8 FILLER_0_19_98 ();
 sg13g2_decap_8 FILLER_0_19_105 ();
 sg13g2_decap_8 FILLER_0_19_112 ();
 sg13g2_decap_8 FILLER_0_19_119 ();
 sg13g2_decap_8 FILLER_0_19_126 ();
 sg13g2_decap_8 FILLER_0_19_133 ();
 sg13g2_decap_8 FILLER_0_19_140 ();
 sg13g2_decap_8 FILLER_0_19_147 ();
 sg13g2_decap_8 FILLER_0_19_154 ();
 sg13g2_decap_8 FILLER_0_19_161 ();
 sg13g2_decap_8 FILLER_0_19_168 ();
 sg13g2_decap_8 FILLER_0_19_175 ();
 sg13g2_decap_8 FILLER_0_19_182 ();
 sg13g2_decap_8 FILLER_0_19_189 ();
 sg13g2_decap_8 FILLER_0_19_196 ();
 sg13g2_decap_8 FILLER_0_19_203 ();
 sg13g2_decap_8 FILLER_0_19_210 ();
 sg13g2_decap_8 FILLER_0_19_217 ();
 sg13g2_decap_8 FILLER_0_19_224 ();
 sg13g2_decap_8 FILLER_0_19_231 ();
 sg13g2_decap_8 FILLER_0_19_238 ();
 sg13g2_decap_8 FILLER_0_19_245 ();
 sg13g2_decap_8 FILLER_0_19_252 ();
 sg13g2_decap_8 FILLER_0_19_259 ();
 sg13g2_decap_8 FILLER_0_19_266 ();
 sg13g2_decap_8 FILLER_0_19_273 ();
 sg13g2_decap_8 FILLER_0_19_280 ();
 sg13g2_decap_8 FILLER_0_19_287 ();
 sg13g2_decap_8 FILLER_0_19_294 ();
 sg13g2_decap_8 FILLER_0_19_301 ();
 sg13g2_decap_8 FILLER_0_19_308 ();
 sg13g2_decap_8 FILLER_0_19_315 ();
 sg13g2_decap_8 FILLER_0_19_322 ();
 sg13g2_decap_8 FILLER_0_19_329 ();
 sg13g2_decap_8 FILLER_0_19_336 ();
 sg13g2_decap_8 FILLER_0_19_343 ();
 sg13g2_decap_8 FILLER_0_19_350 ();
 sg13g2_decap_8 FILLER_0_19_357 ();
 sg13g2_decap_8 FILLER_0_19_364 ();
 sg13g2_decap_8 FILLER_0_19_371 ();
 sg13g2_decap_8 FILLER_0_19_378 ();
 sg13g2_decap_8 FILLER_0_19_385 ();
 sg13g2_decap_8 FILLER_0_19_392 ();
 sg13g2_decap_8 FILLER_0_19_399 ();
 sg13g2_decap_8 FILLER_0_19_406 ();
 sg13g2_decap_8 FILLER_0_19_413 ();
 sg13g2_decap_8 FILLER_0_19_420 ();
 sg13g2_decap_8 FILLER_0_19_427 ();
 sg13g2_decap_8 FILLER_0_19_434 ();
 sg13g2_decap_8 FILLER_0_19_441 ();
 sg13g2_decap_8 FILLER_0_19_448 ();
 sg13g2_decap_8 FILLER_0_19_455 ();
 sg13g2_decap_8 FILLER_0_19_462 ();
 sg13g2_decap_8 FILLER_0_19_469 ();
 sg13g2_decap_8 FILLER_0_19_476 ();
 sg13g2_decap_8 FILLER_0_19_483 ();
 sg13g2_decap_8 FILLER_0_19_490 ();
 sg13g2_decap_8 FILLER_0_19_497 ();
 sg13g2_decap_8 FILLER_0_19_504 ();
 sg13g2_decap_8 FILLER_0_19_511 ();
 sg13g2_decap_8 FILLER_0_19_518 ();
 sg13g2_decap_8 FILLER_0_19_525 ();
 sg13g2_decap_8 FILLER_0_19_532 ();
 sg13g2_decap_8 FILLER_0_19_539 ();
 sg13g2_decap_8 FILLER_0_19_546 ();
 sg13g2_decap_8 FILLER_0_19_553 ();
 sg13g2_decap_8 FILLER_0_19_560 ();
 sg13g2_decap_8 FILLER_0_19_567 ();
 sg13g2_decap_8 FILLER_0_19_574 ();
 sg13g2_decap_8 FILLER_0_19_581 ();
 sg13g2_decap_8 FILLER_0_19_588 ();
 sg13g2_decap_8 FILLER_0_19_595 ();
 sg13g2_decap_8 FILLER_0_19_602 ();
 sg13g2_decap_8 FILLER_0_19_609 ();
 sg13g2_decap_8 FILLER_0_19_616 ();
 sg13g2_decap_8 FILLER_0_19_623 ();
 sg13g2_decap_8 FILLER_0_19_630 ();
 sg13g2_decap_8 FILLER_0_19_637 ();
 sg13g2_decap_8 FILLER_0_19_644 ();
 sg13g2_decap_8 FILLER_0_19_651 ();
 sg13g2_decap_8 FILLER_0_19_658 ();
 sg13g2_decap_8 FILLER_0_19_665 ();
 sg13g2_decap_8 FILLER_0_19_672 ();
 sg13g2_decap_8 FILLER_0_19_679 ();
 sg13g2_decap_8 FILLER_0_19_686 ();
 sg13g2_decap_8 FILLER_0_19_693 ();
 sg13g2_decap_8 FILLER_0_19_700 ();
 sg13g2_decap_8 FILLER_0_19_707 ();
 sg13g2_decap_8 FILLER_0_19_714 ();
 sg13g2_decap_8 FILLER_0_19_721 ();
 sg13g2_decap_8 FILLER_0_19_728 ();
 sg13g2_decap_8 FILLER_0_19_735 ();
 sg13g2_decap_8 FILLER_0_19_742 ();
 sg13g2_decap_8 FILLER_0_19_749 ();
 sg13g2_decap_8 FILLER_0_19_756 ();
 sg13g2_decap_8 FILLER_0_19_763 ();
 sg13g2_decap_8 FILLER_0_19_770 ();
 sg13g2_decap_8 FILLER_0_19_777 ();
 sg13g2_decap_8 FILLER_0_19_784 ();
 sg13g2_decap_8 FILLER_0_19_791 ();
 sg13g2_decap_8 FILLER_0_19_798 ();
 sg13g2_decap_8 FILLER_0_19_805 ();
 sg13g2_decap_8 FILLER_0_19_812 ();
 sg13g2_decap_8 FILLER_0_19_819 ();
 sg13g2_decap_8 FILLER_0_19_826 ();
 sg13g2_decap_8 FILLER_0_19_833 ();
 sg13g2_decap_8 FILLER_0_19_840 ();
 sg13g2_decap_8 FILLER_0_19_847 ();
 sg13g2_decap_8 FILLER_0_19_854 ();
 sg13g2_decap_8 FILLER_0_19_861 ();
 sg13g2_decap_8 FILLER_0_19_868 ();
 sg13g2_decap_8 FILLER_0_19_875 ();
 sg13g2_decap_8 FILLER_0_19_882 ();
 sg13g2_decap_8 FILLER_0_19_889 ();
 sg13g2_decap_8 FILLER_0_19_896 ();
 sg13g2_decap_8 FILLER_0_19_903 ();
 sg13g2_decap_8 FILLER_0_19_910 ();
 sg13g2_decap_8 FILLER_0_19_917 ();
 sg13g2_decap_8 FILLER_0_19_924 ();
 sg13g2_decap_8 FILLER_0_19_931 ();
 sg13g2_decap_8 FILLER_0_19_938 ();
 sg13g2_decap_8 FILLER_0_19_945 ();
 sg13g2_decap_8 FILLER_0_19_952 ();
 sg13g2_decap_8 FILLER_0_19_959 ();
 sg13g2_decap_8 FILLER_0_19_966 ();
 sg13g2_decap_8 FILLER_0_19_973 ();
 sg13g2_decap_8 FILLER_0_19_980 ();
 sg13g2_decap_8 FILLER_0_19_987 ();
 sg13g2_decap_8 FILLER_0_19_994 ();
 sg13g2_decap_8 FILLER_0_19_1001 ();
 sg13g2_decap_8 FILLER_0_19_1008 ();
 sg13g2_decap_8 FILLER_0_19_1015 ();
 sg13g2_decap_8 FILLER_0_19_1022 ();
 sg13g2_decap_8 FILLER_0_19_1029 ();
 sg13g2_decap_8 FILLER_0_19_1036 ();
 sg13g2_decap_8 FILLER_0_19_1043 ();
 sg13g2_decap_8 FILLER_0_19_1050 ();
 sg13g2_decap_8 FILLER_0_19_1057 ();
 sg13g2_decap_8 FILLER_0_19_1064 ();
 sg13g2_decap_8 FILLER_0_19_1071 ();
 sg13g2_decap_8 FILLER_0_19_1078 ();
 sg13g2_decap_8 FILLER_0_19_1085 ();
 sg13g2_decap_8 FILLER_0_19_1092 ();
 sg13g2_decap_8 FILLER_0_19_1099 ();
 sg13g2_decap_8 FILLER_0_19_1106 ();
 sg13g2_decap_8 FILLER_0_19_1113 ();
 sg13g2_decap_8 FILLER_0_19_1120 ();
 sg13g2_decap_8 FILLER_0_19_1127 ();
 sg13g2_decap_8 FILLER_0_19_1134 ();
 sg13g2_decap_8 FILLER_0_19_1141 ();
 sg13g2_decap_8 FILLER_0_19_1148 ();
 sg13g2_decap_8 FILLER_0_19_1155 ();
 sg13g2_decap_8 FILLER_0_19_1162 ();
 sg13g2_decap_8 FILLER_0_19_1169 ();
 sg13g2_decap_8 FILLER_0_19_1176 ();
 sg13g2_decap_8 FILLER_0_19_1183 ();
 sg13g2_decap_8 FILLER_0_19_1190 ();
 sg13g2_decap_8 FILLER_0_19_1197 ();
 sg13g2_decap_8 FILLER_0_19_1204 ();
 sg13g2_decap_8 FILLER_0_19_1211 ();
 sg13g2_decap_8 FILLER_0_19_1218 ();
 sg13g2_fill_2 FILLER_0_19_1225 ();
 sg13g2_fill_1 FILLER_0_19_1227 ();
 sg13g2_decap_8 FILLER_0_20_0 ();
 sg13g2_decap_8 FILLER_0_20_7 ();
 sg13g2_decap_8 FILLER_0_20_14 ();
 sg13g2_decap_8 FILLER_0_20_21 ();
 sg13g2_decap_8 FILLER_0_20_28 ();
 sg13g2_decap_8 FILLER_0_20_35 ();
 sg13g2_decap_8 FILLER_0_20_42 ();
 sg13g2_decap_8 FILLER_0_20_49 ();
 sg13g2_decap_8 FILLER_0_20_56 ();
 sg13g2_decap_8 FILLER_0_20_63 ();
 sg13g2_decap_8 FILLER_0_20_70 ();
 sg13g2_decap_8 FILLER_0_20_77 ();
 sg13g2_decap_8 FILLER_0_20_84 ();
 sg13g2_decap_8 FILLER_0_20_91 ();
 sg13g2_decap_8 FILLER_0_20_98 ();
 sg13g2_decap_8 FILLER_0_20_105 ();
 sg13g2_decap_8 FILLER_0_20_112 ();
 sg13g2_decap_8 FILLER_0_20_119 ();
 sg13g2_decap_8 FILLER_0_20_126 ();
 sg13g2_decap_8 FILLER_0_20_133 ();
 sg13g2_decap_8 FILLER_0_20_140 ();
 sg13g2_decap_8 FILLER_0_20_147 ();
 sg13g2_decap_8 FILLER_0_20_154 ();
 sg13g2_decap_8 FILLER_0_20_161 ();
 sg13g2_decap_8 FILLER_0_20_168 ();
 sg13g2_decap_8 FILLER_0_20_175 ();
 sg13g2_decap_8 FILLER_0_20_182 ();
 sg13g2_decap_8 FILLER_0_20_189 ();
 sg13g2_decap_8 FILLER_0_20_196 ();
 sg13g2_decap_8 FILLER_0_20_203 ();
 sg13g2_decap_8 FILLER_0_20_210 ();
 sg13g2_decap_8 FILLER_0_20_217 ();
 sg13g2_decap_8 FILLER_0_20_224 ();
 sg13g2_decap_8 FILLER_0_20_231 ();
 sg13g2_decap_8 FILLER_0_20_238 ();
 sg13g2_decap_8 FILLER_0_20_245 ();
 sg13g2_decap_8 FILLER_0_20_252 ();
 sg13g2_decap_8 FILLER_0_20_259 ();
 sg13g2_decap_8 FILLER_0_20_266 ();
 sg13g2_decap_8 FILLER_0_20_273 ();
 sg13g2_decap_8 FILLER_0_20_280 ();
 sg13g2_decap_8 FILLER_0_20_287 ();
 sg13g2_decap_8 FILLER_0_20_294 ();
 sg13g2_decap_8 FILLER_0_20_301 ();
 sg13g2_decap_8 FILLER_0_20_308 ();
 sg13g2_decap_8 FILLER_0_20_315 ();
 sg13g2_decap_8 FILLER_0_20_322 ();
 sg13g2_decap_8 FILLER_0_20_329 ();
 sg13g2_decap_8 FILLER_0_20_336 ();
 sg13g2_decap_8 FILLER_0_20_343 ();
 sg13g2_decap_8 FILLER_0_20_350 ();
 sg13g2_decap_8 FILLER_0_20_357 ();
 sg13g2_decap_8 FILLER_0_20_364 ();
 sg13g2_decap_8 FILLER_0_20_371 ();
 sg13g2_decap_8 FILLER_0_20_378 ();
 sg13g2_decap_8 FILLER_0_20_385 ();
 sg13g2_decap_8 FILLER_0_20_392 ();
 sg13g2_decap_8 FILLER_0_20_399 ();
 sg13g2_decap_8 FILLER_0_20_406 ();
 sg13g2_decap_8 FILLER_0_20_413 ();
 sg13g2_decap_8 FILLER_0_20_420 ();
 sg13g2_decap_8 FILLER_0_20_427 ();
 sg13g2_decap_8 FILLER_0_20_434 ();
 sg13g2_decap_8 FILLER_0_20_441 ();
 sg13g2_decap_8 FILLER_0_20_448 ();
 sg13g2_decap_8 FILLER_0_20_455 ();
 sg13g2_decap_8 FILLER_0_20_462 ();
 sg13g2_decap_8 FILLER_0_20_469 ();
 sg13g2_decap_8 FILLER_0_20_476 ();
 sg13g2_decap_8 FILLER_0_20_483 ();
 sg13g2_decap_8 FILLER_0_20_490 ();
 sg13g2_decap_8 FILLER_0_20_497 ();
 sg13g2_decap_8 FILLER_0_20_504 ();
 sg13g2_decap_8 FILLER_0_20_511 ();
 sg13g2_decap_8 FILLER_0_20_518 ();
 sg13g2_decap_8 FILLER_0_20_525 ();
 sg13g2_decap_8 FILLER_0_20_532 ();
 sg13g2_decap_8 FILLER_0_20_539 ();
 sg13g2_decap_8 FILLER_0_20_546 ();
 sg13g2_decap_8 FILLER_0_20_553 ();
 sg13g2_decap_8 FILLER_0_20_560 ();
 sg13g2_decap_8 FILLER_0_20_567 ();
 sg13g2_decap_8 FILLER_0_20_574 ();
 sg13g2_decap_8 FILLER_0_20_581 ();
 sg13g2_decap_8 FILLER_0_20_588 ();
 sg13g2_decap_8 FILLER_0_20_595 ();
 sg13g2_decap_8 FILLER_0_20_602 ();
 sg13g2_decap_8 FILLER_0_20_609 ();
 sg13g2_decap_8 FILLER_0_20_616 ();
 sg13g2_decap_8 FILLER_0_20_623 ();
 sg13g2_decap_8 FILLER_0_20_630 ();
 sg13g2_decap_8 FILLER_0_20_637 ();
 sg13g2_decap_8 FILLER_0_20_644 ();
 sg13g2_decap_8 FILLER_0_20_651 ();
 sg13g2_decap_8 FILLER_0_20_658 ();
 sg13g2_decap_8 FILLER_0_20_665 ();
 sg13g2_decap_8 FILLER_0_20_672 ();
 sg13g2_decap_8 FILLER_0_20_679 ();
 sg13g2_decap_8 FILLER_0_20_686 ();
 sg13g2_decap_8 FILLER_0_20_693 ();
 sg13g2_decap_8 FILLER_0_20_700 ();
 sg13g2_decap_8 FILLER_0_20_707 ();
 sg13g2_decap_8 FILLER_0_20_714 ();
 sg13g2_decap_8 FILLER_0_20_721 ();
 sg13g2_decap_8 FILLER_0_20_728 ();
 sg13g2_decap_8 FILLER_0_20_735 ();
 sg13g2_decap_8 FILLER_0_20_742 ();
 sg13g2_decap_8 FILLER_0_20_749 ();
 sg13g2_decap_8 FILLER_0_20_756 ();
 sg13g2_decap_8 FILLER_0_20_763 ();
 sg13g2_decap_8 FILLER_0_20_770 ();
 sg13g2_decap_8 FILLER_0_20_777 ();
 sg13g2_decap_8 FILLER_0_20_784 ();
 sg13g2_decap_8 FILLER_0_20_791 ();
 sg13g2_decap_8 FILLER_0_20_798 ();
 sg13g2_decap_8 FILLER_0_20_805 ();
 sg13g2_decap_8 FILLER_0_20_812 ();
 sg13g2_decap_8 FILLER_0_20_819 ();
 sg13g2_decap_8 FILLER_0_20_826 ();
 sg13g2_decap_8 FILLER_0_20_833 ();
 sg13g2_decap_8 FILLER_0_20_840 ();
 sg13g2_decap_8 FILLER_0_20_847 ();
 sg13g2_decap_8 FILLER_0_20_854 ();
 sg13g2_decap_8 FILLER_0_20_861 ();
 sg13g2_decap_8 FILLER_0_20_868 ();
 sg13g2_decap_8 FILLER_0_20_875 ();
 sg13g2_decap_8 FILLER_0_20_882 ();
 sg13g2_decap_8 FILLER_0_20_889 ();
 sg13g2_decap_8 FILLER_0_20_896 ();
 sg13g2_decap_8 FILLER_0_20_903 ();
 sg13g2_decap_8 FILLER_0_20_910 ();
 sg13g2_decap_8 FILLER_0_20_917 ();
 sg13g2_decap_8 FILLER_0_20_924 ();
 sg13g2_decap_8 FILLER_0_20_931 ();
 sg13g2_decap_8 FILLER_0_20_938 ();
 sg13g2_decap_8 FILLER_0_20_945 ();
 sg13g2_decap_8 FILLER_0_20_952 ();
 sg13g2_decap_8 FILLER_0_20_959 ();
 sg13g2_decap_8 FILLER_0_20_966 ();
 sg13g2_decap_8 FILLER_0_20_973 ();
 sg13g2_decap_8 FILLER_0_20_980 ();
 sg13g2_decap_8 FILLER_0_20_987 ();
 sg13g2_decap_8 FILLER_0_20_994 ();
 sg13g2_decap_8 FILLER_0_20_1001 ();
 sg13g2_decap_8 FILLER_0_20_1008 ();
 sg13g2_decap_8 FILLER_0_20_1015 ();
 sg13g2_decap_8 FILLER_0_20_1022 ();
 sg13g2_decap_8 FILLER_0_20_1029 ();
 sg13g2_decap_8 FILLER_0_20_1036 ();
 sg13g2_decap_8 FILLER_0_20_1043 ();
 sg13g2_decap_8 FILLER_0_20_1050 ();
 sg13g2_decap_8 FILLER_0_20_1057 ();
 sg13g2_decap_8 FILLER_0_20_1064 ();
 sg13g2_decap_8 FILLER_0_20_1071 ();
 sg13g2_decap_8 FILLER_0_20_1078 ();
 sg13g2_decap_8 FILLER_0_20_1085 ();
 sg13g2_decap_8 FILLER_0_20_1092 ();
 sg13g2_decap_8 FILLER_0_20_1099 ();
 sg13g2_decap_8 FILLER_0_20_1106 ();
 sg13g2_decap_8 FILLER_0_20_1113 ();
 sg13g2_decap_8 FILLER_0_20_1120 ();
 sg13g2_decap_8 FILLER_0_20_1127 ();
 sg13g2_decap_8 FILLER_0_20_1134 ();
 sg13g2_decap_8 FILLER_0_20_1141 ();
 sg13g2_decap_8 FILLER_0_20_1148 ();
 sg13g2_decap_8 FILLER_0_20_1155 ();
 sg13g2_decap_8 FILLER_0_20_1162 ();
 sg13g2_decap_8 FILLER_0_20_1169 ();
 sg13g2_decap_8 FILLER_0_20_1176 ();
 sg13g2_decap_8 FILLER_0_20_1183 ();
 sg13g2_decap_8 FILLER_0_20_1190 ();
 sg13g2_decap_8 FILLER_0_20_1197 ();
 sg13g2_decap_8 FILLER_0_20_1204 ();
 sg13g2_decap_8 FILLER_0_20_1211 ();
 sg13g2_decap_8 FILLER_0_20_1218 ();
 sg13g2_fill_2 FILLER_0_20_1225 ();
 sg13g2_fill_1 FILLER_0_20_1227 ();
 sg13g2_decap_8 FILLER_0_21_0 ();
 sg13g2_decap_8 FILLER_0_21_7 ();
 sg13g2_decap_8 FILLER_0_21_14 ();
 sg13g2_decap_8 FILLER_0_21_21 ();
 sg13g2_decap_8 FILLER_0_21_28 ();
 sg13g2_decap_8 FILLER_0_21_35 ();
 sg13g2_decap_8 FILLER_0_21_42 ();
 sg13g2_decap_8 FILLER_0_21_49 ();
 sg13g2_decap_8 FILLER_0_21_56 ();
 sg13g2_decap_8 FILLER_0_21_63 ();
 sg13g2_decap_8 FILLER_0_21_70 ();
 sg13g2_decap_8 FILLER_0_21_77 ();
 sg13g2_decap_8 FILLER_0_21_84 ();
 sg13g2_decap_8 FILLER_0_21_91 ();
 sg13g2_decap_8 FILLER_0_21_98 ();
 sg13g2_decap_8 FILLER_0_21_105 ();
 sg13g2_decap_8 FILLER_0_21_112 ();
 sg13g2_decap_8 FILLER_0_21_119 ();
 sg13g2_decap_8 FILLER_0_21_126 ();
 sg13g2_decap_8 FILLER_0_21_133 ();
 sg13g2_decap_8 FILLER_0_21_140 ();
 sg13g2_decap_8 FILLER_0_21_147 ();
 sg13g2_decap_8 FILLER_0_21_154 ();
 sg13g2_decap_8 FILLER_0_21_161 ();
 sg13g2_decap_8 FILLER_0_21_168 ();
 sg13g2_decap_8 FILLER_0_21_175 ();
 sg13g2_decap_8 FILLER_0_21_182 ();
 sg13g2_decap_8 FILLER_0_21_189 ();
 sg13g2_decap_8 FILLER_0_21_196 ();
 sg13g2_decap_8 FILLER_0_21_203 ();
 sg13g2_decap_8 FILLER_0_21_210 ();
 sg13g2_decap_8 FILLER_0_21_217 ();
 sg13g2_decap_8 FILLER_0_21_224 ();
 sg13g2_decap_8 FILLER_0_21_231 ();
 sg13g2_decap_8 FILLER_0_21_238 ();
 sg13g2_decap_8 FILLER_0_21_245 ();
 sg13g2_decap_8 FILLER_0_21_252 ();
 sg13g2_decap_8 FILLER_0_21_259 ();
 sg13g2_decap_8 FILLER_0_21_266 ();
 sg13g2_decap_8 FILLER_0_21_273 ();
 sg13g2_decap_8 FILLER_0_21_280 ();
 sg13g2_decap_8 FILLER_0_21_287 ();
 sg13g2_decap_8 FILLER_0_21_294 ();
 sg13g2_decap_8 FILLER_0_21_301 ();
 sg13g2_decap_8 FILLER_0_21_308 ();
 sg13g2_decap_8 FILLER_0_21_315 ();
 sg13g2_decap_8 FILLER_0_21_322 ();
 sg13g2_decap_8 FILLER_0_21_329 ();
 sg13g2_decap_8 FILLER_0_21_336 ();
 sg13g2_decap_8 FILLER_0_21_343 ();
 sg13g2_decap_8 FILLER_0_21_350 ();
 sg13g2_decap_8 FILLER_0_21_357 ();
 sg13g2_decap_8 FILLER_0_21_364 ();
 sg13g2_decap_8 FILLER_0_21_371 ();
 sg13g2_decap_8 FILLER_0_21_378 ();
 sg13g2_decap_8 FILLER_0_21_385 ();
 sg13g2_decap_8 FILLER_0_21_392 ();
 sg13g2_decap_8 FILLER_0_21_399 ();
 sg13g2_decap_8 FILLER_0_21_406 ();
 sg13g2_decap_8 FILLER_0_21_413 ();
 sg13g2_decap_8 FILLER_0_21_420 ();
 sg13g2_decap_8 FILLER_0_21_427 ();
 sg13g2_decap_8 FILLER_0_21_434 ();
 sg13g2_decap_8 FILLER_0_21_441 ();
 sg13g2_decap_8 FILLER_0_21_448 ();
 sg13g2_decap_8 FILLER_0_21_455 ();
 sg13g2_decap_8 FILLER_0_21_462 ();
 sg13g2_decap_8 FILLER_0_21_469 ();
 sg13g2_decap_8 FILLER_0_21_476 ();
 sg13g2_decap_8 FILLER_0_21_483 ();
 sg13g2_decap_8 FILLER_0_21_490 ();
 sg13g2_decap_8 FILLER_0_21_497 ();
 sg13g2_decap_8 FILLER_0_21_504 ();
 sg13g2_decap_8 FILLER_0_21_511 ();
 sg13g2_decap_8 FILLER_0_21_518 ();
 sg13g2_decap_8 FILLER_0_21_525 ();
 sg13g2_decap_8 FILLER_0_21_532 ();
 sg13g2_decap_8 FILLER_0_21_539 ();
 sg13g2_decap_8 FILLER_0_21_546 ();
 sg13g2_decap_8 FILLER_0_21_553 ();
 sg13g2_decap_8 FILLER_0_21_560 ();
 sg13g2_decap_8 FILLER_0_21_567 ();
 sg13g2_decap_8 FILLER_0_21_574 ();
 sg13g2_decap_8 FILLER_0_21_581 ();
 sg13g2_decap_8 FILLER_0_21_588 ();
 sg13g2_decap_8 FILLER_0_21_595 ();
 sg13g2_decap_8 FILLER_0_21_602 ();
 sg13g2_decap_8 FILLER_0_21_609 ();
 sg13g2_decap_8 FILLER_0_21_616 ();
 sg13g2_decap_8 FILLER_0_21_623 ();
 sg13g2_decap_8 FILLER_0_21_630 ();
 sg13g2_decap_8 FILLER_0_21_637 ();
 sg13g2_decap_8 FILLER_0_21_644 ();
 sg13g2_decap_8 FILLER_0_21_651 ();
 sg13g2_decap_8 FILLER_0_21_658 ();
 sg13g2_decap_8 FILLER_0_21_665 ();
 sg13g2_decap_8 FILLER_0_21_672 ();
 sg13g2_decap_8 FILLER_0_21_679 ();
 sg13g2_decap_8 FILLER_0_21_686 ();
 sg13g2_decap_8 FILLER_0_21_693 ();
 sg13g2_decap_8 FILLER_0_21_700 ();
 sg13g2_decap_8 FILLER_0_21_707 ();
 sg13g2_decap_8 FILLER_0_21_714 ();
 sg13g2_decap_8 FILLER_0_21_721 ();
 sg13g2_decap_8 FILLER_0_21_728 ();
 sg13g2_decap_8 FILLER_0_21_735 ();
 sg13g2_decap_8 FILLER_0_21_742 ();
 sg13g2_decap_8 FILLER_0_21_749 ();
 sg13g2_decap_8 FILLER_0_21_756 ();
 sg13g2_decap_8 FILLER_0_21_763 ();
 sg13g2_decap_8 FILLER_0_21_770 ();
 sg13g2_decap_8 FILLER_0_21_777 ();
 sg13g2_decap_8 FILLER_0_21_784 ();
 sg13g2_decap_8 FILLER_0_21_791 ();
 sg13g2_decap_8 FILLER_0_21_798 ();
 sg13g2_decap_8 FILLER_0_21_805 ();
 sg13g2_decap_8 FILLER_0_21_812 ();
 sg13g2_decap_8 FILLER_0_21_819 ();
 sg13g2_decap_8 FILLER_0_21_826 ();
 sg13g2_decap_8 FILLER_0_21_833 ();
 sg13g2_decap_8 FILLER_0_21_840 ();
 sg13g2_decap_8 FILLER_0_21_847 ();
 sg13g2_decap_8 FILLER_0_21_854 ();
 sg13g2_decap_8 FILLER_0_21_861 ();
 sg13g2_decap_8 FILLER_0_21_868 ();
 sg13g2_decap_8 FILLER_0_21_875 ();
 sg13g2_decap_8 FILLER_0_21_882 ();
 sg13g2_decap_8 FILLER_0_21_889 ();
 sg13g2_decap_8 FILLER_0_21_896 ();
 sg13g2_decap_8 FILLER_0_21_903 ();
 sg13g2_decap_8 FILLER_0_21_910 ();
 sg13g2_decap_8 FILLER_0_21_917 ();
 sg13g2_decap_8 FILLER_0_21_924 ();
 sg13g2_decap_8 FILLER_0_21_931 ();
 sg13g2_decap_8 FILLER_0_21_938 ();
 sg13g2_decap_8 FILLER_0_21_945 ();
 sg13g2_decap_8 FILLER_0_21_952 ();
 sg13g2_decap_8 FILLER_0_21_959 ();
 sg13g2_decap_8 FILLER_0_21_966 ();
 sg13g2_decap_8 FILLER_0_21_973 ();
 sg13g2_decap_8 FILLER_0_21_980 ();
 sg13g2_decap_8 FILLER_0_21_987 ();
 sg13g2_decap_8 FILLER_0_21_994 ();
 sg13g2_decap_8 FILLER_0_21_1001 ();
 sg13g2_decap_8 FILLER_0_21_1008 ();
 sg13g2_decap_8 FILLER_0_21_1015 ();
 sg13g2_decap_8 FILLER_0_21_1022 ();
 sg13g2_decap_8 FILLER_0_21_1029 ();
 sg13g2_decap_8 FILLER_0_21_1036 ();
 sg13g2_decap_8 FILLER_0_21_1043 ();
 sg13g2_decap_8 FILLER_0_21_1050 ();
 sg13g2_decap_8 FILLER_0_21_1057 ();
 sg13g2_decap_8 FILLER_0_21_1064 ();
 sg13g2_decap_8 FILLER_0_21_1071 ();
 sg13g2_decap_8 FILLER_0_21_1078 ();
 sg13g2_decap_8 FILLER_0_21_1085 ();
 sg13g2_decap_8 FILLER_0_21_1092 ();
 sg13g2_decap_8 FILLER_0_21_1099 ();
 sg13g2_decap_8 FILLER_0_21_1106 ();
 sg13g2_decap_8 FILLER_0_21_1113 ();
 sg13g2_decap_8 FILLER_0_21_1120 ();
 sg13g2_decap_8 FILLER_0_21_1127 ();
 sg13g2_decap_8 FILLER_0_21_1134 ();
 sg13g2_decap_8 FILLER_0_21_1141 ();
 sg13g2_decap_8 FILLER_0_21_1148 ();
 sg13g2_decap_8 FILLER_0_21_1155 ();
 sg13g2_decap_8 FILLER_0_21_1162 ();
 sg13g2_decap_8 FILLER_0_21_1169 ();
 sg13g2_decap_8 FILLER_0_21_1176 ();
 sg13g2_decap_8 FILLER_0_21_1183 ();
 sg13g2_decap_8 FILLER_0_21_1190 ();
 sg13g2_decap_8 FILLER_0_21_1197 ();
 sg13g2_decap_8 FILLER_0_21_1204 ();
 sg13g2_decap_8 FILLER_0_21_1211 ();
 sg13g2_decap_8 FILLER_0_21_1218 ();
 sg13g2_fill_2 FILLER_0_21_1225 ();
 sg13g2_fill_1 FILLER_0_21_1227 ();
 sg13g2_decap_8 FILLER_0_22_0 ();
 sg13g2_decap_8 FILLER_0_22_7 ();
 sg13g2_decap_8 FILLER_0_22_14 ();
 sg13g2_decap_8 FILLER_0_22_21 ();
 sg13g2_decap_8 FILLER_0_22_28 ();
 sg13g2_decap_8 FILLER_0_22_35 ();
 sg13g2_decap_8 FILLER_0_22_42 ();
 sg13g2_decap_8 FILLER_0_22_49 ();
 sg13g2_decap_8 FILLER_0_22_56 ();
 sg13g2_decap_8 FILLER_0_22_63 ();
 sg13g2_decap_8 FILLER_0_22_70 ();
 sg13g2_decap_8 FILLER_0_22_77 ();
 sg13g2_decap_8 FILLER_0_22_84 ();
 sg13g2_decap_8 FILLER_0_22_91 ();
 sg13g2_decap_8 FILLER_0_22_98 ();
 sg13g2_decap_8 FILLER_0_22_105 ();
 sg13g2_decap_8 FILLER_0_22_112 ();
 sg13g2_decap_8 FILLER_0_22_119 ();
 sg13g2_decap_8 FILLER_0_22_126 ();
 sg13g2_decap_8 FILLER_0_22_133 ();
 sg13g2_decap_8 FILLER_0_22_140 ();
 sg13g2_decap_8 FILLER_0_22_147 ();
 sg13g2_decap_8 FILLER_0_22_154 ();
 sg13g2_decap_8 FILLER_0_22_161 ();
 sg13g2_decap_8 FILLER_0_22_168 ();
 sg13g2_decap_8 FILLER_0_22_175 ();
 sg13g2_decap_8 FILLER_0_22_182 ();
 sg13g2_decap_8 FILLER_0_22_189 ();
 sg13g2_decap_8 FILLER_0_22_196 ();
 sg13g2_decap_8 FILLER_0_22_203 ();
 sg13g2_decap_8 FILLER_0_22_210 ();
 sg13g2_decap_8 FILLER_0_22_217 ();
 sg13g2_decap_8 FILLER_0_22_224 ();
 sg13g2_decap_8 FILLER_0_22_231 ();
 sg13g2_decap_8 FILLER_0_22_238 ();
 sg13g2_decap_8 FILLER_0_22_245 ();
 sg13g2_decap_8 FILLER_0_22_252 ();
 sg13g2_decap_8 FILLER_0_22_259 ();
 sg13g2_decap_8 FILLER_0_22_266 ();
 sg13g2_decap_8 FILLER_0_22_273 ();
 sg13g2_decap_8 FILLER_0_22_280 ();
 sg13g2_decap_8 FILLER_0_22_287 ();
 sg13g2_decap_8 FILLER_0_22_294 ();
 sg13g2_decap_8 FILLER_0_22_301 ();
 sg13g2_decap_8 FILLER_0_22_308 ();
 sg13g2_decap_8 FILLER_0_22_315 ();
 sg13g2_decap_8 FILLER_0_22_322 ();
 sg13g2_decap_8 FILLER_0_22_329 ();
 sg13g2_decap_8 FILLER_0_22_336 ();
 sg13g2_decap_8 FILLER_0_22_343 ();
 sg13g2_decap_8 FILLER_0_22_350 ();
 sg13g2_decap_8 FILLER_0_22_357 ();
 sg13g2_decap_8 FILLER_0_22_364 ();
 sg13g2_decap_8 FILLER_0_22_371 ();
 sg13g2_decap_8 FILLER_0_22_378 ();
 sg13g2_decap_8 FILLER_0_22_385 ();
 sg13g2_decap_8 FILLER_0_22_392 ();
 sg13g2_decap_8 FILLER_0_22_399 ();
 sg13g2_fill_2 FILLER_0_22_406 ();
 sg13g2_decap_4 FILLER_0_22_413 ();
 sg13g2_decap_8 FILLER_0_22_426 ();
 sg13g2_decap_8 FILLER_0_22_433 ();
 sg13g2_decap_8 FILLER_0_22_440 ();
 sg13g2_decap_8 FILLER_0_22_447 ();
 sg13g2_decap_8 FILLER_0_22_454 ();
 sg13g2_decap_8 FILLER_0_22_461 ();
 sg13g2_decap_8 FILLER_0_22_468 ();
 sg13g2_decap_8 FILLER_0_22_475 ();
 sg13g2_decap_8 FILLER_0_22_482 ();
 sg13g2_decap_4 FILLER_0_22_489 ();
 sg13g2_fill_2 FILLER_0_22_493 ();
 sg13g2_decap_8 FILLER_0_22_499 ();
 sg13g2_decap_4 FILLER_0_22_506 ();
 sg13g2_decap_8 FILLER_0_22_515 ();
 sg13g2_decap_8 FILLER_0_22_522 ();
 sg13g2_decap_8 FILLER_0_22_529 ();
 sg13g2_decap_8 FILLER_0_22_536 ();
 sg13g2_decap_8 FILLER_0_22_543 ();
 sg13g2_decap_8 FILLER_0_22_550 ();
 sg13g2_decap_8 FILLER_0_22_557 ();
 sg13g2_decap_8 FILLER_0_22_564 ();
 sg13g2_decap_8 FILLER_0_22_571 ();
 sg13g2_decap_8 FILLER_0_22_578 ();
 sg13g2_decap_8 FILLER_0_22_585 ();
 sg13g2_decap_8 FILLER_0_22_592 ();
 sg13g2_decap_8 FILLER_0_22_599 ();
 sg13g2_decap_8 FILLER_0_22_606 ();
 sg13g2_decap_8 FILLER_0_22_613 ();
 sg13g2_decap_8 FILLER_0_22_620 ();
 sg13g2_decap_8 FILLER_0_22_627 ();
 sg13g2_decap_8 FILLER_0_22_634 ();
 sg13g2_decap_8 FILLER_0_22_641 ();
 sg13g2_decap_8 FILLER_0_22_648 ();
 sg13g2_decap_8 FILLER_0_22_655 ();
 sg13g2_decap_8 FILLER_0_22_662 ();
 sg13g2_decap_8 FILLER_0_22_669 ();
 sg13g2_decap_8 FILLER_0_22_676 ();
 sg13g2_decap_8 FILLER_0_22_683 ();
 sg13g2_decap_8 FILLER_0_22_690 ();
 sg13g2_decap_8 FILLER_0_22_697 ();
 sg13g2_decap_8 FILLER_0_22_704 ();
 sg13g2_decap_8 FILLER_0_22_711 ();
 sg13g2_decap_8 FILLER_0_22_718 ();
 sg13g2_decap_8 FILLER_0_22_725 ();
 sg13g2_decap_8 FILLER_0_22_732 ();
 sg13g2_decap_8 FILLER_0_22_739 ();
 sg13g2_decap_8 FILLER_0_22_746 ();
 sg13g2_decap_8 FILLER_0_22_753 ();
 sg13g2_decap_8 FILLER_0_22_760 ();
 sg13g2_decap_8 FILLER_0_22_767 ();
 sg13g2_decap_8 FILLER_0_22_774 ();
 sg13g2_decap_8 FILLER_0_22_781 ();
 sg13g2_decap_8 FILLER_0_22_788 ();
 sg13g2_decap_8 FILLER_0_22_795 ();
 sg13g2_decap_8 FILLER_0_22_802 ();
 sg13g2_decap_8 FILLER_0_22_809 ();
 sg13g2_decap_8 FILLER_0_22_816 ();
 sg13g2_decap_8 FILLER_0_22_823 ();
 sg13g2_decap_8 FILLER_0_22_830 ();
 sg13g2_decap_8 FILLER_0_22_837 ();
 sg13g2_decap_8 FILLER_0_22_844 ();
 sg13g2_decap_8 FILLER_0_22_851 ();
 sg13g2_decap_8 FILLER_0_22_858 ();
 sg13g2_decap_8 FILLER_0_22_865 ();
 sg13g2_decap_8 FILLER_0_22_872 ();
 sg13g2_decap_8 FILLER_0_22_879 ();
 sg13g2_decap_8 FILLER_0_22_886 ();
 sg13g2_decap_8 FILLER_0_22_893 ();
 sg13g2_decap_8 FILLER_0_22_900 ();
 sg13g2_decap_8 FILLER_0_22_907 ();
 sg13g2_decap_8 FILLER_0_22_914 ();
 sg13g2_decap_8 FILLER_0_22_921 ();
 sg13g2_decap_8 FILLER_0_22_928 ();
 sg13g2_decap_8 FILLER_0_22_935 ();
 sg13g2_decap_8 FILLER_0_22_942 ();
 sg13g2_decap_8 FILLER_0_22_949 ();
 sg13g2_decap_8 FILLER_0_22_956 ();
 sg13g2_decap_8 FILLER_0_22_963 ();
 sg13g2_decap_8 FILLER_0_22_970 ();
 sg13g2_decap_8 FILLER_0_22_977 ();
 sg13g2_decap_8 FILLER_0_22_984 ();
 sg13g2_decap_8 FILLER_0_22_991 ();
 sg13g2_decap_8 FILLER_0_22_998 ();
 sg13g2_decap_8 FILLER_0_22_1005 ();
 sg13g2_decap_8 FILLER_0_22_1012 ();
 sg13g2_decap_8 FILLER_0_22_1019 ();
 sg13g2_decap_8 FILLER_0_22_1026 ();
 sg13g2_decap_8 FILLER_0_22_1033 ();
 sg13g2_decap_8 FILLER_0_22_1040 ();
 sg13g2_decap_8 FILLER_0_22_1047 ();
 sg13g2_decap_8 FILLER_0_22_1054 ();
 sg13g2_decap_8 FILLER_0_22_1061 ();
 sg13g2_decap_8 FILLER_0_22_1068 ();
 sg13g2_decap_8 FILLER_0_22_1075 ();
 sg13g2_decap_8 FILLER_0_22_1082 ();
 sg13g2_decap_8 FILLER_0_22_1089 ();
 sg13g2_decap_8 FILLER_0_22_1096 ();
 sg13g2_decap_8 FILLER_0_22_1103 ();
 sg13g2_decap_8 FILLER_0_22_1110 ();
 sg13g2_decap_8 FILLER_0_22_1117 ();
 sg13g2_decap_8 FILLER_0_22_1124 ();
 sg13g2_decap_8 FILLER_0_22_1131 ();
 sg13g2_decap_8 FILLER_0_22_1138 ();
 sg13g2_decap_8 FILLER_0_22_1145 ();
 sg13g2_decap_8 FILLER_0_22_1152 ();
 sg13g2_decap_8 FILLER_0_22_1159 ();
 sg13g2_decap_8 FILLER_0_22_1166 ();
 sg13g2_decap_8 FILLER_0_22_1173 ();
 sg13g2_decap_8 FILLER_0_22_1180 ();
 sg13g2_decap_8 FILLER_0_22_1187 ();
 sg13g2_decap_8 FILLER_0_22_1194 ();
 sg13g2_decap_8 FILLER_0_22_1201 ();
 sg13g2_decap_8 FILLER_0_22_1208 ();
 sg13g2_decap_8 FILLER_0_22_1215 ();
 sg13g2_decap_4 FILLER_0_22_1222 ();
 sg13g2_fill_2 FILLER_0_22_1226 ();
 sg13g2_decap_8 FILLER_0_23_0 ();
 sg13g2_decap_8 FILLER_0_23_7 ();
 sg13g2_decap_8 FILLER_0_23_14 ();
 sg13g2_decap_8 FILLER_0_23_21 ();
 sg13g2_fill_1 FILLER_0_23_28 ();
 sg13g2_decap_4 FILLER_0_23_33 ();
 sg13g2_fill_1 FILLER_0_23_37 ();
 sg13g2_decap_8 FILLER_0_23_42 ();
 sg13g2_fill_1 FILLER_0_23_49 ();
 sg13g2_decap_8 FILLER_0_23_55 ();
 sg13g2_decap_8 FILLER_0_23_62 ();
 sg13g2_decap_8 FILLER_0_23_69 ();
 sg13g2_decap_8 FILLER_0_23_76 ();
 sg13g2_decap_8 FILLER_0_23_83 ();
 sg13g2_decap_8 FILLER_0_23_90 ();
 sg13g2_decap_8 FILLER_0_23_97 ();
 sg13g2_decap_8 FILLER_0_23_104 ();
 sg13g2_decap_8 FILLER_0_23_111 ();
 sg13g2_decap_8 FILLER_0_23_118 ();
 sg13g2_decap_8 FILLER_0_23_125 ();
 sg13g2_decap_8 FILLER_0_23_132 ();
 sg13g2_decap_8 FILLER_0_23_139 ();
 sg13g2_decap_8 FILLER_0_23_146 ();
 sg13g2_decap_8 FILLER_0_23_153 ();
 sg13g2_decap_8 FILLER_0_23_160 ();
 sg13g2_decap_8 FILLER_0_23_167 ();
 sg13g2_decap_8 FILLER_0_23_174 ();
 sg13g2_decap_8 FILLER_0_23_181 ();
 sg13g2_decap_8 FILLER_0_23_188 ();
 sg13g2_decap_8 FILLER_0_23_195 ();
 sg13g2_decap_8 FILLER_0_23_202 ();
 sg13g2_decap_8 FILLER_0_23_209 ();
 sg13g2_decap_8 FILLER_0_23_216 ();
 sg13g2_decap_8 FILLER_0_23_223 ();
 sg13g2_decap_8 FILLER_0_23_230 ();
 sg13g2_decap_8 FILLER_0_23_237 ();
 sg13g2_decap_8 FILLER_0_23_244 ();
 sg13g2_decap_8 FILLER_0_23_251 ();
 sg13g2_decap_8 FILLER_0_23_258 ();
 sg13g2_decap_8 FILLER_0_23_265 ();
 sg13g2_decap_8 FILLER_0_23_272 ();
 sg13g2_decap_8 FILLER_0_23_279 ();
 sg13g2_decap_4 FILLER_0_23_290 ();
 sg13g2_fill_1 FILLER_0_23_294 ();
 sg13g2_decap_8 FILLER_0_23_321 ();
 sg13g2_decap_8 FILLER_0_23_328 ();
 sg13g2_fill_2 FILLER_0_23_335 ();
 sg13g2_fill_1 FILLER_0_23_337 ();
 sg13g2_decap_4 FILLER_0_23_343 ();
 sg13g2_fill_1 FILLER_0_23_347 ();
 sg13g2_decap_8 FILLER_0_23_353 ();
 sg13g2_decap_8 FILLER_0_23_360 ();
 sg13g2_decap_8 FILLER_0_23_367 ();
 sg13g2_decap_4 FILLER_0_23_374 ();
 sg13g2_fill_2 FILLER_0_23_378 ();
 sg13g2_decap_4 FILLER_0_23_385 ();
 sg13g2_fill_2 FILLER_0_23_389 ();
 sg13g2_decap_4 FILLER_0_23_406 ();
 sg13g2_decap_8 FILLER_0_23_436 ();
 sg13g2_decap_8 FILLER_0_23_443 ();
 sg13g2_decap_8 FILLER_0_23_450 ();
 sg13g2_decap_8 FILLER_0_23_457 ();
 sg13g2_decap_8 FILLER_0_23_464 ();
 sg13g2_fill_2 FILLER_0_23_471 ();
 sg13g2_fill_1 FILLER_0_23_473 ();
 sg13g2_fill_2 FILLER_0_23_514 ();
 sg13g2_fill_1 FILLER_0_23_516 ();
 sg13g2_decap_8 FILLER_0_23_548 ();
 sg13g2_decap_8 FILLER_0_23_555 ();
 sg13g2_decap_8 FILLER_0_23_562 ();
 sg13g2_decap_8 FILLER_0_23_569 ();
 sg13g2_decap_8 FILLER_0_23_576 ();
 sg13g2_decap_8 FILLER_0_23_583 ();
 sg13g2_decap_8 FILLER_0_23_590 ();
 sg13g2_decap_8 FILLER_0_23_597 ();
 sg13g2_decap_8 FILLER_0_23_604 ();
 sg13g2_decap_8 FILLER_0_23_611 ();
 sg13g2_decap_8 FILLER_0_23_618 ();
 sg13g2_decap_8 FILLER_0_23_625 ();
 sg13g2_decap_8 FILLER_0_23_632 ();
 sg13g2_decap_8 FILLER_0_23_639 ();
 sg13g2_decap_8 FILLER_0_23_646 ();
 sg13g2_decap_8 FILLER_0_23_653 ();
 sg13g2_decap_8 FILLER_0_23_660 ();
 sg13g2_decap_8 FILLER_0_23_667 ();
 sg13g2_decap_8 FILLER_0_23_674 ();
 sg13g2_decap_8 FILLER_0_23_681 ();
 sg13g2_decap_8 FILLER_0_23_688 ();
 sg13g2_decap_8 FILLER_0_23_695 ();
 sg13g2_decap_8 FILLER_0_23_702 ();
 sg13g2_decap_8 FILLER_0_23_709 ();
 sg13g2_decap_8 FILLER_0_23_716 ();
 sg13g2_decap_8 FILLER_0_23_723 ();
 sg13g2_decap_8 FILLER_0_23_730 ();
 sg13g2_decap_8 FILLER_0_23_737 ();
 sg13g2_decap_8 FILLER_0_23_744 ();
 sg13g2_decap_8 FILLER_0_23_751 ();
 sg13g2_decap_8 FILLER_0_23_758 ();
 sg13g2_decap_8 FILLER_0_23_765 ();
 sg13g2_decap_8 FILLER_0_23_772 ();
 sg13g2_decap_8 FILLER_0_23_779 ();
 sg13g2_decap_8 FILLER_0_23_786 ();
 sg13g2_decap_8 FILLER_0_23_793 ();
 sg13g2_decap_8 FILLER_0_23_800 ();
 sg13g2_decap_8 FILLER_0_23_807 ();
 sg13g2_decap_8 FILLER_0_23_814 ();
 sg13g2_decap_8 FILLER_0_23_821 ();
 sg13g2_decap_8 FILLER_0_23_828 ();
 sg13g2_decap_8 FILLER_0_23_835 ();
 sg13g2_decap_8 FILLER_0_23_842 ();
 sg13g2_decap_8 FILLER_0_23_849 ();
 sg13g2_decap_8 FILLER_0_23_856 ();
 sg13g2_decap_8 FILLER_0_23_863 ();
 sg13g2_decap_8 FILLER_0_23_870 ();
 sg13g2_decap_8 FILLER_0_23_877 ();
 sg13g2_decap_8 FILLER_0_23_884 ();
 sg13g2_decap_8 FILLER_0_23_891 ();
 sg13g2_decap_8 FILLER_0_23_898 ();
 sg13g2_decap_8 FILLER_0_23_905 ();
 sg13g2_decap_8 FILLER_0_23_912 ();
 sg13g2_decap_8 FILLER_0_23_919 ();
 sg13g2_decap_8 FILLER_0_23_926 ();
 sg13g2_decap_8 FILLER_0_23_933 ();
 sg13g2_decap_8 FILLER_0_23_940 ();
 sg13g2_decap_8 FILLER_0_23_947 ();
 sg13g2_decap_8 FILLER_0_23_954 ();
 sg13g2_decap_8 FILLER_0_23_961 ();
 sg13g2_decap_8 FILLER_0_23_968 ();
 sg13g2_decap_8 FILLER_0_23_975 ();
 sg13g2_decap_8 FILLER_0_23_982 ();
 sg13g2_decap_8 FILLER_0_23_989 ();
 sg13g2_decap_8 FILLER_0_23_996 ();
 sg13g2_decap_8 FILLER_0_23_1003 ();
 sg13g2_decap_8 FILLER_0_23_1010 ();
 sg13g2_decap_8 FILLER_0_23_1017 ();
 sg13g2_decap_8 FILLER_0_23_1029 ();
 sg13g2_decap_8 FILLER_0_23_1036 ();
 sg13g2_fill_2 FILLER_0_23_1043 ();
 sg13g2_decap_4 FILLER_0_23_1071 ();
 sg13g2_fill_2 FILLER_0_23_1075 ();
 sg13g2_decap_8 FILLER_0_23_1103 ();
 sg13g2_decap_8 FILLER_0_23_1110 ();
 sg13g2_decap_8 FILLER_0_23_1117 ();
 sg13g2_decap_8 FILLER_0_23_1124 ();
 sg13g2_decap_8 FILLER_0_23_1131 ();
 sg13g2_decap_8 FILLER_0_23_1138 ();
 sg13g2_decap_8 FILLER_0_23_1145 ();
 sg13g2_decap_8 FILLER_0_23_1152 ();
 sg13g2_decap_8 FILLER_0_23_1159 ();
 sg13g2_decap_8 FILLER_0_23_1166 ();
 sg13g2_decap_8 FILLER_0_23_1173 ();
 sg13g2_decap_8 FILLER_0_23_1180 ();
 sg13g2_decap_8 FILLER_0_23_1187 ();
 sg13g2_decap_8 FILLER_0_23_1194 ();
 sg13g2_decap_8 FILLER_0_23_1201 ();
 sg13g2_decap_8 FILLER_0_23_1208 ();
 sg13g2_decap_8 FILLER_0_23_1215 ();
 sg13g2_decap_4 FILLER_0_23_1222 ();
 sg13g2_fill_2 FILLER_0_23_1226 ();
 sg13g2_decap_8 FILLER_0_24_0 ();
 sg13g2_decap_8 FILLER_0_24_7 ();
 sg13g2_decap_4 FILLER_0_24_14 ();
 sg13g2_fill_1 FILLER_0_24_18 ();
 sg13g2_fill_2 FILLER_0_24_29 ();
 sg13g2_fill_1 FILLER_0_24_31 ();
 sg13g2_decap_4 FILLER_0_24_58 ();
 sg13g2_fill_1 FILLER_0_24_62 ();
 sg13g2_decap_8 FILLER_0_24_67 ();
 sg13g2_decap_8 FILLER_0_24_74 ();
 sg13g2_decap_8 FILLER_0_24_81 ();
 sg13g2_decap_4 FILLER_0_24_88 ();
 sg13g2_fill_2 FILLER_0_24_107 ();
 sg13g2_decap_8 FILLER_0_24_119 ();
 sg13g2_decap_8 FILLER_0_24_161 ();
 sg13g2_fill_2 FILLER_0_24_168 ();
 sg13g2_fill_1 FILLER_0_24_179 ();
 sg13g2_fill_1 FILLER_0_24_185 ();
 sg13g2_decap_4 FILLER_0_24_190 ();
 sg13g2_decap_8 FILLER_0_24_218 ();
 sg13g2_decap_8 FILLER_0_24_225 ();
 sg13g2_decap_8 FILLER_0_24_232 ();
 sg13g2_decap_8 FILLER_0_24_239 ();
 sg13g2_decap_8 FILLER_0_24_246 ();
 sg13g2_decap_8 FILLER_0_24_253 ();
 sg13g2_decap_8 FILLER_0_24_260 ();
 sg13g2_decap_8 FILLER_0_24_267 ();
 sg13g2_decap_4 FILLER_0_24_274 ();
 sg13g2_fill_1 FILLER_0_24_278 ();
 sg13g2_fill_1 FILLER_0_24_309 ();
 sg13g2_fill_2 FILLER_0_24_392 ();
 sg13g2_fill_2 FILLER_0_24_420 ();
 sg13g2_fill_1 FILLER_0_24_422 ();
 sg13g2_decap_8 FILLER_0_24_449 ();
 sg13g2_decap_8 FILLER_0_24_456 ();
 sg13g2_decap_4 FILLER_0_24_463 ();
 sg13g2_fill_1 FILLER_0_24_467 ();
 sg13g2_decap_4 FILLER_0_24_525 ();
 sg13g2_decap_4 FILLER_0_24_555 ();
 sg13g2_decap_8 FILLER_0_24_563 ();
 sg13g2_decap_8 FILLER_0_24_570 ();
 sg13g2_decap_8 FILLER_0_24_577 ();
 sg13g2_decap_8 FILLER_0_24_584 ();
 sg13g2_decap_8 FILLER_0_24_591 ();
 sg13g2_decap_8 FILLER_0_24_598 ();
 sg13g2_decap_8 FILLER_0_24_605 ();
 sg13g2_decap_8 FILLER_0_24_612 ();
 sg13g2_decap_8 FILLER_0_24_619 ();
 sg13g2_decap_8 FILLER_0_24_626 ();
 sg13g2_decap_8 FILLER_0_24_633 ();
 sg13g2_decap_8 FILLER_0_24_640 ();
 sg13g2_decap_8 FILLER_0_24_647 ();
 sg13g2_decap_8 FILLER_0_24_654 ();
 sg13g2_decap_8 FILLER_0_24_661 ();
 sg13g2_decap_8 FILLER_0_24_668 ();
 sg13g2_decap_8 FILLER_0_24_675 ();
 sg13g2_decap_8 FILLER_0_24_682 ();
 sg13g2_decap_8 FILLER_0_24_689 ();
 sg13g2_decap_8 FILLER_0_24_696 ();
 sg13g2_decap_8 FILLER_0_24_703 ();
 sg13g2_decap_8 FILLER_0_24_710 ();
 sg13g2_decap_8 FILLER_0_24_717 ();
 sg13g2_decap_8 FILLER_0_24_724 ();
 sg13g2_decap_8 FILLER_0_24_731 ();
 sg13g2_decap_8 FILLER_0_24_738 ();
 sg13g2_decap_8 FILLER_0_24_745 ();
 sg13g2_decap_8 FILLER_0_24_752 ();
 sg13g2_decap_8 FILLER_0_24_759 ();
 sg13g2_decap_8 FILLER_0_24_766 ();
 sg13g2_decap_8 FILLER_0_24_773 ();
 sg13g2_decap_8 FILLER_0_24_780 ();
 sg13g2_decap_8 FILLER_0_24_787 ();
 sg13g2_decap_8 FILLER_0_24_794 ();
 sg13g2_decap_8 FILLER_0_24_801 ();
 sg13g2_decap_8 FILLER_0_24_808 ();
 sg13g2_decap_8 FILLER_0_24_815 ();
 sg13g2_decap_8 FILLER_0_24_822 ();
 sg13g2_decap_8 FILLER_0_24_829 ();
 sg13g2_decap_8 FILLER_0_24_836 ();
 sg13g2_decap_8 FILLER_0_24_843 ();
 sg13g2_decap_8 FILLER_0_24_850 ();
 sg13g2_decap_8 FILLER_0_24_857 ();
 sg13g2_decap_8 FILLER_0_24_864 ();
 sg13g2_decap_8 FILLER_0_24_871 ();
 sg13g2_decap_8 FILLER_0_24_878 ();
 sg13g2_decap_8 FILLER_0_24_885 ();
 sg13g2_decap_8 FILLER_0_24_892 ();
 sg13g2_decap_8 FILLER_0_24_899 ();
 sg13g2_decap_8 FILLER_0_24_906 ();
 sg13g2_decap_8 FILLER_0_24_913 ();
 sg13g2_decap_8 FILLER_0_24_920 ();
 sg13g2_decap_8 FILLER_0_24_927 ();
 sg13g2_decap_8 FILLER_0_24_934 ();
 sg13g2_decap_8 FILLER_0_24_941 ();
 sg13g2_decap_8 FILLER_0_24_948 ();
 sg13g2_decap_8 FILLER_0_24_955 ();
 sg13g2_decap_8 FILLER_0_24_962 ();
 sg13g2_decap_4 FILLER_0_24_969 ();
 sg13g2_fill_1 FILLER_0_24_973 ();
 sg13g2_decap_4 FILLER_0_24_1052 ();
 sg13g2_fill_2 FILLER_0_24_1056 ();
 sg13g2_fill_2 FILLER_0_24_1063 ();
 sg13g2_decap_8 FILLER_0_24_1111 ();
 sg13g2_decap_8 FILLER_0_24_1118 ();
 sg13g2_decap_8 FILLER_0_24_1125 ();
 sg13g2_decap_8 FILLER_0_24_1132 ();
 sg13g2_decap_8 FILLER_0_24_1139 ();
 sg13g2_decap_8 FILLER_0_24_1146 ();
 sg13g2_decap_8 FILLER_0_24_1153 ();
 sg13g2_decap_8 FILLER_0_24_1160 ();
 sg13g2_decap_8 FILLER_0_24_1167 ();
 sg13g2_decap_8 FILLER_0_24_1174 ();
 sg13g2_decap_8 FILLER_0_24_1181 ();
 sg13g2_decap_8 FILLER_0_24_1188 ();
 sg13g2_decap_8 FILLER_0_24_1195 ();
 sg13g2_decap_8 FILLER_0_24_1202 ();
 sg13g2_decap_8 FILLER_0_24_1209 ();
 sg13g2_decap_8 FILLER_0_24_1216 ();
 sg13g2_decap_4 FILLER_0_24_1223 ();
 sg13g2_fill_1 FILLER_0_24_1227 ();
 sg13g2_decap_8 FILLER_0_25_0 ();
 sg13g2_fill_2 FILLER_0_25_77 ();
 sg13g2_fill_2 FILLER_0_25_161 ();
 sg13g2_decap_4 FILLER_0_25_199 ();
 sg13g2_fill_1 FILLER_0_25_244 ();
 sg13g2_decap_8 FILLER_0_25_249 ();
 sg13g2_decap_8 FILLER_0_25_256 ();
 sg13g2_decap_8 FILLER_0_25_263 ();
 sg13g2_decap_4 FILLER_0_25_270 ();
 sg13g2_fill_2 FILLER_0_25_274 ();
 sg13g2_decap_8 FILLER_0_25_291 ();
 sg13g2_fill_2 FILLER_0_25_349 ();
 sg13g2_fill_2 FILLER_0_25_377 ();
 sg13g2_fill_2 FILLER_0_25_415 ();
 sg13g2_decap_4 FILLER_0_25_427 ();
 sg13g2_decap_4 FILLER_0_25_435 ();
 sg13g2_decap_8 FILLER_0_25_449 ();
 sg13g2_fill_2 FILLER_0_25_456 ();
 sg13g2_fill_1 FILLER_0_25_484 ();
 sg13g2_fill_1 FILLER_0_25_490 ();
 sg13g2_fill_2 FILLER_0_25_501 ();
 sg13g2_decap_4 FILLER_0_25_528 ();
 sg13g2_decap_4 FILLER_0_25_536 ();
 sg13g2_decap_8 FILLER_0_25_617 ();
 sg13g2_decap_8 FILLER_0_25_624 ();
 sg13g2_decap_8 FILLER_0_25_631 ();
 sg13g2_decap_8 FILLER_0_25_638 ();
 sg13g2_decap_8 FILLER_0_25_645 ();
 sg13g2_decap_8 FILLER_0_25_652 ();
 sg13g2_decap_8 FILLER_0_25_659 ();
 sg13g2_decap_8 FILLER_0_25_666 ();
 sg13g2_decap_8 FILLER_0_25_673 ();
 sg13g2_decap_8 FILLER_0_25_680 ();
 sg13g2_decap_8 FILLER_0_25_687 ();
 sg13g2_decap_8 FILLER_0_25_694 ();
 sg13g2_decap_8 FILLER_0_25_701 ();
 sg13g2_decap_8 FILLER_0_25_708 ();
 sg13g2_decap_8 FILLER_0_25_715 ();
 sg13g2_decap_8 FILLER_0_25_722 ();
 sg13g2_decap_8 FILLER_0_25_729 ();
 sg13g2_decap_8 FILLER_0_25_736 ();
 sg13g2_decap_8 FILLER_0_25_743 ();
 sg13g2_decap_8 FILLER_0_25_750 ();
 sg13g2_decap_8 FILLER_0_25_757 ();
 sg13g2_decap_8 FILLER_0_25_764 ();
 sg13g2_decap_8 FILLER_0_25_771 ();
 sg13g2_decap_8 FILLER_0_25_778 ();
 sg13g2_decap_8 FILLER_0_25_785 ();
 sg13g2_decap_8 FILLER_0_25_792 ();
 sg13g2_decap_8 FILLER_0_25_799 ();
 sg13g2_decap_8 FILLER_0_25_806 ();
 sg13g2_decap_8 FILLER_0_25_813 ();
 sg13g2_decap_8 FILLER_0_25_820 ();
 sg13g2_decap_8 FILLER_0_25_827 ();
 sg13g2_decap_8 FILLER_0_25_834 ();
 sg13g2_decap_8 FILLER_0_25_841 ();
 sg13g2_decap_8 FILLER_0_25_848 ();
 sg13g2_decap_8 FILLER_0_25_855 ();
 sg13g2_decap_8 FILLER_0_25_862 ();
 sg13g2_decap_8 FILLER_0_25_869 ();
 sg13g2_decap_8 FILLER_0_25_876 ();
 sg13g2_decap_8 FILLER_0_25_883 ();
 sg13g2_decap_8 FILLER_0_25_890 ();
 sg13g2_decap_8 FILLER_0_25_897 ();
 sg13g2_decap_8 FILLER_0_25_904 ();
 sg13g2_decap_8 FILLER_0_25_911 ();
 sg13g2_decap_8 FILLER_0_25_918 ();
 sg13g2_decap_8 FILLER_0_25_925 ();
 sg13g2_decap_8 FILLER_0_25_932 ();
 sg13g2_decap_8 FILLER_0_25_939 ();
 sg13g2_decap_8 FILLER_0_25_946 ();
 sg13g2_decap_8 FILLER_0_25_953 ();
 sg13g2_decap_8 FILLER_0_25_960 ();
 sg13g2_decap_8 FILLER_0_25_967 ();
 sg13g2_decap_8 FILLER_0_25_974 ();
 sg13g2_decap_4 FILLER_0_25_981 ();
 sg13g2_fill_1 FILLER_0_25_1009 ();
 sg13g2_decap_4 FILLER_0_25_1014 ();
 sg13g2_decap_4 FILLER_0_25_1028 ();
 sg13g2_fill_1 FILLER_0_25_1032 ();
 sg13g2_decap_4 FILLER_0_25_1037 ();
 sg13g2_fill_2 FILLER_0_25_1041 ();
 sg13g2_fill_1 FILLER_0_25_1078 ();
 sg13g2_fill_1 FILLER_0_25_1088 ();
 sg13g2_decap_4 FILLER_0_25_1094 ();
 sg13g2_decap_8 FILLER_0_25_1138 ();
 sg13g2_decap_8 FILLER_0_25_1145 ();
 sg13g2_decap_8 FILLER_0_25_1152 ();
 sg13g2_decap_8 FILLER_0_25_1159 ();
 sg13g2_decap_8 FILLER_0_25_1166 ();
 sg13g2_decap_8 FILLER_0_25_1173 ();
 sg13g2_decap_8 FILLER_0_25_1180 ();
 sg13g2_decap_8 FILLER_0_25_1187 ();
 sg13g2_decap_8 FILLER_0_25_1194 ();
 sg13g2_decap_8 FILLER_0_25_1201 ();
 sg13g2_decap_8 FILLER_0_25_1208 ();
 sg13g2_decap_8 FILLER_0_25_1215 ();
 sg13g2_decap_4 FILLER_0_25_1222 ();
 sg13g2_fill_2 FILLER_0_25_1226 ();
 sg13g2_fill_1 FILLER_0_26_0 ();
 sg13g2_fill_2 FILLER_0_26_45 ();
 sg13g2_fill_1 FILLER_0_26_51 ();
 sg13g2_fill_1 FILLER_0_26_78 ();
 sg13g2_fill_1 FILLER_0_26_105 ();
 sg13g2_fill_1 FILLER_0_26_126 ();
 sg13g2_fill_1 FILLER_0_26_137 ();
 sg13g2_fill_1 FILLER_0_26_148 ();
 sg13g2_fill_2 FILLER_0_26_175 ();
 sg13g2_fill_1 FILLER_0_26_229 ();
 sg13g2_decap_8 FILLER_0_26_256 ();
 sg13g2_decap_8 FILLER_0_26_309 ();
 sg13g2_fill_1 FILLER_0_26_316 ();
 sg13g2_fill_2 FILLER_0_26_397 ();
 sg13g2_decap_8 FILLER_0_26_445 ();
 sg13g2_decap_8 FILLER_0_26_452 ();
 sg13g2_decap_4 FILLER_0_26_459 ();
 sg13g2_fill_2 FILLER_0_26_463 ();
 sg13g2_fill_2 FILLER_0_26_469 ();
 sg13g2_fill_2 FILLER_0_26_476 ();
 sg13g2_fill_1 FILLER_0_26_478 ();
 sg13g2_decap_8 FILLER_0_26_489 ();
 sg13g2_decap_8 FILLER_0_26_496 ();
 sg13g2_fill_2 FILLER_0_26_503 ();
 sg13g2_fill_1 FILLER_0_26_505 ();
 sg13g2_decap_8 FILLER_0_26_518 ();
 sg13g2_fill_2 FILLER_0_26_525 ();
 sg13g2_decap_8 FILLER_0_26_531 ();
 sg13g2_fill_2 FILLER_0_26_563 ();
 sg13g2_fill_1 FILLER_0_26_565 ();
 sg13g2_decap_8 FILLER_0_26_601 ();
 sg13g2_decap_8 FILLER_0_26_608 ();
 sg13g2_decap_8 FILLER_0_26_615 ();
 sg13g2_decap_8 FILLER_0_26_622 ();
 sg13g2_decap_8 FILLER_0_26_629 ();
 sg13g2_decap_8 FILLER_0_26_636 ();
 sg13g2_decap_8 FILLER_0_26_643 ();
 sg13g2_decap_8 FILLER_0_26_650 ();
 sg13g2_decap_8 FILLER_0_26_657 ();
 sg13g2_decap_8 FILLER_0_26_664 ();
 sg13g2_decap_8 FILLER_0_26_671 ();
 sg13g2_decap_8 FILLER_0_26_678 ();
 sg13g2_decap_8 FILLER_0_26_685 ();
 sg13g2_decap_8 FILLER_0_26_692 ();
 sg13g2_decap_8 FILLER_0_26_699 ();
 sg13g2_decap_8 FILLER_0_26_706 ();
 sg13g2_decap_8 FILLER_0_26_713 ();
 sg13g2_decap_8 FILLER_0_26_720 ();
 sg13g2_decap_8 FILLER_0_26_727 ();
 sg13g2_decap_8 FILLER_0_26_734 ();
 sg13g2_decap_8 FILLER_0_26_741 ();
 sg13g2_decap_8 FILLER_0_26_748 ();
 sg13g2_decap_8 FILLER_0_26_755 ();
 sg13g2_decap_8 FILLER_0_26_762 ();
 sg13g2_decap_8 FILLER_0_26_769 ();
 sg13g2_decap_4 FILLER_0_26_776 ();
 sg13g2_decap_8 FILLER_0_26_811 ();
 sg13g2_decap_8 FILLER_0_26_818 ();
 sg13g2_decap_8 FILLER_0_26_825 ();
 sg13g2_decap_8 FILLER_0_26_832 ();
 sg13g2_decap_8 FILLER_0_26_839 ();
 sg13g2_decap_8 FILLER_0_26_846 ();
 sg13g2_decap_8 FILLER_0_26_853 ();
 sg13g2_decap_8 FILLER_0_26_860 ();
 sg13g2_decap_8 FILLER_0_26_867 ();
 sg13g2_decap_8 FILLER_0_26_874 ();
 sg13g2_decap_8 FILLER_0_26_881 ();
 sg13g2_decap_8 FILLER_0_26_888 ();
 sg13g2_decap_8 FILLER_0_26_895 ();
 sg13g2_decap_8 FILLER_0_26_902 ();
 sg13g2_decap_8 FILLER_0_26_909 ();
 sg13g2_decap_8 FILLER_0_26_916 ();
 sg13g2_decap_8 FILLER_0_26_923 ();
 sg13g2_decap_8 FILLER_0_26_930 ();
 sg13g2_decap_8 FILLER_0_26_937 ();
 sg13g2_decap_8 FILLER_0_26_944 ();
 sg13g2_decap_8 FILLER_0_26_951 ();
 sg13g2_decap_8 FILLER_0_26_958 ();
 sg13g2_decap_8 FILLER_0_26_965 ();
 sg13g2_fill_2 FILLER_0_26_972 ();
 sg13g2_fill_2 FILLER_0_26_979 ();
 sg13g2_fill_1 FILLER_0_26_985 ();
 sg13g2_fill_2 FILLER_0_26_996 ();
 sg13g2_decap_8 FILLER_0_26_1008 ();
 sg13g2_fill_2 FILLER_0_26_1027 ();
 sg13g2_decap_8 FILLER_0_26_1039 ();
 sg13g2_decap_4 FILLER_0_26_1046 ();
 sg13g2_fill_1 FILLER_0_26_1050 ();
 sg13g2_fill_2 FILLER_0_26_1055 ();
 sg13g2_fill_2 FILLER_0_26_1062 ();
 sg13g2_fill_1 FILLER_0_26_1064 ();
 sg13g2_decap_4 FILLER_0_26_1096 ();
 sg13g2_fill_2 FILLER_0_26_1100 ();
 sg13g2_fill_2 FILLER_0_26_1117 ();
 sg13g2_decap_8 FILLER_0_26_1123 ();
 sg13g2_decap_8 FILLER_0_26_1130 ();
 sg13g2_decap_8 FILLER_0_26_1137 ();
 sg13g2_decap_8 FILLER_0_26_1144 ();
 sg13g2_decap_8 FILLER_0_26_1151 ();
 sg13g2_decap_8 FILLER_0_26_1158 ();
 sg13g2_decap_8 FILLER_0_26_1165 ();
 sg13g2_decap_8 FILLER_0_26_1172 ();
 sg13g2_decap_8 FILLER_0_26_1179 ();
 sg13g2_decap_8 FILLER_0_26_1186 ();
 sg13g2_decap_8 FILLER_0_26_1193 ();
 sg13g2_decap_8 FILLER_0_26_1200 ();
 sg13g2_decap_8 FILLER_0_26_1207 ();
 sg13g2_decap_8 FILLER_0_26_1214 ();
 sg13g2_decap_8 FILLER_0_26_1221 ();
 sg13g2_decap_4 FILLER_0_27_0 ();
 sg13g2_fill_1 FILLER_0_27_4 ();
 sg13g2_fill_1 FILLER_0_27_34 ();
 sg13g2_fill_2 FILLER_0_27_40 ();
 sg13g2_fill_1 FILLER_0_27_47 ();
 sg13g2_fill_2 FILLER_0_27_63 ();
 sg13g2_fill_1 FILLER_0_27_65 ();
 sg13g2_decap_8 FILLER_0_27_76 ();
 sg13g2_decap_4 FILLER_0_27_83 ();
 sg13g2_decap_8 FILLER_0_27_91 ();
 sg13g2_decap_4 FILLER_0_27_98 ();
 sg13g2_fill_1 FILLER_0_27_102 ();
 sg13g2_decap_8 FILLER_0_27_118 ();
 sg13g2_fill_2 FILLER_0_27_125 ();
 sg13g2_fill_1 FILLER_0_27_127 ();
 sg13g2_decap_8 FILLER_0_27_133 ();
 sg13g2_fill_1 FILLER_0_27_140 ();
 sg13g2_fill_2 FILLER_0_27_164 ();
 sg13g2_fill_1 FILLER_0_27_166 ();
 sg13g2_fill_2 FILLER_0_27_177 ();
 sg13g2_fill_1 FILLER_0_27_189 ();
 sg13g2_decap_4 FILLER_0_27_229 ();
 sg13g2_fill_2 FILLER_0_27_233 ();
 sg13g2_decap_8 FILLER_0_27_265 ();
 sg13g2_fill_2 FILLER_0_27_272 ();
 sg13g2_fill_1 FILLER_0_27_281 ();
 sg13g2_decap_8 FILLER_0_27_308 ();
 sg13g2_decap_8 FILLER_0_27_315 ();
 sg13g2_decap_8 FILLER_0_27_322 ();
 sg13g2_decap_8 FILLER_0_27_329 ();
 sg13g2_decap_4 FILLER_0_27_336 ();
 sg13g2_decap_8 FILLER_0_27_351 ();
 sg13g2_decap_8 FILLER_0_27_358 ();
 sg13g2_decap_8 FILLER_0_27_365 ();
 sg13g2_decap_8 FILLER_0_27_372 ();
 sg13g2_decap_8 FILLER_0_27_379 ();
 sg13g2_decap_4 FILLER_0_27_386 ();
 sg13g2_fill_2 FILLER_0_27_390 ();
 sg13g2_decap_4 FILLER_0_27_397 ();
 sg13g2_fill_2 FILLER_0_27_401 ();
 sg13g2_decap_8 FILLER_0_27_423 ();
 sg13g2_decap_8 FILLER_0_27_430 ();
 sg13g2_decap_8 FILLER_0_27_441 ();
 sg13g2_decap_8 FILLER_0_27_448 ();
 sg13g2_decap_8 FILLER_0_27_455 ();
 sg13g2_decap_8 FILLER_0_27_462 ();
 sg13g2_decap_4 FILLER_0_27_469 ();
 sg13g2_fill_2 FILLER_0_27_473 ();
 sg13g2_fill_2 FILLER_0_27_480 ();
 sg13g2_decap_8 FILLER_0_27_508 ();
 sg13g2_fill_2 FILLER_0_27_515 ();
 sg13g2_fill_1 FILLER_0_27_517 ();
 sg13g2_decap_8 FILLER_0_27_523 ();
 sg13g2_fill_2 FILLER_0_27_530 ();
 sg13g2_fill_1 FILLER_0_27_532 ();
 sg13g2_fill_1 FILLER_0_27_569 ();
 sg13g2_fill_2 FILLER_0_27_580 ();
 sg13g2_decap_8 FILLER_0_27_586 ();
 sg13g2_decap_8 FILLER_0_27_593 ();
 sg13g2_decap_8 FILLER_0_27_600 ();
 sg13g2_decap_8 FILLER_0_27_607 ();
 sg13g2_decap_8 FILLER_0_27_614 ();
 sg13g2_decap_8 FILLER_0_27_621 ();
 sg13g2_decap_8 FILLER_0_27_628 ();
 sg13g2_decap_8 FILLER_0_27_635 ();
 sg13g2_decap_8 FILLER_0_27_642 ();
 sg13g2_decap_8 FILLER_0_27_649 ();
 sg13g2_decap_8 FILLER_0_27_656 ();
 sg13g2_decap_8 FILLER_0_27_663 ();
 sg13g2_decap_8 FILLER_0_27_670 ();
 sg13g2_decap_8 FILLER_0_27_677 ();
 sg13g2_decap_8 FILLER_0_27_684 ();
 sg13g2_decap_8 FILLER_0_27_691 ();
 sg13g2_decap_8 FILLER_0_27_698 ();
 sg13g2_decap_8 FILLER_0_27_705 ();
 sg13g2_decap_8 FILLER_0_27_712 ();
 sg13g2_decap_8 FILLER_0_27_719 ();
 sg13g2_decap_8 FILLER_0_27_726 ();
 sg13g2_decap_8 FILLER_0_27_733 ();
 sg13g2_decap_8 FILLER_0_27_740 ();
 sg13g2_decap_4 FILLER_0_27_747 ();
 sg13g2_fill_2 FILLER_0_27_782 ();
 sg13g2_decap_8 FILLER_0_27_828 ();
 sg13g2_decap_8 FILLER_0_27_835 ();
 sg13g2_decap_8 FILLER_0_27_842 ();
 sg13g2_decap_8 FILLER_0_27_849 ();
 sg13g2_decap_8 FILLER_0_27_856 ();
 sg13g2_decap_8 FILLER_0_27_863 ();
 sg13g2_decap_8 FILLER_0_27_870 ();
 sg13g2_decap_8 FILLER_0_27_877 ();
 sg13g2_decap_8 FILLER_0_27_884 ();
 sg13g2_decap_8 FILLER_0_27_891 ();
 sg13g2_decap_8 FILLER_0_27_898 ();
 sg13g2_decap_8 FILLER_0_27_905 ();
 sg13g2_decap_8 FILLER_0_27_912 ();
 sg13g2_decap_8 FILLER_0_27_919 ();
 sg13g2_decap_8 FILLER_0_27_926 ();
 sg13g2_decap_8 FILLER_0_27_933 ();
 sg13g2_decap_8 FILLER_0_27_940 ();
 sg13g2_decap_8 FILLER_0_27_947 ();
 sg13g2_decap_8 FILLER_0_27_954 ();
 sg13g2_decap_8 FILLER_0_27_961 ();
 sg13g2_decap_8 FILLER_0_27_968 ();
 sg13g2_fill_2 FILLER_0_27_975 ();
 sg13g2_fill_1 FILLER_0_27_977 ();
 sg13g2_decap_8 FILLER_0_27_1004 ();
 sg13g2_decap_8 FILLER_0_27_1037 ();
 sg13g2_decap_8 FILLER_0_27_1044 ();
 sg13g2_fill_2 FILLER_0_27_1051 ();
 sg13g2_decap_8 FILLER_0_27_1083 ();
 sg13g2_decap_8 FILLER_0_27_1090 ();
 sg13g2_decap_4 FILLER_0_27_1097 ();
 sg13g2_decap_8 FILLER_0_27_1132 ();
 sg13g2_decap_8 FILLER_0_27_1139 ();
 sg13g2_decap_8 FILLER_0_27_1146 ();
 sg13g2_decap_8 FILLER_0_27_1153 ();
 sg13g2_decap_8 FILLER_0_27_1160 ();
 sg13g2_decap_8 FILLER_0_27_1167 ();
 sg13g2_decap_8 FILLER_0_27_1174 ();
 sg13g2_decap_8 FILLER_0_27_1181 ();
 sg13g2_decap_8 FILLER_0_27_1188 ();
 sg13g2_decap_8 FILLER_0_27_1195 ();
 sg13g2_decap_8 FILLER_0_27_1202 ();
 sg13g2_decap_8 FILLER_0_27_1209 ();
 sg13g2_decap_8 FILLER_0_27_1216 ();
 sg13g2_decap_4 FILLER_0_27_1223 ();
 sg13g2_fill_1 FILLER_0_27_1227 ();
 sg13g2_fill_1 FILLER_0_28_4 ();
 sg13g2_fill_2 FILLER_0_28_36 ();
 sg13g2_fill_1 FILLER_0_28_38 ();
 sg13g2_decap_8 FILLER_0_28_65 ();
 sg13g2_decap_8 FILLER_0_28_72 ();
 sg13g2_decap_4 FILLER_0_28_79 ();
 sg13g2_fill_1 FILLER_0_28_87 ();
 sg13g2_fill_2 FILLER_0_28_114 ();
 sg13g2_decap_8 FILLER_0_28_147 ();
 sg13g2_decap_8 FILLER_0_28_154 ();
 sg13g2_decap_8 FILLER_0_28_161 ();
 sg13g2_decap_8 FILLER_0_28_168 ();
 sg13g2_decap_4 FILLER_0_28_175 ();
 sg13g2_fill_2 FILLER_0_28_179 ();
 sg13g2_decap_8 FILLER_0_28_184 ();
 sg13g2_decap_4 FILLER_0_28_191 ();
 sg13g2_decap_4 FILLER_0_28_204 ();
 sg13g2_decap_8 FILLER_0_28_220 ();
 sg13g2_decap_8 FILLER_0_28_256 ();
 sg13g2_fill_2 FILLER_0_28_263 ();
 sg13g2_fill_1 FILLER_0_28_265 ();
 sg13g2_decap_8 FILLER_0_28_289 ();
 sg13g2_fill_2 FILLER_0_28_296 ();
 sg13g2_fill_1 FILLER_0_28_298 ();
 sg13g2_decap_8 FILLER_0_28_303 ();
 sg13g2_decap_8 FILLER_0_28_310 ();
 sg13g2_decap_8 FILLER_0_28_317 ();
 sg13g2_fill_1 FILLER_0_28_344 ();
 sg13g2_decap_8 FILLER_0_28_359 ();
 sg13g2_decap_8 FILLER_0_28_366 ();
 sg13g2_decap_8 FILLER_0_28_373 ();
 sg13g2_decap_4 FILLER_0_28_385 ();
 sg13g2_fill_1 FILLER_0_28_389 ();
 sg13g2_fill_1 FILLER_0_28_416 ();
 sg13g2_decap_8 FILLER_0_28_443 ();
 sg13g2_decap_8 FILLER_0_28_450 ();
 sg13g2_decap_8 FILLER_0_28_457 ();
 sg13g2_fill_1 FILLER_0_28_464 ();
 sg13g2_fill_2 FILLER_0_28_476 ();
 sg13g2_fill_1 FILLER_0_28_478 ();
 sg13g2_decap_8 FILLER_0_28_493 ();
 sg13g2_decap_8 FILLER_0_28_500 ();
 sg13g2_decap_8 FILLER_0_28_507 ();
 sg13g2_fill_1 FILLER_0_28_549 ();
 sg13g2_decap_8 FILLER_0_28_562 ();
 sg13g2_decap_8 FILLER_0_28_569 ();
 sg13g2_decap_8 FILLER_0_28_576 ();
 sg13g2_decap_8 FILLER_0_28_583 ();
 sg13g2_decap_4 FILLER_0_28_590 ();
 sg13g2_fill_2 FILLER_0_28_594 ();
 sg13g2_decap_8 FILLER_0_28_601 ();
 sg13g2_decap_8 FILLER_0_28_608 ();
 sg13g2_decap_8 FILLER_0_28_615 ();
 sg13g2_decap_8 FILLER_0_28_622 ();
 sg13g2_decap_8 FILLER_0_28_629 ();
 sg13g2_decap_8 FILLER_0_28_636 ();
 sg13g2_decap_8 FILLER_0_28_643 ();
 sg13g2_decap_8 FILLER_0_28_650 ();
 sg13g2_decap_8 FILLER_0_28_657 ();
 sg13g2_decap_8 FILLER_0_28_664 ();
 sg13g2_decap_8 FILLER_0_28_671 ();
 sg13g2_decap_8 FILLER_0_28_678 ();
 sg13g2_decap_8 FILLER_0_28_685 ();
 sg13g2_decap_8 FILLER_0_28_692 ();
 sg13g2_decap_8 FILLER_0_28_699 ();
 sg13g2_decap_8 FILLER_0_28_706 ();
 sg13g2_decap_8 FILLER_0_28_713 ();
 sg13g2_decap_8 FILLER_0_28_720 ();
 sg13g2_decap_8 FILLER_0_28_727 ();
 sg13g2_decap_8 FILLER_0_28_734 ();
 sg13g2_decap_4 FILLER_0_28_741 ();
 sg13g2_fill_1 FILLER_0_28_745 ();
 sg13g2_fill_2 FILLER_0_28_751 ();
 sg13g2_fill_1 FILLER_0_28_767 ();
 sg13g2_fill_2 FILLER_0_28_812 ();
 sg13g2_fill_1 FILLER_0_28_814 ();
 sg13g2_decap_8 FILLER_0_28_841 ();
 sg13g2_decap_8 FILLER_0_28_848 ();
 sg13g2_decap_8 FILLER_0_28_855 ();
 sg13g2_decap_8 FILLER_0_28_862 ();
 sg13g2_decap_8 FILLER_0_28_869 ();
 sg13g2_decap_8 FILLER_0_28_876 ();
 sg13g2_decap_8 FILLER_0_28_883 ();
 sg13g2_decap_8 FILLER_0_28_890 ();
 sg13g2_decap_8 FILLER_0_28_897 ();
 sg13g2_decap_8 FILLER_0_28_904 ();
 sg13g2_decap_8 FILLER_0_28_911 ();
 sg13g2_decap_8 FILLER_0_28_918 ();
 sg13g2_decap_8 FILLER_0_28_925 ();
 sg13g2_decap_8 FILLER_0_28_932 ();
 sg13g2_decap_8 FILLER_0_28_939 ();
 sg13g2_decap_8 FILLER_0_28_946 ();
 sg13g2_decap_8 FILLER_0_28_953 ();
 sg13g2_decap_8 FILLER_0_28_960 ();
 sg13g2_decap_8 FILLER_0_28_967 ();
 sg13g2_decap_4 FILLER_0_28_1005 ();
 sg13g2_fill_1 FILLER_0_28_1009 ();
 sg13g2_decap_8 FILLER_0_28_1052 ();
 sg13g2_fill_1 FILLER_0_28_1059 ();
 sg13g2_fill_1 FILLER_0_28_1065 ();
 sg13g2_decap_8 FILLER_0_28_1121 ();
 sg13g2_decap_8 FILLER_0_28_1128 ();
 sg13g2_decap_8 FILLER_0_28_1135 ();
 sg13g2_decap_8 FILLER_0_28_1142 ();
 sg13g2_decap_8 FILLER_0_28_1149 ();
 sg13g2_decap_8 FILLER_0_28_1156 ();
 sg13g2_decap_8 FILLER_0_28_1163 ();
 sg13g2_decap_8 FILLER_0_28_1170 ();
 sg13g2_decap_8 FILLER_0_28_1177 ();
 sg13g2_decap_8 FILLER_0_28_1184 ();
 sg13g2_decap_8 FILLER_0_28_1191 ();
 sg13g2_decap_8 FILLER_0_28_1198 ();
 sg13g2_decap_8 FILLER_0_28_1205 ();
 sg13g2_decap_8 FILLER_0_28_1212 ();
 sg13g2_decap_8 FILLER_0_28_1219 ();
 sg13g2_fill_2 FILLER_0_28_1226 ();
 sg13g2_decap_8 FILLER_0_29_0 ();
 sg13g2_fill_2 FILLER_0_29_7 ();
 sg13g2_fill_1 FILLER_0_29_9 ();
 sg13g2_decap_8 FILLER_0_29_14 ();
 sg13g2_decap_4 FILLER_0_29_21 ();
 sg13g2_fill_2 FILLER_0_29_35 ();
 sg13g2_fill_1 FILLER_0_29_37 ();
 sg13g2_fill_2 FILLER_0_29_42 ();
 sg13g2_fill_1 FILLER_0_29_44 ();
 sg13g2_decap_8 FILLER_0_29_69 ();
 sg13g2_decap_8 FILLER_0_29_76 ();
 sg13g2_fill_1 FILLER_0_29_103 ();
 sg13g2_fill_2 FILLER_0_29_114 ();
 sg13g2_fill_2 FILLER_0_29_126 ();
 sg13g2_fill_2 FILLER_0_29_133 ();
 sg13g2_fill_1 FILLER_0_29_135 ();
 sg13g2_decap_8 FILLER_0_29_201 ();
 sg13g2_decap_4 FILLER_0_29_208 ();
 sg13g2_decap_4 FILLER_0_29_222 ();
 sg13g2_fill_1 FILLER_0_29_226 ();
 sg13g2_fill_1 FILLER_0_29_267 ();
 sg13g2_decap_8 FILLER_0_29_298 ();
 sg13g2_decap_8 FILLER_0_29_305 ();
 sg13g2_fill_1 FILLER_0_29_312 ();
 sg13g2_fill_2 FILLER_0_29_365 ();
 sg13g2_decap_4 FILLER_0_29_422 ();
 sg13g2_decap_8 FILLER_0_29_430 ();
 sg13g2_decap_8 FILLER_0_29_437 ();
 sg13g2_decap_8 FILLER_0_29_444 ();
 sg13g2_decap_8 FILLER_0_29_451 ();
 sg13g2_decap_8 FILLER_0_29_458 ();
 sg13g2_decap_8 FILLER_0_29_465 ();
 sg13g2_fill_2 FILLER_0_29_513 ();
 sg13g2_fill_2 FILLER_0_29_545 ();
 sg13g2_fill_1 FILLER_0_29_555 ();
 sg13g2_decap_8 FILLER_0_29_560 ();
 sg13g2_fill_1 FILLER_0_29_567 ();
 sg13g2_decap_8 FILLER_0_29_625 ();
 sg13g2_decap_8 FILLER_0_29_632 ();
 sg13g2_decap_8 FILLER_0_29_639 ();
 sg13g2_decap_8 FILLER_0_29_646 ();
 sg13g2_decap_8 FILLER_0_29_653 ();
 sg13g2_decap_8 FILLER_0_29_660 ();
 sg13g2_decap_8 FILLER_0_29_667 ();
 sg13g2_decap_8 FILLER_0_29_674 ();
 sg13g2_decap_8 FILLER_0_29_681 ();
 sg13g2_decap_8 FILLER_0_29_688 ();
 sg13g2_decap_8 FILLER_0_29_695 ();
 sg13g2_decap_8 FILLER_0_29_702 ();
 sg13g2_decap_8 FILLER_0_29_709 ();
 sg13g2_decap_8 FILLER_0_29_716 ();
 sg13g2_decap_8 FILLER_0_29_723 ();
 sg13g2_decap_8 FILLER_0_29_730 ();
 sg13g2_decap_4 FILLER_0_29_737 ();
 sg13g2_fill_2 FILLER_0_29_741 ();
 sg13g2_decap_8 FILLER_0_29_748 ();
 sg13g2_fill_2 FILLER_0_29_755 ();
 sg13g2_decap_8 FILLER_0_29_767 ();
 sg13g2_decap_8 FILLER_0_29_778 ();
 sg13g2_decap_4 FILLER_0_29_785 ();
 sg13g2_fill_2 FILLER_0_29_794 ();
 sg13g2_decap_8 FILLER_0_29_829 ();
 sg13g2_decap_8 FILLER_0_29_836 ();
 sg13g2_decap_8 FILLER_0_29_843 ();
 sg13g2_decap_8 FILLER_0_29_850 ();
 sg13g2_decap_8 FILLER_0_29_857 ();
 sg13g2_decap_8 FILLER_0_29_864 ();
 sg13g2_decap_8 FILLER_0_29_871 ();
 sg13g2_decap_8 FILLER_0_29_878 ();
 sg13g2_decap_8 FILLER_0_29_885 ();
 sg13g2_decap_8 FILLER_0_29_892 ();
 sg13g2_decap_8 FILLER_0_29_899 ();
 sg13g2_decap_8 FILLER_0_29_906 ();
 sg13g2_decap_8 FILLER_0_29_913 ();
 sg13g2_decap_8 FILLER_0_29_920 ();
 sg13g2_decap_8 FILLER_0_29_927 ();
 sg13g2_decap_8 FILLER_0_29_934 ();
 sg13g2_decap_8 FILLER_0_29_941 ();
 sg13g2_decap_8 FILLER_0_29_948 ();
 sg13g2_decap_8 FILLER_0_29_955 ();
 sg13g2_decap_8 FILLER_0_29_962 ();
 sg13g2_fill_2 FILLER_0_29_969 ();
 sg13g2_fill_1 FILLER_0_29_971 ();
 sg13g2_decap_4 FILLER_0_29_982 ();
 sg13g2_decap_8 FILLER_0_29_990 ();
 sg13g2_fill_1 FILLER_0_29_1059 ();
 sg13g2_decap_8 FILLER_0_29_1079 ();
 sg13g2_decap_8 FILLER_0_29_1116 ();
 sg13g2_decap_8 FILLER_0_29_1123 ();
 sg13g2_decap_8 FILLER_0_29_1130 ();
 sg13g2_decap_8 FILLER_0_29_1137 ();
 sg13g2_decap_8 FILLER_0_29_1144 ();
 sg13g2_decap_8 FILLER_0_29_1151 ();
 sg13g2_decap_8 FILLER_0_29_1158 ();
 sg13g2_decap_8 FILLER_0_29_1165 ();
 sg13g2_decap_8 FILLER_0_29_1172 ();
 sg13g2_decap_8 FILLER_0_29_1179 ();
 sg13g2_decap_8 FILLER_0_29_1186 ();
 sg13g2_decap_8 FILLER_0_29_1193 ();
 sg13g2_decap_8 FILLER_0_29_1200 ();
 sg13g2_decap_8 FILLER_0_29_1207 ();
 sg13g2_decap_8 FILLER_0_29_1214 ();
 sg13g2_decap_8 FILLER_0_29_1221 ();
 sg13g2_fill_2 FILLER_0_30_0 ();
 sg13g2_fill_1 FILLER_0_30_2 ();
 sg13g2_fill_2 FILLER_0_30_34 ();
 sg13g2_fill_1 FILLER_0_30_41 ();
 sg13g2_fill_2 FILLER_0_30_126 ();
 sg13g2_fill_2 FILLER_0_30_148 ();
 sg13g2_fill_1 FILLER_0_30_198 ();
 sg13g2_fill_1 FILLER_0_30_225 ();
 sg13g2_fill_1 FILLER_0_30_262 ();
 sg13g2_fill_2 FILLER_0_30_273 ();
 sg13g2_fill_1 FILLER_0_30_275 ();
 sg13g2_decap_8 FILLER_0_30_291 ();
 sg13g2_fill_2 FILLER_0_30_298 ();
 sg13g2_fill_1 FILLER_0_30_335 ();
 sg13g2_decap_4 FILLER_0_30_341 ();
 sg13g2_fill_2 FILLER_0_30_376 ();
 sg13g2_fill_1 FILLER_0_30_387 ();
 sg13g2_fill_2 FILLER_0_30_396 ();
 sg13g2_decap_8 FILLER_0_30_417 ();
 sg13g2_decap_8 FILLER_0_30_424 ();
 sg13g2_decap_8 FILLER_0_30_431 ();
 sg13g2_decap_8 FILLER_0_30_438 ();
 sg13g2_decap_8 FILLER_0_30_445 ();
 sg13g2_decap_8 FILLER_0_30_452 ();
 sg13g2_decap_8 FILLER_0_30_459 ();
 sg13g2_decap_4 FILLER_0_30_466 ();
 sg13g2_decap_8 FILLER_0_30_505 ();
 sg13g2_decap_8 FILLER_0_30_512 ();
 sg13g2_fill_1 FILLER_0_30_575 ();
 sg13g2_fill_1 FILLER_0_30_586 ();
 sg13g2_decap_8 FILLER_0_30_597 ();
 sg13g2_fill_1 FILLER_0_30_604 ();
 sg13g2_decap_8 FILLER_0_30_609 ();
 sg13g2_decap_4 FILLER_0_30_616 ();
 sg13g2_fill_2 FILLER_0_30_620 ();
 sg13g2_decap_8 FILLER_0_30_634 ();
 sg13g2_decap_8 FILLER_0_30_641 ();
 sg13g2_decap_8 FILLER_0_30_648 ();
 sg13g2_decap_8 FILLER_0_30_655 ();
 sg13g2_decap_8 FILLER_0_30_662 ();
 sg13g2_decap_8 FILLER_0_30_669 ();
 sg13g2_decap_8 FILLER_0_30_676 ();
 sg13g2_decap_8 FILLER_0_30_683 ();
 sg13g2_decap_8 FILLER_0_30_690 ();
 sg13g2_decap_8 FILLER_0_30_697 ();
 sg13g2_decap_8 FILLER_0_30_704 ();
 sg13g2_decap_8 FILLER_0_30_711 ();
 sg13g2_decap_8 FILLER_0_30_718 ();
 sg13g2_decap_8 FILLER_0_30_725 ();
 sg13g2_decap_8 FILLER_0_30_732 ();
 sg13g2_decap_4 FILLER_0_30_739 ();
 sg13g2_decap_8 FILLER_0_30_769 ();
 sg13g2_decap_8 FILLER_0_30_776 ();
 sg13g2_decap_8 FILLER_0_30_783 ();
 sg13g2_decap_8 FILLER_0_30_790 ();
 sg13g2_decap_8 FILLER_0_30_797 ();
 sg13g2_fill_2 FILLER_0_30_804 ();
 sg13g2_fill_1 FILLER_0_30_806 ();
 sg13g2_decap_8 FILLER_0_30_822 ();
 sg13g2_decap_8 FILLER_0_30_829 ();
 sg13g2_decap_8 FILLER_0_30_836 ();
 sg13g2_decap_8 FILLER_0_30_843 ();
 sg13g2_decap_8 FILLER_0_30_850 ();
 sg13g2_decap_8 FILLER_0_30_857 ();
 sg13g2_decap_8 FILLER_0_30_864 ();
 sg13g2_decap_8 FILLER_0_30_871 ();
 sg13g2_decap_8 FILLER_0_30_878 ();
 sg13g2_decap_8 FILLER_0_30_885 ();
 sg13g2_decap_8 FILLER_0_30_892 ();
 sg13g2_decap_8 FILLER_0_30_899 ();
 sg13g2_decap_8 FILLER_0_30_906 ();
 sg13g2_decap_8 FILLER_0_30_913 ();
 sg13g2_decap_8 FILLER_0_30_920 ();
 sg13g2_decap_8 FILLER_0_30_927 ();
 sg13g2_decap_8 FILLER_0_30_934 ();
 sg13g2_decap_8 FILLER_0_30_941 ();
 sg13g2_decap_8 FILLER_0_30_948 ();
 sg13g2_decap_4 FILLER_0_30_955 ();
 sg13g2_decap_4 FILLER_0_30_1000 ();
 sg13g2_fill_1 FILLER_0_30_1004 ();
 sg13g2_decap_8 FILLER_0_30_1009 ();
 sg13g2_decap_4 FILLER_0_30_1016 ();
 sg13g2_fill_1 FILLER_0_30_1064 ();
 sg13g2_decap_4 FILLER_0_30_1077 ();
 sg13g2_fill_1 FILLER_0_30_1081 ();
 sg13g2_decap_8 FILLER_0_30_1108 ();
 sg13g2_decap_8 FILLER_0_30_1115 ();
 sg13g2_decap_8 FILLER_0_30_1122 ();
 sg13g2_decap_8 FILLER_0_30_1129 ();
 sg13g2_decap_8 FILLER_0_30_1136 ();
 sg13g2_decap_8 FILLER_0_30_1143 ();
 sg13g2_decap_8 FILLER_0_30_1150 ();
 sg13g2_decap_8 FILLER_0_30_1157 ();
 sg13g2_decap_8 FILLER_0_30_1164 ();
 sg13g2_decap_8 FILLER_0_30_1171 ();
 sg13g2_decap_8 FILLER_0_30_1178 ();
 sg13g2_decap_8 FILLER_0_30_1185 ();
 sg13g2_decap_8 FILLER_0_30_1192 ();
 sg13g2_decap_8 FILLER_0_30_1199 ();
 sg13g2_decap_8 FILLER_0_30_1206 ();
 sg13g2_decap_8 FILLER_0_30_1213 ();
 sg13g2_decap_8 FILLER_0_30_1220 ();
 sg13g2_fill_1 FILLER_0_30_1227 ();
 sg13g2_decap_4 FILLER_0_31_0 ();
 sg13g2_fill_1 FILLER_0_31_4 ();
 sg13g2_fill_1 FILLER_0_31_9 ();
 sg13g2_fill_1 FILLER_0_31_75 ();
 sg13g2_fill_1 FILLER_0_31_102 ();
 sg13g2_fill_1 FILLER_0_31_111 ();
 sg13g2_decap_8 FILLER_0_31_147 ();
 sg13g2_decap_8 FILLER_0_31_154 ();
 sg13g2_decap_4 FILLER_0_31_166 ();
 sg13g2_fill_1 FILLER_0_31_170 ();
 sg13g2_fill_2 FILLER_0_31_190 ();
 sg13g2_decap_4 FILLER_0_31_223 ();
 sg13g2_fill_2 FILLER_0_31_227 ();
 sg13g2_decap_8 FILLER_0_31_237 ();
 sg13g2_fill_1 FILLER_0_31_244 ();
 sg13g2_decap_8 FILLER_0_31_249 ();
 sg13g2_decap_4 FILLER_0_31_256 ();
 sg13g2_fill_1 FILLER_0_31_265 ();
 sg13g2_decap_8 FILLER_0_31_302 ();
 sg13g2_fill_1 FILLER_0_31_309 ();
 sg13g2_fill_1 FILLER_0_31_318 ();
 sg13g2_fill_1 FILLER_0_31_327 ();
 sg13g2_decap_4 FILLER_0_31_338 ();
 sg13g2_fill_1 FILLER_0_31_342 ();
 sg13g2_decap_8 FILLER_0_31_351 ();
 sg13g2_decap_4 FILLER_0_31_358 ();
 sg13g2_fill_1 FILLER_0_31_362 ();
 sg13g2_fill_2 FILLER_0_31_381 ();
 sg13g2_decap_4 FILLER_0_31_409 ();
 sg13g2_fill_1 FILLER_0_31_413 ();
 sg13g2_decap_8 FILLER_0_31_418 ();
 sg13g2_decap_4 FILLER_0_31_425 ();
 sg13g2_fill_2 FILLER_0_31_429 ();
 sg13g2_decap_4 FILLER_0_31_435 ();
 sg13g2_fill_2 FILLER_0_31_439 ();
 sg13g2_decap_8 FILLER_0_31_445 ();
 sg13g2_fill_2 FILLER_0_31_452 ();
 sg13g2_fill_1 FILLER_0_31_454 ();
 sg13g2_decap_8 FILLER_0_31_490 ();
 sg13g2_decap_8 FILLER_0_31_497 ();
 sg13g2_decap_8 FILLER_0_31_504 ();
 sg13g2_fill_1 FILLER_0_31_511 ();
 sg13g2_decap_4 FILLER_0_31_520 ();
 sg13g2_fill_1 FILLER_0_31_524 ();
 sg13g2_fill_2 FILLER_0_31_627 ();
 sg13g2_decap_8 FILLER_0_31_634 ();
 sg13g2_decap_8 FILLER_0_31_641 ();
 sg13g2_decap_8 FILLER_0_31_648 ();
 sg13g2_decap_8 FILLER_0_31_655 ();
 sg13g2_decap_8 FILLER_0_31_662 ();
 sg13g2_decap_8 FILLER_0_31_669 ();
 sg13g2_decap_8 FILLER_0_31_676 ();
 sg13g2_decap_8 FILLER_0_31_683 ();
 sg13g2_decap_8 FILLER_0_31_690 ();
 sg13g2_decap_8 FILLER_0_31_697 ();
 sg13g2_decap_8 FILLER_0_31_704 ();
 sg13g2_decap_8 FILLER_0_31_711 ();
 sg13g2_decap_8 FILLER_0_31_718 ();
 sg13g2_decap_8 FILLER_0_31_725 ();
 sg13g2_decap_8 FILLER_0_31_732 ();
 sg13g2_decap_8 FILLER_0_31_739 ();
 sg13g2_decap_4 FILLER_0_31_746 ();
 sg13g2_fill_2 FILLER_0_31_750 ();
 sg13g2_fill_1 FILLER_0_31_756 ();
 sg13g2_decap_8 FILLER_0_31_767 ();
 sg13g2_decap_8 FILLER_0_31_774 ();
 sg13g2_decap_8 FILLER_0_31_781 ();
 sg13g2_decap_4 FILLER_0_31_788 ();
 sg13g2_fill_2 FILLER_0_31_792 ();
 sg13g2_decap_8 FILLER_0_31_824 ();
 sg13g2_decap_8 FILLER_0_31_831 ();
 sg13g2_decap_8 FILLER_0_31_838 ();
 sg13g2_decap_8 FILLER_0_31_845 ();
 sg13g2_decap_8 FILLER_0_31_852 ();
 sg13g2_decap_8 FILLER_0_31_859 ();
 sg13g2_decap_8 FILLER_0_31_866 ();
 sg13g2_decap_8 FILLER_0_31_873 ();
 sg13g2_decap_8 FILLER_0_31_880 ();
 sg13g2_decap_8 FILLER_0_31_887 ();
 sg13g2_decap_8 FILLER_0_31_894 ();
 sg13g2_decap_8 FILLER_0_31_901 ();
 sg13g2_decap_8 FILLER_0_31_908 ();
 sg13g2_decap_8 FILLER_0_31_915 ();
 sg13g2_decap_8 FILLER_0_31_922 ();
 sg13g2_decap_8 FILLER_0_31_929 ();
 sg13g2_decap_4 FILLER_0_31_936 ();
 sg13g2_fill_1 FILLER_0_31_940 ();
 sg13g2_decap_4 FILLER_0_31_951 ();
 sg13g2_fill_2 FILLER_0_31_955 ();
 sg13g2_decap_4 FILLER_0_31_962 ();
 sg13g2_fill_2 FILLER_0_31_966 ();
 sg13g2_fill_2 FILLER_0_31_979 ();
 sg13g2_decap_8 FILLER_0_31_985 ();
 sg13g2_decap_8 FILLER_0_31_992 ();
 sg13g2_decap_4 FILLER_0_31_999 ();
 sg13g2_fill_1 FILLER_0_31_1012 ();
 sg13g2_decap_8 FILLER_0_31_1023 ();
 sg13g2_decap_8 FILLER_0_31_1030 ();
 sg13g2_decap_4 FILLER_0_31_1037 ();
 sg13g2_fill_2 FILLER_0_31_1041 ();
 sg13g2_decap_8 FILLER_0_31_1058 ();
 sg13g2_decap_8 FILLER_0_31_1065 ();
 sg13g2_decap_8 FILLER_0_31_1072 ();
 sg13g2_fill_1 FILLER_0_31_1079 ();
 sg13g2_decap_8 FILLER_0_31_1111 ();
 sg13g2_decap_8 FILLER_0_31_1118 ();
 sg13g2_decap_8 FILLER_0_31_1125 ();
 sg13g2_decap_8 FILLER_0_31_1132 ();
 sg13g2_decap_8 FILLER_0_31_1139 ();
 sg13g2_decap_8 FILLER_0_31_1146 ();
 sg13g2_decap_8 FILLER_0_31_1153 ();
 sg13g2_decap_8 FILLER_0_31_1160 ();
 sg13g2_decap_8 FILLER_0_31_1167 ();
 sg13g2_decap_8 FILLER_0_31_1174 ();
 sg13g2_decap_8 FILLER_0_31_1181 ();
 sg13g2_decap_8 FILLER_0_31_1188 ();
 sg13g2_decap_8 FILLER_0_31_1195 ();
 sg13g2_decap_8 FILLER_0_31_1202 ();
 sg13g2_decap_8 FILLER_0_31_1209 ();
 sg13g2_decap_8 FILLER_0_31_1216 ();
 sg13g2_decap_4 FILLER_0_31_1223 ();
 sg13g2_fill_1 FILLER_0_31_1227 ();
 sg13g2_decap_4 FILLER_0_32_0 ();
 sg13g2_fill_1 FILLER_0_32_4 ();
 sg13g2_fill_2 FILLER_0_32_20 ();
 sg13g2_fill_2 FILLER_0_32_32 ();
 sg13g2_fill_1 FILLER_0_32_34 ();
 sg13g2_fill_2 FILLER_0_32_42 ();
 sg13g2_fill_1 FILLER_0_32_44 ();
 sg13g2_decap_4 FILLER_0_32_65 ();
 sg13g2_fill_2 FILLER_0_32_69 ();
 sg13g2_decap_8 FILLER_0_32_76 ();
 sg13g2_fill_2 FILLER_0_32_83 ();
 sg13g2_decap_8 FILLER_0_32_89 ();
 sg13g2_decap_8 FILLER_0_32_96 ();
 sg13g2_decap_8 FILLER_0_32_103 ();
 sg13g2_fill_2 FILLER_0_32_110 ();
 sg13g2_fill_2 FILLER_0_32_125 ();
 sg13g2_fill_1 FILLER_0_32_127 ();
 sg13g2_decap_8 FILLER_0_32_143 ();
 sg13g2_decap_8 FILLER_0_32_150 ();
 sg13g2_decap_4 FILLER_0_32_157 ();
 sg13g2_fill_1 FILLER_0_32_161 ();
 sg13g2_fill_1 FILLER_0_32_171 ();
 sg13g2_fill_2 FILLER_0_32_182 ();
 sg13g2_decap_4 FILLER_0_32_192 ();
 sg13g2_fill_2 FILLER_0_32_209 ();
 sg13g2_fill_1 FILLER_0_32_211 ();
 sg13g2_decap_4 FILLER_0_32_232 ();
 sg13g2_fill_2 FILLER_0_32_236 ();
 sg13g2_fill_1 FILLER_0_32_242 ();
 sg13g2_decap_4 FILLER_0_32_269 ();
 sg13g2_decap_4 FILLER_0_32_278 ();
 sg13g2_fill_1 FILLER_0_32_282 ();
 sg13g2_fill_2 FILLER_0_32_287 ();
 sg13g2_fill_1 FILLER_0_32_289 ();
 sg13g2_decap_8 FILLER_0_32_294 ();
 sg13g2_decap_8 FILLER_0_32_301 ();
 sg13g2_fill_2 FILLER_0_32_308 ();
 sg13g2_decap_4 FILLER_0_32_315 ();
 sg13g2_decap_8 FILLER_0_32_323 ();
 sg13g2_decap_8 FILLER_0_32_340 ();
 sg13g2_fill_1 FILLER_0_32_347 ();
 sg13g2_fill_1 FILLER_0_32_383 ();
 sg13g2_fill_1 FILLER_0_32_433 ();
 sg13g2_fill_2 FILLER_0_32_465 ();
 sg13g2_fill_1 FILLER_0_32_467 ();
 sg13g2_fill_2 FILLER_0_32_478 ();
 sg13g2_fill_1 FILLER_0_32_480 ();
 sg13g2_decap_8 FILLER_0_32_491 ();
 sg13g2_fill_1 FILLER_0_32_498 ();
 sg13g2_fill_1 FILLER_0_32_534 ();
 sg13g2_decap_8 FILLER_0_32_539 ();
 sg13g2_decap_8 FILLER_0_32_546 ();
 sg13g2_fill_1 FILLER_0_32_553 ();
 sg13g2_fill_2 FILLER_0_32_559 ();
 sg13g2_fill_1 FILLER_0_32_561 ();
 sg13g2_fill_2 FILLER_0_32_566 ();
 sg13g2_fill_1 FILLER_0_32_568 ();
 sg13g2_decap_8 FILLER_0_32_579 ();
 sg13g2_decap_8 FILLER_0_32_586 ();
 sg13g2_decap_8 FILLER_0_32_593 ();
 sg13g2_fill_2 FILLER_0_32_600 ();
 sg13g2_fill_2 FILLER_0_32_628 ();
 sg13g2_decap_8 FILLER_0_32_656 ();
 sg13g2_decap_8 FILLER_0_32_663 ();
 sg13g2_decap_8 FILLER_0_32_722 ();
 sg13g2_decap_8 FILLER_0_32_729 ();
 sg13g2_fill_2 FILLER_0_32_736 ();
 sg13g2_fill_1 FILLER_0_32_741 ();
 sg13g2_decap_8 FILLER_0_32_783 ();
 sg13g2_decap_8 FILLER_0_32_790 ();
 sg13g2_decap_4 FILLER_0_32_797 ();
 sg13g2_fill_2 FILLER_0_32_801 ();
 sg13g2_decap_8 FILLER_0_32_834 ();
 sg13g2_decap_8 FILLER_0_32_841 ();
 sg13g2_decap_8 FILLER_0_32_848 ();
 sg13g2_decap_8 FILLER_0_32_855 ();
 sg13g2_decap_8 FILLER_0_32_862 ();
 sg13g2_decap_8 FILLER_0_32_869 ();
 sg13g2_decap_8 FILLER_0_32_876 ();
 sg13g2_decap_8 FILLER_0_32_883 ();
 sg13g2_decap_8 FILLER_0_32_890 ();
 sg13g2_decap_8 FILLER_0_32_897 ();
 sg13g2_decap_8 FILLER_0_32_904 ();
 sg13g2_decap_8 FILLER_0_32_911 ();
 sg13g2_decap_8 FILLER_0_32_918 ();
 sg13g2_decap_4 FILLER_0_32_925 ();
 sg13g2_fill_1 FILLER_0_32_929 ();
 sg13g2_fill_2 FILLER_0_32_961 ();
 sg13g2_fill_1 FILLER_0_32_963 ();
 sg13g2_decap_8 FILLER_0_32_994 ();
 sg13g2_fill_1 FILLER_0_32_1001 ();
 sg13g2_decap_4 FILLER_0_32_1031 ();
 sg13g2_fill_1 FILLER_0_32_1035 ();
 sg13g2_decap_8 FILLER_0_32_1066 ();
 sg13g2_decap_8 FILLER_0_32_1073 ();
 sg13g2_fill_1 FILLER_0_32_1080 ();
 sg13g2_decap_8 FILLER_0_32_1107 ();
 sg13g2_decap_8 FILLER_0_32_1114 ();
 sg13g2_decap_8 FILLER_0_32_1121 ();
 sg13g2_decap_8 FILLER_0_32_1128 ();
 sg13g2_decap_8 FILLER_0_32_1135 ();
 sg13g2_decap_8 FILLER_0_32_1142 ();
 sg13g2_decap_8 FILLER_0_32_1149 ();
 sg13g2_decap_8 FILLER_0_32_1156 ();
 sg13g2_decap_8 FILLER_0_32_1163 ();
 sg13g2_decap_8 FILLER_0_32_1170 ();
 sg13g2_decap_8 FILLER_0_32_1177 ();
 sg13g2_decap_8 FILLER_0_32_1184 ();
 sg13g2_decap_8 FILLER_0_32_1191 ();
 sg13g2_decap_8 FILLER_0_32_1198 ();
 sg13g2_decap_8 FILLER_0_32_1205 ();
 sg13g2_decap_8 FILLER_0_32_1212 ();
 sg13g2_decap_8 FILLER_0_32_1219 ();
 sg13g2_fill_2 FILLER_0_32_1226 ();
 sg13g2_decap_8 FILLER_0_33_0 ();
 sg13g2_decap_8 FILLER_0_33_47 ();
 sg13g2_fill_2 FILLER_0_33_54 ();
 sg13g2_fill_1 FILLER_0_33_56 ();
 sg13g2_decap_8 FILLER_0_33_61 ();
 sg13g2_fill_2 FILLER_0_33_68 ();
 sg13g2_fill_2 FILLER_0_33_80 ();
 sg13g2_fill_1 FILLER_0_33_82 ();
 sg13g2_fill_1 FILLER_0_33_93 ();
 sg13g2_fill_2 FILLER_0_33_120 ();
 sg13g2_decap_8 FILLER_0_33_153 ();
 sg13g2_fill_2 FILLER_0_33_160 ();
 sg13g2_fill_1 FILLER_0_33_162 ();
 sg13g2_decap_8 FILLER_0_33_189 ();
 sg13g2_decap_8 FILLER_0_33_226 ();
 sg13g2_decap_8 FILLER_0_33_233 ();
 sg13g2_decap_4 FILLER_0_33_240 ();
 sg13g2_fill_1 FILLER_0_33_244 ();
 sg13g2_fill_2 FILLER_0_33_271 ();
 sg13g2_fill_1 FILLER_0_33_273 ();
 sg13g2_decap_8 FILLER_0_33_304 ();
 sg13g2_fill_2 FILLER_0_33_347 ();
 sg13g2_decap_8 FILLER_0_33_379 ();
 sg13g2_decap_4 FILLER_0_33_386 ();
 sg13g2_fill_1 FILLER_0_33_390 ();
 sg13g2_decap_4 FILLER_0_33_417 ();
 sg13g2_fill_1 FILLER_0_33_421 ();
 sg13g2_fill_2 FILLER_0_33_478 ();
 sg13g2_decap_4 FILLER_0_33_523 ();
 sg13g2_fill_1 FILLER_0_33_527 ();
 sg13g2_decap_8 FILLER_0_33_538 ();
 sg13g2_decap_8 FILLER_0_33_545 ();
 sg13g2_decap_8 FILLER_0_33_552 ();
 sg13g2_fill_1 FILLER_0_33_559 ();
 sg13g2_decap_8 FILLER_0_33_570 ();
 sg13g2_decap_8 FILLER_0_33_577 ();
 sg13g2_decap_8 FILLER_0_33_584 ();
 sg13g2_decap_8 FILLER_0_33_591 ();
 sg13g2_fill_1 FILLER_0_33_678 ();
 sg13g2_fill_2 FILLER_0_33_710 ();
 sg13g2_fill_1 FILLER_0_33_751 ();
 sg13g2_fill_1 FILLER_0_33_787 ();
 sg13g2_fill_2 FILLER_0_33_798 ();
 sg13g2_fill_2 FILLER_0_33_805 ();
 sg13g2_fill_2 FILLER_0_33_811 ();
 sg13g2_fill_2 FILLER_0_33_823 ();
 sg13g2_decap_8 FILLER_0_33_859 ();
 sg13g2_decap_8 FILLER_0_33_866 ();
 sg13g2_decap_8 FILLER_0_33_873 ();
 sg13g2_decap_8 FILLER_0_33_880 ();
 sg13g2_decap_8 FILLER_0_33_887 ();
 sg13g2_decap_8 FILLER_0_33_894 ();
 sg13g2_decap_8 FILLER_0_33_901 ();
 sg13g2_decap_8 FILLER_0_33_908 ();
 sg13g2_decap_8 FILLER_0_33_915 ();
 sg13g2_decap_8 FILLER_0_33_922 ();
 sg13g2_decap_4 FILLER_0_33_929 ();
 sg13g2_fill_2 FILLER_0_33_933 ();
 sg13g2_fill_2 FILLER_0_33_1041 ();
 sg13g2_fill_1 FILLER_0_33_1043 ();
 sg13g2_decap_4 FILLER_0_33_1059 ();
 sg13g2_decap_8 FILLER_0_33_1073 ();
 sg13g2_decap_8 FILLER_0_33_1109 ();
 sg13g2_decap_8 FILLER_0_33_1116 ();
 sg13g2_decap_8 FILLER_0_33_1123 ();
 sg13g2_decap_8 FILLER_0_33_1130 ();
 sg13g2_decap_8 FILLER_0_33_1137 ();
 sg13g2_decap_8 FILLER_0_33_1144 ();
 sg13g2_decap_8 FILLER_0_33_1151 ();
 sg13g2_decap_8 FILLER_0_33_1158 ();
 sg13g2_decap_8 FILLER_0_33_1165 ();
 sg13g2_decap_8 FILLER_0_33_1172 ();
 sg13g2_decap_8 FILLER_0_33_1179 ();
 sg13g2_decap_8 FILLER_0_33_1186 ();
 sg13g2_decap_8 FILLER_0_33_1193 ();
 sg13g2_decap_8 FILLER_0_33_1200 ();
 sg13g2_decap_8 FILLER_0_33_1207 ();
 sg13g2_decap_8 FILLER_0_33_1214 ();
 sg13g2_decap_8 FILLER_0_33_1221 ();
 sg13g2_decap_4 FILLER_0_34_0 ();
 sg13g2_decap_8 FILLER_0_34_40 ();
 sg13g2_fill_1 FILLER_0_34_47 ();
 sg13g2_fill_1 FILLER_0_34_53 ();
 sg13g2_fill_1 FILLER_0_34_106 ();
 sg13g2_fill_1 FILLER_0_34_159 ();
 sg13g2_decap_8 FILLER_0_34_190 ();
 sg13g2_fill_1 FILLER_0_34_197 ();
 sg13g2_decap_8 FILLER_0_34_238 ();
 sg13g2_fill_2 FILLER_0_34_245 ();
 sg13g2_fill_1 FILLER_0_34_274 ();
 sg13g2_fill_2 FILLER_0_34_280 ();
 sg13g2_fill_1 FILLER_0_34_282 ();
 sg13g2_decap_8 FILLER_0_34_309 ();
 sg13g2_fill_1 FILLER_0_34_316 ();
 sg13g2_fill_2 FILLER_0_34_348 ();
 sg13g2_decap_8 FILLER_0_34_380 ();
 sg13g2_decap_8 FILLER_0_34_387 ();
 sg13g2_fill_2 FILLER_0_34_394 ();
 sg13g2_fill_1 FILLER_0_34_396 ();
 sg13g2_fill_2 FILLER_0_34_401 ();
 sg13g2_fill_1 FILLER_0_34_403 ();
 sg13g2_fill_2 FILLER_0_34_424 ();
 sg13g2_fill_2 FILLER_0_34_436 ();
 sg13g2_fill_1 FILLER_0_34_438 ();
 sg13g2_decap_4 FILLER_0_34_458 ();
 sg13g2_decap_8 FILLER_0_34_477 ();
 sg13g2_decap_8 FILLER_0_34_484 ();
 sg13g2_fill_2 FILLER_0_34_491 ();
 sg13g2_fill_1 FILLER_0_34_512 ();
 sg13g2_decap_8 FILLER_0_34_523 ();
 sg13g2_decap_4 FILLER_0_34_530 ();
 sg13g2_decap_8 FILLER_0_34_551 ();
 sg13g2_fill_1 FILLER_0_34_558 ();
 sg13g2_decap_8 FILLER_0_34_569 ();
 sg13g2_decap_8 FILLER_0_34_576 ();
 sg13g2_decap_8 FILLER_0_34_583 ();
 sg13g2_decap_8 FILLER_0_34_590 ();
 sg13g2_fill_2 FILLER_0_34_597 ();
 sg13g2_fill_1 FILLER_0_34_599 ();
 sg13g2_fill_2 FILLER_0_34_680 ();
 sg13g2_fill_2 FILLER_0_34_691 ();
 sg13g2_fill_2 FILLER_0_34_703 ();
 sg13g2_fill_1 FILLER_0_34_705 ();
 sg13g2_fill_2 FILLER_0_34_725 ();
 sg13g2_decap_4 FILLER_0_34_757 ();
 sg13g2_fill_1 FILLER_0_34_761 ();
 sg13g2_decap_8 FILLER_0_34_766 ();
 sg13g2_decap_4 FILLER_0_34_773 ();
 sg13g2_fill_2 FILLER_0_34_777 ();
 sg13g2_decap_4 FILLER_0_34_789 ();
 sg13g2_fill_2 FILLER_0_34_793 ();
 sg13g2_fill_2 FILLER_0_34_800 ();
 sg13g2_fill_2 FILLER_0_34_806 ();
 sg13g2_fill_1 FILLER_0_34_808 ();
 sg13g2_fill_1 FILLER_0_34_823 ();
 sg13g2_fill_1 FILLER_0_34_829 ();
 sg13g2_fill_1 FILLER_0_34_856 ();
 sg13g2_fill_2 FILLER_0_34_861 ();
 sg13g2_fill_2 FILLER_0_34_873 ();
 sg13g2_decap_4 FILLER_0_34_880 ();
 sg13g2_fill_2 FILLER_0_34_884 ();
 sg13g2_fill_2 FILLER_0_34_891 ();
 sg13g2_decap_8 FILLER_0_34_905 ();
 sg13g2_decap_8 FILLER_0_34_912 ();
 sg13g2_fill_2 FILLER_0_34_950 ();
 sg13g2_fill_1 FILLER_0_34_977 ();
 sg13g2_decap_8 FILLER_0_34_993 ();
 sg13g2_decap_4 FILLER_0_34_1000 ();
 sg13g2_fill_1 FILLER_0_34_1004 ();
 sg13g2_fill_2 FILLER_0_34_1037 ();
 sg13g2_fill_1 FILLER_0_34_1039 ();
 sg13g2_fill_1 FILLER_0_34_1111 ();
 sg13g2_decap_8 FILLER_0_34_1142 ();
 sg13g2_decap_8 FILLER_0_34_1149 ();
 sg13g2_decap_8 FILLER_0_34_1156 ();
 sg13g2_decap_8 FILLER_0_34_1163 ();
 sg13g2_decap_8 FILLER_0_34_1170 ();
 sg13g2_decap_8 FILLER_0_34_1177 ();
 sg13g2_decap_8 FILLER_0_34_1184 ();
 sg13g2_decap_8 FILLER_0_34_1191 ();
 sg13g2_decap_8 FILLER_0_34_1198 ();
 sg13g2_decap_8 FILLER_0_34_1205 ();
 sg13g2_decap_8 FILLER_0_34_1212 ();
 sg13g2_decap_8 FILLER_0_34_1219 ();
 sg13g2_fill_2 FILLER_0_34_1226 ();
 sg13g2_decap_4 FILLER_0_35_0 ();
 sg13g2_fill_2 FILLER_0_35_13 ();
 sg13g2_fill_1 FILLER_0_35_15 ();
 sg13g2_fill_1 FILLER_0_35_24 ();
 sg13g2_decap_8 FILLER_0_35_35 ();
 sg13g2_decap_4 FILLER_0_35_42 ();
 sg13g2_fill_1 FILLER_0_35_46 ();
 sg13g2_decap_4 FILLER_0_35_82 ();
 sg13g2_fill_1 FILLER_0_35_86 ();
 sg13g2_fill_2 FILLER_0_35_115 ();
 sg13g2_fill_1 FILLER_0_35_127 ();
 sg13g2_fill_1 FILLER_0_35_133 ();
 sg13g2_fill_1 FILLER_0_35_138 ();
 sg13g2_decap_4 FILLER_0_35_161 ();
 sg13g2_fill_1 FILLER_0_35_165 ();
 sg13g2_decap_8 FILLER_0_35_181 ();
 sg13g2_decap_8 FILLER_0_35_188 ();
 sg13g2_decap_8 FILLER_0_35_195 ();
 sg13g2_fill_1 FILLER_0_35_202 ();
 sg13g2_decap_4 FILLER_0_35_208 ();
 sg13g2_fill_1 FILLER_0_35_212 ();
 sg13g2_decap_8 FILLER_0_35_244 ();
 sg13g2_decap_8 FILLER_0_35_251 ();
 sg13g2_decap_4 FILLER_0_35_258 ();
 sg13g2_fill_1 FILLER_0_35_262 ();
 sg13g2_decap_4 FILLER_0_35_270 ();
 sg13g2_decap_8 FILLER_0_35_284 ();
 sg13g2_decap_8 FILLER_0_35_291 ();
 sg13g2_fill_2 FILLER_0_35_298 ();
 sg13g2_fill_1 FILLER_0_35_300 ();
 sg13g2_decap_8 FILLER_0_35_316 ();
 sg13g2_decap_8 FILLER_0_35_327 ();
 sg13g2_decap_8 FILLER_0_35_334 ();
 sg13g2_decap_8 FILLER_0_35_341 ();
 sg13g2_decap_8 FILLER_0_35_382 ();
 sg13g2_fill_2 FILLER_0_35_389 ();
 sg13g2_decap_8 FILLER_0_35_396 ();
 sg13g2_decap_8 FILLER_0_35_403 ();
 sg13g2_decap_8 FILLER_0_35_410 ();
 sg13g2_decap_8 FILLER_0_35_417 ();
 sg13g2_decap_8 FILLER_0_35_424 ();
 sg13g2_decap_8 FILLER_0_35_439 ();
 sg13g2_decap_8 FILLER_0_35_446 ();
 sg13g2_decap_8 FILLER_0_35_453 ();
 sg13g2_decap_8 FILLER_0_35_460 ();
 sg13g2_decap_8 FILLER_0_35_467 ();
 sg13g2_decap_8 FILLER_0_35_474 ();
 sg13g2_decap_8 FILLER_0_35_481 ();
 sg13g2_fill_1 FILLER_0_35_488 ();
 sg13g2_decap_8 FILLER_0_35_515 ();
 sg13g2_decap_8 FILLER_0_35_522 ();
 sg13g2_decap_8 FILLER_0_35_529 ();
 sg13g2_decap_4 FILLER_0_35_536 ();
 sg13g2_fill_1 FILLER_0_35_566 ();
 sg13g2_fill_2 FILLER_0_35_593 ();
 sg13g2_fill_1 FILLER_0_35_600 ();
 sg13g2_fill_2 FILLER_0_35_606 ();
 sg13g2_fill_1 FILLER_0_35_608 ();
 sg13g2_decap_8 FILLER_0_35_622 ();
 sg13g2_decap_8 FILLER_0_35_629 ();
 sg13g2_fill_1 FILLER_0_35_636 ();
 sg13g2_decap_8 FILLER_0_35_641 ();
 sg13g2_fill_1 FILLER_0_35_657 ();
 sg13g2_fill_1 FILLER_0_35_662 ();
 sg13g2_fill_1 FILLER_0_35_673 ();
 sg13g2_fill_2 FILLER_0_35_684 ();
 sg13g2_fill_1 FILLER_0_35_691 ();
 sg13g2_decap_8 FILLER_0_35_702 ();
 sg13g2_decap_4 FILLER_0_35_709 ();
 sg13g2_fill_2 FILLER_0_35_713 ();
 sg13g2_decap_8 FILLER_0_35_719 ();
 sg13g2_fill_2 FILLER_0_35_726 ();
 sg13g2_fill_1 FILLER_0_35_728 ();
 sg13g2_decap_8 FILLER_0_35_753 ();
 sg13g2_fill_2 FILLER_0_35_791 ();
 sg13g2_fill_2 FILLER_0_35_819 ();
 sg13g2_fill_2 FILLER_0_35_831 ();
 sg13g2_decap_8 FILLER_0_35_841 ();
 sg13g2_fill_2 FILLER_0_35_848 ();
 sg13g2_fill_1 FILLER_0_35_850 ();
 sg13g2_decap_8 FILLER_0_35_903 ();
 sg13g2_decap_8 FILLER_0_35_910 ();
 sg13g2_decap_8 FILLER_0_35_917 ();
 sg13g2_decap_8 FILLER_0_35_924 ();
 sg13g2_fill_2 FILLER_0_35_931 ();
 sg13g2_fill_1 FILLER_0_35_933 ();
 sg13g2_decap_8 FILLER_0_35_938 ();
 sg13g2_decap_8 FILLER_0_35_945 ();
 sg13g2_decap_4 FILLER_0_35_952 ();
 sg13g2_fill_1 FILLER_0_35_956 ();
 sg13g2_decap_8 FILLER_0_35_961 ();
 sg13g2_fill_2 FILLER_0_35_968 ();
 sg13g2_fill_1 FILLER_0_35_970 ();
 sg13g2_decap_8 FILLER_0_35_975 ();
 sg13g2_decap_8 FILLER_0_35_982 ();
 sg13g2_decap_8 FILLER_0_35_989 ();
 sg13g2_decap_8 FILLER_0_35_996 ();
 sg13g2_decap_8 FILLER_0_35_1003 ();
 sg13g2_decap_8 FILLER_0_35_1036 ();
 sg13g2_decap_8 FILLER_0_35_1043 ();
 sg13g2_fill_1 FILLER_0_35_1050 ();
 sg13g2_decap_4 FILLER_0_35_1077 ();
 sg13g2_decap_4 FILLER_0_35_1085 ();
 sg13g2_fill_1 FILLER_0_35_1089 ();
 sg13g2_decap_8 FILLER_0_35_1094 ();
 sg13g2_fill_2 FILLER_0_35_1101 ();
 sg13g2_decap_8 FILLER_0_35_1128 ();
 sg13g2_decap_8 FILLER_0_35_1135 ();
 sg13g2_decap_8 FILLER_0_35_1142 ();
 sg13g2_decap_8 FILLER_0_35_1149 ();
 sg13g2_decap_8 FILLER_0_35_1156 ();
 sg13g2_decap_8 FILLER_0_35_1163 ();
 sg13g2_decap_8 FILLER_0_35_1170 ();
 sg13g2_decap_8 FILLER_0_35_1177 ();
 sg13g2_decap_8 FILLER_0_35_1184 ();
 sg13g2_decap_8 FILLER_0_35_1191 ();
 sg13g2_decap_8 FILLER_0_35_1198 ();
 sg13g2_decap_8 FILLER_0_35_1205 ();
 sg13g2_decap_8 FILLER_0_35_1212 ();
 sg13g2_decap_8 FILLER_0_35_1219 ();
 sg13g2_fill_2 FILLER_0_35_1226 ();
 sg13g2_fill_2 FILLER_0_36_0 ();
 sg13g2_fill_1 FILLER_0_36_2 ();
 sg13g2_fill_1 FILLER_0_36_43 ();
 sg13g2_fill_1 FILLER_0_36_49 ();
 sg13g2_fill_2 FILLER_0_36_70 ();
 sg13g2_decap_4 FILLER_0_36_80 ();
 sg13g2_fill_1 FILLER_0_36_84 ();
 sg13g2_decap_8 FILLER_0_36_90 ();
 sg13g2_decap_8 FILLER_0_36_97 ();
 sg13g2_decap_8 FILLER_0_36_104 ();
 sg13g2_decap_4 FILLER_0_36_111 ();
 sg13g2_fill_1 FILLER_0_36_115 ();
 sg13g2_decap_8 FILLER_0_36_120 ();
 sg13g2_decap_8 FILLER_0_36_127 ();
 sg13g2_decap_8 FILLER_0_36_134 ();
 sg13g2_decap_8 FILLER_0_36_141 ();
 sg13g2_decap_4 FILLER_0_36_148 ();
 sg13g2_fill_2 FILLER_0_36_152 ();
 sg13g2_decap_8 FILLER_0_36_184 ();
 sg13g2_decap_8 FILLER_0_36_191 ();
 sg13g2_decap_4 FILLER_0_36_198 ();
 sg13g2_fill_2 FILLER_0_36_202 ();
 sg13g2_fill_1 FILLER_0_36_258 ();
 sg13g2_decap_8 FILLER_0_36_285 ();
 sg13g2_decap_8 FILLER_0_36_292 ();
 sg13g2_decap_8 FILLER_0_36_299 ();
 sg13g2_decap_8 FILLER_0_36_306 ();
 sg13g2_decap_8 FILLER_0_36_313 ();
 sg13g2_decap_8 FILLER_0_36_320 ();
 sg13g2_decap_8 FILLER_0_36_327 ();
 sg13g2_decap_4 FILLER_0_36_334 ();
 sg13g2_fill_1 FILLER_0_36_338 ();
 sg13g2_decap_4 FILLER_0_36_369 ();
 sg13g2_fill_2 FILLER_0_36_373 ();
 sg13g2_fill_2 FILLER_0_36_401 ();
 sg13g2_fill_1 FILLER_0_36_403 ();
 sg13g2_fill_2 FILLER_0_36_430 ();
 sg13g2_fill_2 FILLER_0_36_458 ();
 sg13g2_fill_1 FILLER_0_36_460 ();
 sg13g2_decap_8 FILLER_0_36_465 ();
 sg13g2_decap_8 FILLER_0_36_472 ();
 sg13g2_decap_8 FILLER_0_36_479 ();
 sg13g2_fill_2 FILLER_0_36_486 ();
 sg13g2_fill_1 FILLER_0_36_488 ();
 sg13g2_decap_8 FILLER_0_36_512 ();
 sg13g2_fill_2 FILLER_0_36_519 ();
 sg13g2_decap_8 FILLER_0_36_529 ();
 sg13g2_decap_8 FILLER_0_36_536 ();
 sg13g2_decap_8 FILLER_0_36_543 ();
 sg13g2_decap_4 FILLER_0_36_550 ();
 sg13g2_fill_1 FILLER_0_36_554 ();
 sg13g2_decap_8 FILLER_0_36_622 ();
 sg13g2_decap_8 FILLER_0_36_629 ();
 sg13g2_decap_8 FILLER_0_36_636 ();
 sg13g2_decap_8 FILLER_0_36_643 ();
 sg13g2_decap_8 FILLER_0_36_650 ();
 sg13g2_decap_8 FILLER_0_36_657 ();
 sg13g2_decap_4 FILLER_0_36_664 ();
 sg13g2_fill_2 FILLER_0_36_668 ();
 sg13g2_decap_8 FILLER_0_36_687 ();
 sg13g2_decap_8 FILLER_0_36_694 ();
 sg13g2_decap_8 FILLER_0_36_701 ();
 sg13g2_decap_8 FILLER_0_36_708 ();
 sg13g2_fill_2 FILLER_0_36_715 ();
 sg13g2_fill_1 FILLER_0_36_717 ();
 sg13g2_decap_8 FILLER_0_36_766 ();
 sg13g2_decap_8 FILLER_0_36_773 ();
 sg13g2_decap_8 FILLER_0_36_780 ();
 sg13g2_decap_4 FILLER_0_36_787 ();
 sg13g2_decap_8 FILLER_0_36_827 ();
 sg13g2_decap_8 FILLER_0_36_834 ();
 sg13g2_decap_4 FILLER_0_36_841 ();
 sg13g2_fill_2 FILLER_0_36_876 ();
 sg13g2_decap_8 FILLER_0_36_909 ();
 sg13g2_decap_4 FILLER_0_36_916 ();
 sg13g2_fill_2 FILLER_0_36_920 ();
 sg13g2_decap_8 FILLER_0_36_948 ();
 sg13g2_decap_8 FILLER_0_36_955 ();
 sg13g2_decap_8 FILLER_0_36_962 ();
 sg13g2_decap_8 FILLER_0_36_969 ();
 sg13g2_decap_8 FILLER_0_36_976 ();
 sg13g2_decap_8 FILLER_0_36_983 ();
 sg13g2_decap_8 FILLER_0_36_990 ();
 sg13g2_decap_8 FILLER_0_36_997 ();
 sg13g2_decap_8 FILLER_0_36_1004 ();
 sg13g2_decap_8 FILLER_0_36_1011 ();
 sg13g2_decap_4 FILLER_0_36_1018 ();
 sg13g2_fill_2 FILLER_0_36_1022 ();
 sg13g2_fill_1 FILLER_0_36_1028 ();
 sg13g2_fill_2 FILLER_0_36_1044 ();
 sg13g2_decap_4 FILLER_0_36_1049 ();
 sg13g2_fill_2 FILLER_0_36_1053 ();
 sg13g2_decap_4 FILLER_0_36_1059 ();
 sg13g2_decap_4 FILLER_0_36_1099 ();
 sg13g2_decap_8 FILLER_0_36_1134 ();
 sg13g2_decap_8 FILLER_0_36_1141 ();
 sg13g2_decap_8 FILLER_0_36_1148 ();
 sg13g2_decap_8 FILLER_0_36_1155 ();
 sg13g2_decap_8 FILLER_0_36_1162 ();
 sg13g2_decap_8 FILLER_0_36_1169 ();
 sg13g2_decap_8 FILLER_0_36_1176 ();
 sg13g2_decap_8 FILLER_0_36_1183 ();
 sg13g2_decap_8 FILLER_0_36_1190 ();
 sg13g2_decap_8 FILLER_0_36_1197 ();
 sg13g2_decap_8 FILLER_0_36_1204 ();
 sg13g2_decap_8 FILLER_0_36_1211 ();
 sg13g2_decap_8 FILLER_0_36_1218 ();
 sg13g2_fill_2 FILLER_0_36_1225 ();
 sg13g2_fill_1 FILLER_0_36_1227 ();
 sg13g2_fill_2 FILLER_0_37_67 ();
 sg13g2_decap_8 FILLER_0_37_98 ();
 sg13g2_decap_8 FILLER_0_37_105 ();
 sg13g2_decap_8 FILLER_0_37_112 ();
 sg13g2_decap_8 FILLER_0_37_119 ();
 sg13g2_decap_8 FILLER_0_37_126 ();
 sg13g2_decap_8 FILLER_0_37_133 ();
 sg13g2_decap_8 FILLER_0_37_140 ();
 sg13g2_decap_8 FILLER_0_37_147 ();
 sg13g2_decap_4 FILLER_0_37_154 ();
 sg13g2_fill_1 FILLER_0_37_158 ();
 sg13g2_fill_1 FILLER_0_37_164 ();
 sg13g2_fill_2 FILLER_0_37_175 ();
 sg13g2_fill_2 FILLER_0_37_187 ();
 sg13g2_fill_2 FILLER_0_37_215 ();
 sg13g2_fill_1 FILLER_0_37_221 ();
 sg13g2_fill_1 FILLER_0_37_230 ();
 sg13g2_fill_1 FILLER_0_37_241 ();
 sg13g2_fill_1 FILLER_0_37_268 ();
 sg13g2_decap_8 FILLER_0_37_300 ();
 sg13g2_decap_8 FILLER_0_37_307 ();
 sg13g2_decap_8 FILLER_0_37_314 ();
 sg13g2_decap_8 FILLER_0_37_321 ();
 sg13g2_decap_8 FILLER_0_37_328 ();
 sg13g2_decap_4 FILLER_0_37_335 ();
 sg13g2_fill_1 FILLER_0_37_339 ();
 sg13g2_decap_4 FILLER_0_37_356 ();
 sg13g2_fill_1 FILLER_0_37_360 ();
 sg13g2_decap_8 FILLER_0_37_371 ();
 sg13g2_decap_4 FILLER_0_37_378 ();
 sg13g2_fill_2 FILLER_0_37_386 ();
 sg13g2_fill_1 FILLER_0_37_393 ();
 sg13g2_fill_1 FILLER_0_37_404 ();
 sg13g2_fill_1 FILLER_0_37_410 ();
 sg13g2_fill_2 FILLER_0_37_415 ();
 sg13g2_fill_2 FILLER_0_37_443 ();
 sg13g2_fill_1 FILLER_0_37_445 ();
 sg13g2_fill_2 FILLER_0_37_451 ();
 sg13g2_fill_1 FILLER_0_37_453 ();
 sg13g2_decap_4 FILLER_0_37_480 ();
 sg13g2_fill_1 FILLER_0_37_484 ();
 sg13g2_fill_1 FILLER_0_37_511 ();
 sg13g2_fill_2 FILLER_0_37_517 ();
 sg13g2_fill_2 FILLER_0_37_529 ();
 sg13g2_fill_2 FILLER_0_37_541 ();
 sg13g2_fill_2 FILLER_0_37_574 ();
 sg13g2_fill_1 FILLER_0_37_586 ();
 sg13g2_fill_1 FILLER_0_37_597 ();
 sg13g2_fill_2 FILLER_0_37_608 ();
 sg13g2_decap_8 FILLER_0_37_633 ();
 sg13g2_decap_8 FILLER_0_37_640 ();
 sg13g2_decap_8 FILLER_0_37_647 ();
 sg13g2_fill_2 FILLER_0_37_659 ();
 sg13g2_fill_1 FILLER_0_37_661 ();
 sg13g2_fill_1 FILLER_0_37_696 ();
 sg13g2_decap_8 FILLER_0_37_707 ();
 sg13g2_decap_8 FILLER_0_37_714 ();
 sg13g2_fill_1 FILLER_0_37_730 ();
 sg13g2_fill_1 FILLER_0_37_736 ();
 sg13g2_fill_2 FILLER_0_37_777 ();
 sg13g2_fill_2 FILLER_0_37_784 ();
 sg13g2_fill_1 FILLER_0_37_786 ();
 sg13g2_fill_2 FILLER_0_37_827 ();
 sg13g2_decap_8 FILLER_0_37_834 ();
 sg13g2_decap_8 FILLER_0_37_841 ();
 sg13g2_fill_2 FILLER_0_37_848 ();
 sg13g2_fill_2 FILLER_0_37_854 ();
 sg13g2_fill_1 FILLER_0_37_856 ();
 sg13g2_decap_4 FILLER_0_37_918 ();
 sg13g2_decap_4 FILLER_0_37_954 ();
 sg13g2_fill_1 FILLER_0_37_958 ();
 sg13g2_decap_8 FILLER_0_37_969 ();
 sg13g2_decap_8 FILLER_0_37_976 ();
 sg13g2_decap_8 FILLER_0_37_983 ();
 sg13g2_decap_8 FILLER_0_37_990 ();
 sg13g2_decap_8 FILLER_0_37_997 ();
 sg13g2_decap_8 FILLER_0_37_1004 ();
 sg13g2_decap_4 FILLER_0_37_1011 ();
 sg13g2_decap_4 FILLER_0_37_1059 ();
 sg13g2_fill_2 FILLER_0_37_1063 ();
 sg13g2_decap_8 FILLER_0_37_1093 ();
 sg13g2_decap_8 FILLER_0_37_1130 ();
 sg13g2_decap_8 FILLER_0_37_1137 ();
 sg13g2_decap_8 FILLER_0_37_1144 ();
 sg13g2_decap_8 FILLER_0_37_1151 ();
 sg13g2_decap_8 FILLER_0_37_1158 ();
 sg13g2_decap_8 FILLER_0_37_1165 ();
 sg13g2_decap_8 FILLER_0_37_1172 ();
 sg13g2_decap_8 FILLER_0_37_1179 ();
 sg13g2_decap_8 FILLER_0_37_1186 ();
 sg13g2_decap_8 FILLER_0_37_1193 ();
 sg13g2_decap_8 FILLER_0_37_1200 ();
 sg13g2_decap_8 FILLER_0_37_1207 ();
 sg13g2_decap_8 FILLER_0_37_1214 ();
 sg13g2_decap_8 FILLER_0_37_1221 ();
 sg13g2_decap_4 FILLER_0_38_0 ();
 sg13g2_fill_1 FILLER_0_38_4 ();
 sg13g2_decap_8 FILLER_0_38_35 ();
 sg13g2_fill_1 FILLER_0_38_42 ();
 sg13g2_fill_1 FILLER_0_38_51 ();
 sg13g2_decap_4 FILLER_0_38_65 ();
 sg13g2_fill_2 FILLER_0_38_74 ();
 sg13g2_fill_1 FILLER_0_38_76 ();
 sg13g2_decap_8 FILLER_0_38_112 ();
 sg13g2_decap_8 FILLER_0_38_119 ();
 sg13g2_decap_8 FILLER_0_38_126 ();
 sg13g2_decap_8 FILLER_0_38_133 ();
 sg13g2_decap_8 FILLER_0_38_140 ();
 sg13g2_decap_8 FILLER_0_38_147 ();
 sg13g2_fill_1 FILLER_0_38_185 ();
 sg13g2_fill_2 FILLER_0_38_191 ();
 sg13g2_fill_1 FILLER_0_38_197 ();
 sg13g2_fill_1 FILLER_0_38_202 ();
 sg13g2_decap_8 FILLER_0_38_213 ();
 sg13g2_fill_2 FILLER_0_38_220 ();
 sg13g2_fill_2 FILLER_0_38_226 ();
 sg13g2_fill_1 FILLER_0_38_233 ();
 sg13g2_fill_2 FILLER_0_38_238 ();
 sg13g2_fill_1 FILLER_0_38_240 ();
 sg13g2_fill_1 FILLER_0_38_251 ();
 sg13g2_fill_2 FILLER_0_38_256 ();
 sg13g2_fill_2 FILLER_0_38_263 ();
 sg13g2_fill_2 FILLER_0_38_275 ();
 sg13g2_fill_1 FILLER_0_38_277 ();
 sg13g2_fill_2 FILLER_0_38_292 ();
 sg13g2_fill_2 FILLER_0_38_308 ();
 sg13g2_decap_8 FILLER_0_38_315 ();
 sg13g2_decap_8 FILLER_0_38_322 ();
 sg13g2_decap_8 FILLER_0_38_329 ();
 sg13g2_decap_8 FILLER_0_38_336 ();
 sg13g2_fill_1 FILLER_0_38_343 ();
 sg13g2_fill_1 FILLER_0_38_349 ();
 sg13g2_decap_8 FILLER_0_38_364 ();
 sg13g2_decap_8 FILLER_0_38_371 ();
 sg13g2_fill_1 FILLER_0_38_378 ();
 sg13g2_decap_8 FILLER_0_38_384 ();
 sg13g2_fill_2 FILLER_0_38_401 ();
 sg13g2_fill_1 FILLER_0_38_403 ();
 sg13g2_fill_2 FILLER_0_38_414 ();
 sg13g2_fill_1 FILLER_0_38_416 ();
 sg13g2_fill_2 FILLER_0_38_427 ();
 sg13g2_fill_1 FILLER_0_38_439 ();
 sg13g2_fill_1 FILLER_0_38_450 ();
 sg13g2_fill_2 FILLER_0_38_460 ();
 sg13g2_fill_2 FILLER_0_38_492 ();
 sg13g2_fill_1 FILLER_0_38_498 ();
 sg13g2_decap_8 FILLER_0_38_549 ();
 sg13g2_decap_8 FILLER_0_38_560 ();
 sg13g2_fill_1 FILLER_0_38_567 ();
 sg13g2_fill_1 FILLER_0_38_580 ();
 sg13g2_fill_2 FILLER_0_38_585 ();
 sg13g2_decap_8 FILLER_0_38_630 ();
 sg13g2_decap_4 FILLER_0_38_637 ();
 sg13g2_fill_1 FILLER_0_38_641 ();
 sg13g2_decap_8 FILLER_0_38_651 ();
 sg13g2_decap_8 FILLER_0_38_658 ();
 sg13g2_decap_4 FILLER_0_38_665 ();
 sg13g2_fill_1 FILLER_0_38_669 ();
 sg13g2_fill_2 FILLER_0_38_725 ();
 sg13g2_fill_1 FILLER_0_38_727 ();
 sg13g2_decap_4 FILLER_0_38_738 ();
 sg13g2_fill_1 FILLER_0_38_742 ();
 sg13g2_fill_1 FILLER_0_38_788 ();
 sg13g2_decap_8 FILLER_0_38_819 ();
 sg13g2_fill_1 FILLER_0_38_831 ();
 sg13g2_decap_8 FILLER_0_38_858 ();
 sg13g2_decap_4 FILLER_0_38_865 ();
 sg13g2_fill_1 FILLER_0_38_882 ();
 sg13g2_fill_2 FILLER_0_38_887 ();
 sg13g2_fill_1 FILLER_0_38_889 ();
 sg13g2_fill_1 FILLER_0_38_926 ();
 sg13g2_fill_1 FILLER_0_38_934 ();
 sg13g2_fill_1 FILLER_0_38_965 ();
 sg13g2_decap_8 FILLER_0_38_971 ();
 sg13g2_decap_8 FILLER_0_38_978 ();
 sg13g2_decap_8 FILLER_0_38_985 ();
 sg13g2_decap_8 FILLER_0_38_992 ();
 sg13g2_decap_8 FILLER_0_38_999 ();
 sg13g2_decap_8 FILLER_0_38_1006 ();
 sg13g2_fill_2 FILLER_0_38_1013 ();
 sg13g2_decap_4 FILLER_0_38_1020 ();
 sg13g2_fill_1 FILLER_0_38_1024 ();
 sg13g2_fill_1 FILLER_0_38_1030 ();
 sg13g2_fill_1 FILLER_0_38_1036 ();
 sg13g2_fill_1 FILLER_0_38_1063 ();
 sg13g2_fill_1 FILLER_0_38_1074 ();
 sg13g2_decap_8 FILLER_0_38_1101 ();
 sg13g2_decap_8 FILLER_0_38_1134 ();
 sg13g2_decap_8 FILLER_0_38_1141 ();
 sg13g2_decap_8 FILLER_0_38_1148 ();
 sg13g2_decap_8 FILLER_0_38_1155 ();
 sg13g2_decap_8 FILLER_0_38_1162 ();
 sg13g2_decap_8 FILLER_0_38_1169 ();
 sg13g2_decap_8 FILLER_0_38_1176 ();
 sg13g2_decap_8 FILLER_0_38_1183 ();
 sg13g2_decap_8 FILLER_0_38_1190 ();
 sg13g2_decap_8 FILLER_0_38_1197 ();
 sg13g2_decap_8 FILLER_0_38_1204 ();
 sg13g2_decap_8 FILLER_0_38_1211 ();
 sg13g2_decap_8 FILLER_0_38_1218 ();
 sg13g2_fill_2 FILLER_0_38_1225 ();
 sg13g2_fill_1 FILLER_0_38_1227 ();
 sg13g2_decap_8 FILLER_0_39_0 ();
 sg13g2_decap_8 FILLER_0_39_7 ();
 sg13g2_fill_1 FILLER_0_39_14 ();
 sg13g2_fill_2 FILLER_0_39_23 ();
 sg13g2_decap_8 FILLER_0_39_30 ();
 sg13g2_fill_2 FILLER_0_39_37 ();
 sg13g2_fill_2 FILLER_0_39_86 ();
 sg13g2_decap_4 FILLER_0_39_124 ();
 sg13g2_decap_8 FILLER_0_39_133 ();
 sg13g2_decap_8 FILLER_0_39_140 ();
 sg13g2_decap_8 FILLER_0_39_147 ();
 sg13g2_decap_8 FILLER_0_39_154 ();
 sg13g2_fill_2 FILLER_0_39_161 ();
 sg13g2_fill_2 FILLER_0_39_175 ();
 sg13g2_fill_2 FILLER_0_39_182 ();
 sg13g2_decap_8 FILLER_0_39_230 ();
 sg13g2_decap_8 FILLER_0_39_237 ();
 sg13g2_decap_8 FILLER_0_39_244 ();
 sg13g2_decap_8 FILLER_0_39_251 ();
 sg13g2_decap_8 FILLER_0_39_258 ();
 sg13g2_decap_8 FILLER_0_39_265 ();
 sg13g2_decap_8 FILLER_0_39_272 ();
 sg13g2_decap_8 FILLER_0_39_279 ();
 sg13g2_fill_2 FILLER_0_39_286 ();
 sg13g2_decap_4 FILLER_0_39_314 ();
 sg13g2_fill_1 FILLER_0_39_318 ();
 sg13g2_decap_8 FILLER_0_39_328 ();
 sg13g2_fill_2 FILLER_0_39_335 ();
 sg13g2_decap_8 FILLER_0_39_368 ();
 sg13g2_decap_4 FILLER_0_39_375 ();
 sg13g2_decap_8 FILLER_0_39_409 ();
 sg13g2_decap_8 FILLER_0_39_416 ();
 sg13g2_fill_1 FILLER_0_39_423 ();
 sg13g2_decap_8 FILLER_0_39_428 ();
 sg13g2_fill_2 FILLER_0_39_435 ();
 sg13g2_fill_1 FILLER_0_39_437 ();
 sg13g2_fill_2 FILLER_0_39_447 ();
 sg13g2_fill_1 FILLER_0_39_449 ();
 sg13g2_fill_2 FILLER_0_39_465 ();
 sg13g2_decap_8 FILLER_0_39_482 ();
 sg13g2_decap_8 FILLER_0_39_489 ();
 sg13g2_decap_4 FILLER_0_39_496 ();
 sg13g2_fill_1 FILLER_0_39_500 ();
 sg13g2_fill_2 FILLER_0_39_505 ();
 sg13g2_fill_1 FILLER_0_39_507 ();
 sg13g2_fill_2 FILLER_0_39_512 ();
 sg13g2_fill_1 FILLER_0_39_514 ();
 sg13g2_decap_4 FILLER_0_39_519 ();
 sg13g2_fill_2 FILLER_0_39_523 ();
 sg13g2_fill_1 FILLER_0_39_551 ();
 sg13g2_decap_8 FILLER_0_39_562 ();
 sg13g2_fill_2 FILLER_0_39_569 ();
 sg13g2_decap_8 FILLER_0_39_575 ();
 sg13g2_decap_8 FILLER_0_39_582 ();
 sg13g2_fill_2 FILLER_0_39_589 ();
 sg13g2_fill_1 FILLER_0_39_591 ();
 sg13g2_fill_1 FILLER_0_39_626 ();
 sg13g2_decap_4 FILLER_0_39_632 ();
 sg13g2_fill_2 FILLER_0_39_636 ();
 sg13g2_fill_1 FILLER_0_39_664 ();
 sg13g2_fill_1 FILLER_0_39_696 ();
 sg13g2_decap_4 FILLER_0_39_741 ();
 sg13g2_fill_1 FILLER_0_39_745 ();
 sg13g2_decap_8 FILLER_0_39_765 ();
 sg13g2_decap_8 FILLER_0_39_772 ();
 sg13g2_decap_4 FILLER_0_39_779 ();
 sg13g2_fill_1 FILLER_0_39_783 ();
 sg13g2_decap_8 FILLER_0_39_792 ();
 sg13g2_decap_4 FILLER_0_39_799 ();
 sg13g2_fill_2 FILLER_0_39_834 ();
 sg13g2_fill_1 FILLER_0_39_836 ();
 sg13g2_fill_2 FILLER_0_39_873 ();
 sg13g2_decap_4 FILLER_0_39_880 ();
 sg13g2_fill_1 FILLER_0_39_884 ();
 sg13g2_decap_4 FILLER_0_39_889 ();
 sg13g2_fill_1 FILLER_0_39_893 ();
 sg13g2_fill_1 FILLER_0_39_898 ();
 sg13g2_fill_2 FILLER_0_39_904 ();
 sg13g2_fill_2 FILLER_0_39_910 ();
 sg13g2_decap_8 FILLER_0_39_932 ();
 sg13g2_fill_1 FILLER_0_39_970 ();
 sg13g2_decap_8 FILLER_0_39_979 ();
 sg13g2_decap_8 FILLER_0_39_986 ();
 sg13g2_decap_8 FILLER_0_39_993 ();
 sg13g2_decap_8 FILLER_0_39_1000 ();
 sg13g2_decap_8 FILLER_0_39_1007 ();
 sg13g2_decap_8 FILLER_0_39_1014 ();
 sg13g2_fill_2 FILLER_0_39_1021 ();
 sg13g2_fill_1 FILLER_0_39_1023 ();
 sg13g2_decap_4 FILLER_0_39_1081 ();
 sg13g2_fill_2 FILLER_0_39_1085 ();
 sg13g2_fill_1 FILLER_0_39_1097 ();
 sg13g2_decap_8 FILLER_0_39_1106 ();
 sg13g2_fill_1 FILLER_0_39_1113 ();
 sg13g2_decap_8 FILLER_0_39_1144 ();
 sg13g2_decap_8 FILLER_0_39_1151 ();
 sg13g2_decap_8 FILLER_0_39_1158 ();
 sg13g2_decap_8 FILLER_0_39_1165 ();
 sg13g2_decap_8 FILLER_0_39_1172 ();
 sg13g2_decap_8 FILLER_0_39_1179 ();
 sg13g2_decap_8 FILLER_0_39_1186 ();
 sg13g2_decap_8 FILLER_0_39_1193 ();
 sg13g2_decap_8 FILLER_0_39_1200 ();
 sg13g2_decap_8 FILLER_0_39_1207 ();
 sg13g2_decap_8 FILLER_0_39_1214 ();
 sg13g2_decap_8 FILLER_0_39_1221 ();
 sg13g2_decap_8 FILLER_0_40_0 ();
 sg13g2_decap_8 FILLER_0_40_7 ();
 sg13g2_decap_8 FILLER_0_40_14 ();
 sg13g2_decap_8 FILLER_0_40_21 ();
 sg13g2_decap_8 FILLER_0_40_28 ();
 sg13g2_decap_8 FILLER_0_40_35 ();
 sg13g2_decap_8 FILLER_0_40_42 ();
 sg13g2_decap_4 FILLER_0_40_49 ();
 sg13g2_fill_2 FILLER_0_40_61 ();
 sg13g2_fill_1 FILLER_0_40_63 ();
 sg13g2_fill_1 FILLER_0_40_111 ();
 sg13g2_decap_8 FILLER_0_40_116 ();
 sg13g2_decap_8 FILLER_0_40_123 ();
 sg13g2_decap_8 FILLER_0_40_130 ();
 sg13g2_decap_8 FILLER_0_40_137 ();
 sg13g2_decap_8 FILLER_0_40_144 ();
 sg13g2_decap_8 FILLER_0_40_151 ();
 sg13g2_decap_8 FILLER_0_40_158 ();
 sg13g2_decap_8 FILLER_0_40_169 ();
 sg13g2_decap_8 FILLER_0_40_176 ();
 sg13g2_fill_1 FILLER_0_40_199 ();
 sg13g2_fill_2 FILLER_0_40_256 ();
 sg13g2_fill_1 FILLER_0_40_258 ();
 sg13g2_decap_4 FILLER_0_40_294 ();
 sg13g2_fill_2 FILLER_0_40_298 ();
 sg13g2_fill_2 FILLER_0_40_310 ();
 sg13g2_fill_2 FILLER_0_40_317 ();
 sg13g2_decap_4 FILLER_0_40_345 ();
 sg13g2_decap_4 FILLER_0_40_359 ();
 sg13g2_decap_8 FILLER_0_40_418 ();
 sg13g2_decap_8 FILLER_0_40_425 ();
 sg13g2_decap_8 FILLER_0_40_432 ();
 sg13g2_decap_8 FILLER_0_40_439 ();
 sg13g2_decap_8 FILLER_0_40_446 ();
 sg13g2_decap_8 FILLER_0_40_453 ();
 sg13g2_decap_8 FILLER_0_40_460 ();
 sg13g2_decap_8 FILLER_0_40_467 ();
 sg13g2_decap_4 FILLER_0_40_474 ();
 sg13g2_fill_1 FILLER_0_40_478 ();
 sg13g2_decap_4 FILLER_0_40_505 ();
 sg13g2_fill_1 FILLER_0_40_509 ();
 sg13g2_decap_8 FILLER_0_40_515 ();
 sg13g2_decap_4 FILLER_0_40_522 ();
 sg13g2_fill_2 FILLER_0_40_526 ();
 sg13g2_decap_4 FILLER_0_40_613 ();
 sg13g2_fill_2 FILLER_0_40_617 ();
 sg13g2_decap_8 FILLER_0_40_629 ();
 sg13g2_fill_1 FILLER_0_40_636 ();
 sg13g2_decap_8 FILLER_0_40_647 ();
 sg13g2_decap_8 FILLER_0_40_654 ();
 sg13g2_fill_2 FILLER_0_40_661 ();
 sg13g2_fill_1 FILLER_0_40_671 ();
 sg13g2_fill_1 FILLER_0_40_676 ();
 sg13g2_decap_4 FILLER_0_40_701 ();
 sg13g2_fill_2 FILLER_0_40_715 ();
 sg13g2_decap_4 FILLER_0_40_743 ();
 sg13g2_fill_1 FILLER_0_40_747 ();
 sg13g2_decap_8 FILLER_0_40_774 ();
 sg13g2_decap_8 FILLER_0_40_781 ();
 sg13g2_decap_8 FILLER_0_40_788 ();
 sg13g2_decap_8 FILLER_0_40_795 ();
 sg13g2_decap_8 FILLER_0_40_802 ();
 sg13g2_fill_2 FILLER_0_40_878 ();
 sg13g2_decap_8 FILLER_0_40_890 ();
 sg13g2_decap_4 FILLER_0_40_932 ();
 sg13g2_fill_1 FILLER_0_40_936 ();
 sg13g2_decap_8 FILLER_0_40_982 ();
 sg13g2_decap_8 FILLER_0_40_989 ();
 sg13g2_fill_2 FILLER_0_40_1020 ();
 sg13g2_fill_1 FILLER_0_40_1022 ();
 sg13g2_decap_8 FILLER_0_40_1055 ();
 sg13g2_fill_1 FILLER_0_40_1062 ();
 sg13g2_decap_8 FILLER_0_40_1103 ();
 sg13g2_fill_1 FILLER_0_40_1110 ();
 sg13g2_fill_1 FILLER_0_40_1126 ();
 sg13g2_decap_8 FILLER_0_40_1131 ();
 sg13g2_decap_8 FILLER_0_40_1138 ();
 sg13g2_decap_8 FILLER_0_40_1145 ();
 sg13g2_decap_8 FILLER_0_40_1152 ();
 sg13g2_decap_8 FILLER_0_40_1159 ();
 sg13g2_decap_8 FILLER_0_40_1166 ();
 sg13g2_decap_8 FILLER_0_40_1173 ();
 sg13g2_decap_8 FILLER_0_40_1180 ();
 sg13g2_decap_8 FILLER_0_40_1187 ();
 sg13g2_decap_8 FILLER_0_40_1194 ();
 sg13g2_decap_8 FILLER_0_40_1201 ();
 sg13g2_decap_8 FILLER_0_40_1208 ();
 sg13g2_decap_8 FILLER_0_40_1215 ();
 sg13g2_decap_4 FILLER_0_40_1222 ();
 sg13g2_fill_2 FILLER_0_40_1226 ();
 sg13g2_decap_8 FILLER_0_41_0 ();
 sg13g2_decap_8 FILLER_0_41_7 ();
 sg13g2_decap_8 FILLER_0_41_14 ();
 sg13g2_decap_8 FILLER_0_41_21 ();
 sg13g2_decap_8 FILLER_0_41_28 ();
 sg13g2_decap_8 FILLER_0_41_35 ();
 sg13g2_decap_8 FILLER_0_41_42 ();
 sg13g2_decap_4 FILLER_0_41_49 ();
 sg13g2_fill_2 FILLER_0_41_53 ();
 sg13g2_decap_8 FILLER_0_41_59 ();
 sg13g2_fill_2 FILLER_0_41_66 ();
 sg13g2_fill_1 FILLER_0_41_68 ();
 sg13g2_decap_8 FILLER_0_41_73 ();
 sg13g2_fill_1 FILLER_0_41_80 ();
 sg13g2_decap_4 FILLER_0_41_106 ();
 sg13g2_fill_1 FILLER_0_41_120 ();
 sg13g2_decap_8 FILLER_0_41_131 ();
 sg13g2_decap_8 FILLER_0_41_138 ();
 sg13g2_decap_8 FILLER_0_41_145 ();
 sg13g2_decap_8 FILLER_0_41_152 ();
 sg13g2_decap_8 FILLER_0_41_159 ();
 sg13g2_decap_8 FILLER_0_41_166 ();
 sg13g2_decap_8 FILLER_0_41_173 ();
 sg13g2_decap_8 FILLER_0_41_180 ();
 sg13g2_decap_8 FILLER_0_41_187 ();
 sg13g2_fill_2 FILLER_0_41_194 ();
 sg13g2_fill_1 FILLER_0_41_196 ();
 sg13g2_decap_8 FILLER_0_41_222 ();
 sg13g2_decap_4 FILLER_0_41_229 ();
 sg13g2_fill_1 FILLER_0_41_233 ();
 sg13g2_fill_1 FILLER_0_41_242 ();
 sg13g2_fill_2 FILLER_0_41_300 ();
 sg13g2_decap_4 FILLER_0_41_332 ();
 sg13g2_fill_2 FILLER_0_41_336 ();
 sg13g2_fill_1 FILLER_0_41_343 ();
 sg13g2_fill_2 FILLER_0_41_404 ();
 sg13g2_fill_1 FILLER_0_41_437 ();
 sg13g2_fill_1 FILLER_0_41_442 ();
 sg13g2_fill_2 FILLER_0_41_453 ();
 sg13g2_fill_1 FILLER_0_41_455 ();
 sg13g2_decap_4 FILLER_0_41_491 ();
 sg13g2_fill_1 FILLER_0_41_495 ();
 sg13g2_decap_4 FILLER_0_41_522 ();
 sg13g2_fill_1 FILLER_0_41_526 ();
 sg13g2_fill_2 FILLER_0_41_532 ();
 sg13g2_fill_1 FILLER_0_41_556 ();
 sg13g2_decap_8 FILLER_0_41_619 ();
 sg13g2_fill_2 FILLER_0_41_626 ();
 sg13g2_decap_8 FILLER_0_41_654 ();
 sg13g2_fill_1 FILLER_0_41_661 ();
 sg13g2_decap_8 FILLER_0_41_693 ();
 sg13g2_decap_8 FILLER_0_41_700 ();
 sg13g2_fill_2 FILLER_0_41_707 ();
 sg13g2_fill_1 FILLER_0_41_709 ();
 sg13g2_fill_1 FILLER_0_41_715 ();
 sg13g2_decap_8 FILLER_0_41_730 ();
 sg13g2_decap_8 FILLER_0_41_737 ();
 sg13g2_decap_4 FILLER_0_41_744 ();
 sg13g2_fill_2 FILLER_0_41_748 ();
 sg13g2_fill_1 FILLER_0_41_768 ();
 sg13g2_decap_8 FILLER_0_41_795 ();
 sg13g2_decap_8 FILLER_0_41_802 ();
 sg13g2_decap_8 FILLER_0_41_809 ();
 sg13g2_decap_8 FILLER_0_41_816 ();
 sg13g2_decap_8 FILLER_0_41_823 ();
 sg13g2_decap_8 FILLER_0_41_830 ();
 sg13g2_decap_8 FILLER_0_41_837 ();
 sg13g2_fill_2 FILLER_0_41_844 ();
 sg13g2_fill_1 FILLER_0_41_850 ();
 sg13g2_fill_2 FILLER_0_41_881 ();
 sg13g2_fill_1 FILLER_0_41_883 ();
 sg13g2_decap_8 FILLER_0_41_889 ();
 sg13g2_fill_1 FILLER_0_41_896 ();
 sg13g2_decap_4 FILLER_0_41_901 ();
 sg13g2_decap_4 FILLER_0_41_931 ();
 sg13g2_fill_1 FILLER_0_41_935 ();
 sg13g2_decap_8 FILLER_0_41_967 ();
 sg13g2_fill_2 FILLER_0_41_974 ();
 sg13g2_fill_1 FILLER_0_41_980 ();
 sg13g2_fill_2 FILLER_0_41_1007 ();
 sg13g2_fill_1 FILLER_0_41_1009 ();
 sg13g2_decap_8 FILLER_0_41_1046 ();
 sg13g2_decap_8 FILLER_0_41_1053 ();
 sg13g2_decap_8 FILLER_0_41_1060 ();
 sg13g2_decap_8 FILLER_0_41_1067 ();
 sg13g2_fill_1 FILLER_0_41_1074 ();
 sg13g2_decap_8 FILLER_0_41_1131 ();
 sg13g2_decap_8 FILLER_0_41_1138 ();
 sg13g2_decap_8 FILLER_0_41_1145 ();
 sg13g2_decap_8 FILLER_0_41_1152 ();
 sg13g2_decap_8 FILLER_0_41_1159 ();
 sg13g2_decap_8 FILLER_0_41_1166 ();
 sg13g2_decap_8 FILLER_0_41_1173 ();
 sg13g2_decap_8 FILLER_0_41_1180 ();
 sg13g2_decap_8 FILLER_0_41_1187 ();
 sg13g2_decap_8 FILLER_0_41_1194 ();
 sg13g2_decap_8 FILLER_0_41_1201 ();
 sg13g2_decap_8 FILLER_0_41_1208 ();
 sg13g2_decap_8 FILLER_0_41_1215 ();
 sg13g2_decap_4 FILLER_0_41_1222 ();
 sg13g2_fill_2 FILLER_0_41_1226 ();
 sg13g2_decap_8 FILLER_0_42_0 ();
 sg13g2_decap_8 FILLER_0_42_7 ();
 sg13g2_decap_8 FILLER_0_42_14 ();
 sg13g2_decap_8 FILLER_0_42_21 ();
 sg13g2_decap_8 FILLER_0_42_28 ();
 sg13g2_decap_8 FILLER_0_42_35 ();
 sg13g2_decap_4 FILLER_0_42_42 ();
 sg13g2_fill_1 FILLER_0_42_99 ();
 sg13g2_fill_2 FILLER_0_42_126 ();
 sg13g2_decap_8 FILLER_0_42_132 ();
 sg13g2_decap_8 FILLER_0_42_139 ();
 sg13g2_decap_8 FILLER_0_42_146 ();
 sg13g2_decap_8 FILLER_0_42_153 ();
 sg13g2_decap_8 FILLER_0_42_160 ();
 sg13g2_decap_8 FILLER_0_42_167 ();
 sg13g2_decap_8 FILLER_0_42_174 ();
 sg13g2_decap_8 FILLER_0_42_181 ();
 sg13g2_decap_8 FILLER_0_42_223 ();
 sg13g2_decap_4 FILLER_0_42_230 ();
 sg13g2_fill_2 FILLER_0_42_234 ();
 sg13g2_fill_1 FILLER_0_42_265 ();
 sg13g2_fill_2 FILLER_0_42_271 ();
 sg13g2_fill_1 FILLER_0_42_283 ();
 sg13g2_fill_2 FILLER_0_42_294 ();
 sg13g2_fill_1 FILLER_0_42_311 ();
 sg13g2_decap_8 FILLER_0_42_316 ();
 sg13g2_decap_8 FILLER_0_42_323 ();
 sg13g2_decap_4 FILLER_0_42_330 ();
 sg13g2_decap_8 FILLER_0_42_338 ();
 sg13g2_decap_8 FILLER_0_42_345 ();
 sg13g2_fill_1 FILLER_0_42_352 ();
 sg13g2_decap_4 FILLER_0_42_357 ();
 sg13g2_decap_8 FILLER_0_42_366 ();
 sg13g2_fill_2 FILLER_0_42_373 ();
 sg13g2_fill_1 FILLER_0_42_375 ();
 sg13g2_fill_1 FILLER_0_42_399 ();
 sg13g2_fill_1 FILLER_0_42_430 ();
 sg13g2_fill_1 FILLER_0_42_461 ();
 sg13g2_decap_4 FILLER_0_42_470 ();
 sg13g2_fill_2 FILLER_0_42_479 ();
 sg13g2_fill_1 FILLER_0_42_481 ();
 sg13g2_fill_1 FILLER_0_42_502 ();
 sg13g2_fill_1 FILLER_0_42_507 ();
 sg13g2_decap_8 FILLER_0_42_518 ();
 sg13g2_fill_1 FILLER_0_42_525 ();
 sg13g2_decap_8 FILLER_0_42_536 ();
 sg13g2_fill_1 FILLER_0_42_576 ();
 sg13g2_fill_1 FILLER_0_42_587 ();
 sg13g2_fill_1 FILLER_0_42_593 ();
 sg13g2_decap_8 FILLER_0_42_608 ();
 sg13g2_decap_8 FILLER_0_42_615 ();
 sg13g2_decap_4 FILLER_0_42_622 ();
 sg13g2_fill_1 FILLER_0_42_626 ();
 sg13g2_fill_1 FILLER_0_42_632 ();
 sg13g2_fill_2 FILLER_0_42_665 ();
 sg13g2_fill_1 FILLER_0_42_676 ();
 sg13g2_decap_8 FILLER_0_42_687 ();
 sg13g2_decap_8 FILLER_0_42_694 ();
 sg13g2_fill_1 FILLER_0_42_701 ();
 sg13g2_fill_2 FILLER_0_42_762 ();
 sg13g2_fill_1 FILLER_0_42_769 ();
 sg13g2_decap_8 FILLER_0_42_774 ();
 sg13g2_decap_8 FILLER_0_42_781 ();
 sg13g2_decap_8 FILLER_0_42_788 ();
 sg13g2_decap_8 FILLER_0_42_795 ();
 sg13g2_decap_8 FILLER_0_42_802 ();
 sg13g2_decap_8 FILLER_0_42_809 ();
 sg13g2_decap_4 FILLER_0_42_816 ();
 sg13g2_fill_2 FILLER_0_42_820 ();
 sg13g2_decap_8 FILLER_0_42_831 ();
 sg13g2_decap_8 FILLER_0_42_838 ();
 sg13g2_decap_8 FILLER_0_42_845 ();
 sg13g2_fill_2 FILLER_0_42_852 ();
 sg13g2_fill_1 FILLER_0_42_854 ();
 sg13g2_decap_4 FILLER_0_42_907 ();
 sg13g2_fill_2 FILLER_0_42_915 ();
 sg13g2_decap_4 FILLER_0_42_922 ();
 sg13g2_fill_1 FILLER_0_42_956 ();
 sg13g2_fill_2 FILLER_0_42_962 ();
 sg13g2_decap_8 FILLER_0_42_1005 ();
 sg13g2_decap_4 FILLER_0_42_1012 ();
 sg13g2_fill_1 FILLER_0_42_1016 ();
 sg13g2_decap_4 FILLER_0_42_1021 ();
 sg13g2_fill_1 FILLER_0_42_1025 ();
 sg13g2_decap_8 FILLER_0_42_1057 ();
 sg13g2_decap_8 FILLER_0_42_1064 ();
 sg13g2_decap_8 FILLER_0_42_1071 ();
 sg13g2_fill_2 FILLER_0_42_1078 ();
 sg13g2_fill_1 FILLER_0_42_1080 ();
 sg13g2_decap_4 FILLER_0_42_1090 ();
 sg13g2_fill_1 FILLER_0_42_1094 ();
 sg13g2_fill_1 FILLER_0_42_1120 ();
 sg13g2_decap_8 FILLER_0_42_1125 ();
 sg13g2_decap_8 FILLER_0_42_1132 ();
 sg13g2_decap_8 FILLER_0_42_1139 ();
 sg13g2_decap_8 FILLER_0_42_1146 ();
 sg13g2_decap_8 FILLER_0_42_1153 ();
 sg13g2_decap_8 FILLER_0_42_1160 ();
 sg13g2_decap_8 FILLER_0_42_1167 ();
 sg13g2_decap_8 FILLER_0_42_1174 ();
 sg13g2_decap_8 FILLER_0_42_1181 ();
 sg13g2_decap_8 FILLER_0_42_1188 ();
 sg13g2_decap_8 FILLER_0_42_1195 ();
 sg13g2_decap_8 FILLER_0_42_1202 ();
 sg13g2_decap_8 FILLER_0_42_1209 ();
 sg13g2_decap_8 FILLER_0_42_1216 ();
 sg13g2_decap_4 FILLER_0_42_1223 ();
 sg13g2_fill_1 FILLER_0_42_1227 ();
 sg13g2_decap_8 FILLER_0_43_0 ();
 sg13g2_decap_8 FILLER_0_43_7 ();
 sg13g2_decap_8 FILLER_0_43_14 ();
 sg13g2_decap_8 FILLER_0_43_21 ();
 sg13g2_decap_8 FILLER_0_43_28 ();
 sg13g2_decap_8 FILLER_0_43_35 ();
 sg13g2_decap_8 FILLER_0_43_42 ();
 sg13g2_decap_4 FILLER_0_43_49 ();
 sg13g2_fill_1 FILLER_0_43_53 ();
 sg13g2_decap_8 FILLER_0_43_130 ();
 sg13g2_decap_8 FILLER_0_43_137 ();
 sg13g2_decap_8 FILLER_0_43_144 ();
 sg13g2_decap_8 FILLER_0_43_151 ();
 sg13g2_decap_8 FILLER_0_43_158 ();
 sg13g2_decap_8 FILLER_0_43_165 ();
 sg13g2_decap_8 FILLER_0_43_172 ();
 sg13g2_fill_2 FILLER_0_43_179 ();
 sg13g2_fill_1 FILLER_0_43_181 ();
 sg13g2_decap_8 FILLER_0_43_212 ();
 sg13g2_decap_8 FILLER_0_43_219 ();
 sg13g2_decap_4 FILLER_0_43_226 ();
 sg13g2_fill_2 FILLER_0_43_230 ();
 sg13g2_fill_2 FILLER_0_43_252 ();
 sg13g2_fill_1 FILLER_0_43_265 ();
 sg13g2_decap_4 FILLER_0_43_271 ();
 sg13g2_decap_8 FILLER_0_43_280 ();
 sg13g2_decap_8 FILLER_0_43_287 ();
 sg13g2_decap_8 FILLER_0_43_294 ();
 sg13g2_decap_8 FILLER_0_43_301 ();
 sg13g2_decap_8 FILLER_0_43_308 ();
 sg13g2_decap_8 FILLER_0_43_315 ();
 sg13g2_fill_1 FILLER_0_43_322 ();
 sg13g2_decap_8 FILLER_0_43_339 ();
 sg13g2_decap_8 FILLER_0_43_346 ();
 sg13g2_decap_4 FILLER_0_43_353 ();
 sg13g2_fill_1 FILLER_0_43_357 ();
 sg13g2_decap_8 FILLER_0_43_362 ();
 sg13g2_fill_2 FILLER_0_43_369 ();
 sg13g2_decap_4 FILLER_0_43_375 ();
 sg13g2_fill_2 FILLER_0_43_379 ();
 sg13g2_decap_4 FILLER_0_43_393 ();
 sg13g2_fill_1 FILLER_0_43_417 ();
 sg13g2_decap_4 FILLER_0_43_422 ();
 sg13g2_decap_8 FILLER_0_43_460 ();
 sg13g2_decap_8 FILLER_0_43_467 ();
 sg13g2_decap_8 FILLER_0_43_474 ();
 sg13g2_decap_8 FILLER_0_43_481 ();
 sg13g2_decap_4 FILLER_0_43_488 ();
 sg13g2_decap_4 FILLER_0_43_518 ();
 sg13g2_fill_1 FILLER_0_43_522 ();
 sg13g2_decap_8 FILLER_0_43_538 ();
 sg13g2_decap_8 FILLER_0_43_545 ();
 sg13g2_decap_4 FILLER_0_43_552 ();
 sg13g2_decap_4 FILLER_0_43_560 ();
 sg13g2_fill_1 FILLER_0_43_564 ();
 sg13g2_fill_2 FILLER_0_43_569 ();
 sg13g2_fill_2 FILLER_0_43_606 ();
 sg13g2_fill_1 FILLER_0_43_608 ();
 sg13g2_decap_4 FILLER_0_43_619 ();
 sg13g2_fill_1 FILLER_0_43_623 ();
 sg13g2_fill_2 FILLER_0_43_663 ();
 sg13g2_decap_8 FILLER_0_43_695 ();
 sg13g2_decap_8 FILLER_0_43_702 ();
 sg13g2_fill_1 FILLER_0_43_713 ();
 sg13g2_fill_1 FILLER_0_43_750 ();
 sg13g2_decap_4 FILLER_0_43_777 ();
 sg13g2_fill_2 FILLER_0_43_781 ();
 sg13g2_fill_2 FILLER_0_43_793 ();
 sg13g2_fill_1 FILLER_0_43_795 ();
 sg13g2_fill_1 FILLER_0_43_806 ();
 sg13g2_fill_2 FILLER_0_43_817 ();
 sg13g2_fill_1 FILLER_0_43_819 ();
 sg13g2_decap_8 FILLER_0_43_855 ();
 sg13g2_fill_2 FILLER_0_43_906 ();
 sg13g2_fill_2 FILLER_0_43_913 ();
 sg13g2_decap_8 FILLER_0_43_1006 ();
 sg13g2_fill_2 FILLER_0_43_1013 ();
 sg13g2_decap_8 FILLER_0_43_1019 ();
 sg13g2_fill_1 FILLER_0_43_1035 ();
 sg13g2_decap_4 FILLER_0_43_1040 ();
 sg13g2_fill_1 FILLER_0_43_1056 ();
 sg13g2_decap_8 FILLER_0_43_1062 ();
 sg13g2_decap_4 FILLER_0_43_1069 ();
 sg13g2_fill_1 FILLER_0_43_1073 ();
 sg13g2_decap_8 FILLER_0_43_1079 ();
 sg13g2_decap_8 FILLER_0_43_1086 ();
 sg13g2_decap_4 FILLER_0_43_1093 ();
 sg13g2_decap_8 FILLER_0_43_1118 ();
 sg13g2_decap_8 FILLER_0_43_1125 ();
 sg13g2_decap_8 FILLER_0_43_1132 ();
 sg13g2_decap_8 FILLER_0_43_1139 ();
 sg13g2_decap_8 FILLER_0_43_1146 ();
 sg13g2_decap_8 FILLER_0_43_1153 ();
 sg13g2_decap_8 FILLER_0_43_1160 ();
 sg13g2_decap_8 FILLER_0_43_1167 ();
 sg13g2_decap_8 FILLER_0_43_1174 ();
 sg13g2_decap_8 FILLER_0_43_1181 ();
 sg13g2_decap_8 FILLER_0_43_1188 ();
 sg13g2_decap_8 FILLER_0_43_1195 ();
 sg13g2_decap_8 FILLER_0_43_1202 ();
 sg13g2_decap_8 FILLER_0_43_1209 ();
 sg13g2_decap_8 FILLER_0_43_1216 ();
 sg13g2_decap_4 FILLER_0_43_1223 ();
 sg13g2_fill_1 FILLER_0_43_1227 ();
 sg13g2_decap_8 FILLER_0_44_0 ();
 sg13g2_decap_8 FILLER_0_44_7 ();
 sg13g2_decap_8 FILLER_0_44_14 ();
 sg13g2_decap_8 FILLER_0_44_21 ();
 sg13g2_decap_8 FILLER_0_44_28 ();
 sg13g2_decap_8 FILLER_0_44_35 ();
 sg13g2_decap_8 FILLER_0_44_42 ();
 sg13g2_decap_8 FILLER_0_44_49 ();
 sg13g2_decap_4 FILLER_0_44_56 ();
 sg13g2_fill_1 FILLER_0_44_60 ();
 sg13g2_decap_8 FILLER_0_44_65 ();
 sg13g2_decap_8 FILLER_0_44_98 ();
 sg13g2_fill_1 FILLER_0_44_105 ();
 sg13g2_fill_2 FILLER_0_44_110 ();
 sg13g2_decap_8 FILLER_0_44_127 ();
 sg13g2_decap_8 FILLER_0_44_134 ();
 sg13g2_decap_8 FILLER_0_44_141 ();
 sg13g2_decap_8 FILLER_0_44_148 ();
 sg13g2_decap_8 FILLER_0_44_155 ();
 sg13g2_decap_4 FILLER_0_44_162 ();
 sg13g2_fill_2 FILLER_0_44_166 ();
 sg13g2_fill_1 FILLER_0_44_178 ();
 sg13g2_decap_4 FILLER_0_44_183 ();
 sg13g2_fill_2 FILLER_0_44_187 ();
 sg13g2_decap_8 FILLER_0_44_193 ();
 sg13g2_decap_4 FILLER_0_44_215 ();
 sg13g2_fill_2 FILLER_0_44_249 ();
 sg13g2_fill_2 FILLER_0_44_266 ();
 sg13g2_decap_8 FILLER_0_44_314 ();
 sg13g2_decap_8 FILLER_0_44_321 ();
 sg13g2_decap_8 FILLER_0_44_328 ();
 sg13g2_decap_8 FILLER_0_44_335 ();
 sg13g2_decap_8 FILLER_0_44_342 ();
 sg13g2_decap_8 FILLER_0_44_349 ();
 sg13g2_fill_2 FILLER_0_44_356 ();
 sg13g2_fill_1 FILLER_0_44_358 ();
 sg13g2_decap_4 FILLER_0_44_421 ();
 sg13g2_fill_1 FILLER_0_44_438 ();
 sg13g2_decap_8 FILLER_0_44_465 ();
 sg13g2_decap_8 FILLER_0_44_472 ();
 sg13g2_fill_2 FILLER_0_44_479 ();
 sg13g2_fill_1 FILLER_0_44_481 ();
 sg13g2_decap_8 FILLER_0_44_507 ();
 sg13g2_decap_8 FILLER_0_44_514 ();
 sg13g2_fill_2 FILLER_0_44_521 ();
 sg13g2_fill_1 FILLER_0_44_523 ();
 sg13g2_decap_8 FILLER_0_44_555 ();
 sg13g2_decap_8 FILLER_0_44_562 ();
 sg13g2_decap_8 FILLER_0_44_569 ();
 sg13g2_fill_1 FILLER_0_44_576 ();
 sg13g2_decap_8 FILLER_0_44_693 ();
 sg13g2_decap_8 FILLER_0_44_700 ();
 sg13g2_decap_8 FILLER_0_44_707 ();
 sg13g2_decap_8 FILLER_0_44_714 ();
 sg13g2_fill_1 FILLER_0_44_721 ();
 sg13g2_fill_2 FILLER_0_44_771 ();
 sg13g2_fill_1 FILLER_0_44_773 ();
 sg13g2_fill_1 FILLER_0_44_805 ();
 sg13g2_fill_1 FILLER_0_44_837 ();
 sg13g2_decap_8 FILLER_0_44_864 ();
 sg13g2_decap_8 FILLER_0_44_871 ();
 sg13g2_fill_2 FILLER_0_44_948 ();
 sg13g2_fill_1 FILLER_0_44_950 ();
 sg13g2_decap_4 FILLER_0_44_963 ();
 sg13g2_fill_1 FILLER_0_44_967 ();
 sg13g2_decap_8 FILLER_0_44_972 ();
 sg13g2_fill_1 FILLER_0_44_979 ();
 sg13g2_decap_8 FILLER_0_44_990 ();
 sg13g2_decap_8 FILLER_0_44_997 ();
 sg13g2_decap_8 FILLER_0_44_1004 ();
 sg13g2_decap_8 FILLER_0_44_1011 ();
 sg13g2_decap_8 FILLER_0_44_1018 ();
 sg13g2_decap_8 FILLER_0_44_1025 ();
 sg13g2_decap_4 FILLER_0_44_1032 ();
 sg13g2_fill_1 FILLER_0_44_1036 ();
 sg13g2_fill_1 FILLER_0_44_1073 ();
 sg13g2_fill_2 FILLER_0_44_1079 ();
 sg13g2_decap_8 FILLER_0_44_1112 ();
 sg13g2_decap_8 FILLER_0_44_1119 ();
 sg13g2_decap_8 FILLER_0_44_1126 ();
 sg13g2_decap_8 FILLER_0_44_1133 ();
 sg13g2_decap_8 FILLER_0_44_1140 ();
 sg13g2_decap_8 FILLER_0_44_1147 ();
 sg13g2_decap_8 FILLER_0_44_1154 ();
 sg13g2_decap_8 FILLER_0_44_1161 ();
 sg13g2_decap_8 FILLER_0_44_1168 ();
 sg13g2_decap_8 FILLER_0_44_1175 ();
 sg13g2_decap_8 FILLER_0_44_1182 ();
 sg13g2_decap_8 FILLER_0_44_1189 ();
 sg13g2_decap_8 FILLER_0_44_1196 ();
 sg13g2_decap_8 FILLER_0_44_1203 ();
 sg13g2_decap_8 FILLER_0_44_1210 ();
 sg13g2_decap_8 FILLER_0_44_1217 ();
 sg13g2_decap_4 FILLER_0_44_1224 ();
 sg13g2_decap_8 FILLER_0_45_0 ();
 sg13g2_decap_8 FILLER_0_45_7 ();
 sg13g2_decap_8 FILLER_0_45_14 ();
 sg13g2_decap_8 FILLER_0_45_21 ();
 sg13g2_decap_8 FILLER_0_45_28 ();
 sg13g2_decap_8 FILLER_0_45_35 ();
 sg13g2_decap_8 FILLER_0_45_42 ();
 sg13g2_decap_8 FILLER_0_45_49 ();
 sg13g2_decap_8 FILLER_0_45_56 ();
 sg13g2_decap_8 FILLER_0_45_63 ();
 sg13g2_decap_4 FILLER_0_45_75 ();
 sg13g2_fill_2 FILLER_0_45_79 ();
 sg13g2_decap_8 FILLER_0_45_95 ();
 sg13g2_decap_8 FILLER_0_45_102 ();
 sg13g2_fill_2 FILLER_0_45_109 ();
 sg13g2_fill_1 FILLER_0_45_111 ();
 sg13g2_decap_4 FILLER_0_45_138 ();
 sg13g2_fill_1 FILLER_0_45_142 ();
 sg13g2_decap_8 FILLER_0_45_148 ();
 sg13g2_decap_8 FILLER_0_45_155 ();
 sg13g2_fill_1 FILLER_0_45_172 ();
 sg13g2_decap_8 FILLER_0_45_199 ();
 sg13g2_decap_8 FILLER_0_45_206 ();
 sg13g2_decap_8 FILLER_0_45_213 ();
 sg13g2_decap_8 FILLER_0_45_220 ();
 sg13g2_fill_2 FILLER_0_45_227 ();
 sg13g2_decap_8 FILLER_0_45_320 ();
 sg13g2_decap_8 FILLER_0_45_347 ();
 sg13g2_decap_8 FILLER_0_45_354 ();
 sg13g2_decap_4 FILLER_0_45_361 ();
 sg13g2_fill_2 FILLER_0_45_365 ();
 sg13g2_fill_2 FILLER_0_45_403 ();
 sg13g2_fill_2 FILLER_0_45_431 ();
 sg13g2_fill_2 FILLER_0_45_441 ();
 sg13g2_fill_2 FILLER_0_45_469 ();
 sg13g2_fill_2 FILLER_0_45_486 ();
 sg13g2_decap_4 FILLER_0_45_519 ();
 sg13g2_decap_4 FILLER_0_45_533 ();
 sg13g2_decap_4 FILLER_0_45_541 ();
 sg13g2_decap_8 FILLER_0_45_571 ();
 sg13g2_decap_8 FILLER_0_45_578 ();
 sg13g2_decap_4 FILLER_0_45_585 ();
 sg13g2_fill_1 FILLER_0_45_589 ();
 sg13g2_fill_1 FILLER_0_45_598 ();
 sg13g2_fill_2 FILLER_0_45_635 ();
 sg13g2_fill_1 FILLER_0_45_637 ();
 sg13g2_decap_8 FILLER_0_45_656 ();
 sg13g2_fill_2 FILLER_0_45_663 ();
 sg13g2_fill_1 FILLER_0_45_665 ();
 sg13g2_fill_2 FILLER_0_45_681 ();
 sg13g2_fill_1 FILLER_0_45_683 ();
 sg13g2_decap_8 FILLER_0_45_694 ();
 sg13g2_decap_8 FILLER_0_45_701 ();
 sg13g2_decap_8 FILLER_0_45_708 ();
 sg13g2_decap_8 FILLER_0_45_715 ();
 sg13g2_decap_8 FILLER_0_45_722 ();
 sg13g2_decap_8 FILLER_0_45_729 ();
 sg13g2_decap_8 FILLER_0_45_736 ();
 sg13g2_decap_8 FILLER_0_45_743 ();
 sg13g2_fill_2 FILLER_0_45_750 ();
 sg13g2_decap_8 FILLER_0_45_756 ();
 sg13g2_decap_8 FILLER_0_45_763 ();
 sg13g2_fill_2 FILLER_0_45_770 ();
 sg13g2_fill_2 FILLER_0_45_776 ();
 sg13g2_fill_1 FILLER_0_45_793 ();
 sg13g2_fill_1 FILLER_0_45_825 ();
 sg13g2_fill_2 FILLER_0_45_836 ();
 sg13g2_fill_1 FILLER_0_45_838 ();
 sg13g2_decap_8 FILLER_0_45_859 ();
 sg13g2_decap_8 FILLER_0_45_866 ();
 sg13g2_decap_8 FILLER_0_45_873 ();
 sg13g2_decap_8 FILLER_0_45_880 ();
 sg13g2_decap_8 FILLER_0_45_910 ();
 sg13g2_decap_8 FILLER_0_45_917 ();
 sg13g2_decap_4 FILLER_0_45_924 ();
 sg13g2_decap_8 FILLER_0_45_933 ();
 sg13g2_decap_8 FILLER_0_45_940 ();
 sg13g2_fill_1 FILLER_0_45_947 ();
 sg13g2_decap_8 FILLER_0_45_952 ();
 sg13g2_fill_2 FILLER_0_45_959 ();
 sg13g2_fill_1 FILLER_0_45_961 ();
 sg13g2_decap_8 FILLER_0_45_993 ();
 sg13g2_decap_8 FILLER_0_45_1000 ();
 sg13g2_decap_8 FILLER_0_45_1007 ();
 sg13g2_decap_4 FILLER_0_45_1018 ();
 sg13g2_fill_2 FILLER_0_45_1084 ();
 sg13g2_fill_2 FILLER_0_45_1096 ();
 sg13g2_decap_8 FILLER_0_45_1128 ();
 sg13g2_decap_8 FILLER_0_45_1135 ();
 sg13g2_decap_8 FILLER_0_45_1142 ();
 sg13g2_decap_8 FILLER_0_45_1149 ();
 sg13g2_decap_8 FILLER_0_45_1156 ();
 sg13g2_decap_8 FILLER_0_45_1163 ();
 sg13g2_decap_8 FILLER_0_45_1170 ();
 sg13g2_decap_8 FILLER_0_45_1177 ();
 sg13g2_decap_8 FILLER_0_45_1184 ();
 sg13g2_decap_8 FILLER_0_45_1191 ();
 sg13g2_decap_8 FILLER_0_45_1198 ();
 sg13g2_decap_8 FILLER_0_45_1205 ();
 sg13g2_decap_8 FILLER_0_45_1212 ();
 sg13g2_decap_8 FILLER_0_45_1219 ();
 sg13g2_fill_2 FILLER_0_45_1226 ();
 sg13g2_decap_8 FILLER_0_46_0 ();
 sg13g2_decap_8 FILLER_0_46_7 ();
 sg13g2_decap_8 FILLER_0_46_14 ();
 sg13g2_decap_8 FILLER_0_46_21 ();
 sg13g2_decap_8 FILLER_0_46_28 ();
 sg13g2_decap_4 FILLER_0_46_35 ();
 sg13g2_fill_1 FILLER_0_46_39 ();
 sg13g2_decap_4 FILLER_0_46_50 ();
 sg13g2_decap_8 FILLER_0_46_58 ();
 sg13g2_decap_4 FILLER_0_46_65 ();
 sg13g2_decap_8 FILLER_0_46_74 ();
 sg13g2_fill_1 FILLER_0_46_81 ();
 sg13g2_decap_8 FILLER_0_46_86 ();
 sg13g2_decap_8 FILLER_0_46_93 ();
 sg13g2_decap_4 FILLER_0_46_100 ();
 sg13g2_fill_1 FILLER_0_46_104 ();
 sg13g2_fill_2 FILLER_0_46_124 ();
 sg13g2_decap_8 FILLER_0_46_131 ();
 sg13g2_fill_1 FILLER_0_46_138 ();
 sg13g2_decap_4 FILLER_0_46_144 ();
 sg13g2_fill_2 FILLER_0_46_184 ();
 sg13g2_decap_8 FILLER_0_46_212 ();
 sg13g2_decap_8 FILLER_0_46_219 ();
 sg13g2_decap_8 FILLER_0_46_226 ();
 sg13g2_fill_2 FILLER_0_46_233 ();
 sg13g2_fill_1 FILLER_0_46_235 ();
 sg13g2_fill_1 FILLER_0_46_241 ();
 sg13g2_fill_1 FILLER_0_46_252 ();
 sg13g2_fill_1 FILLER_0_46_279 ();
 sg13g2_fill_1 FILLER_0_46_294 ();
 sg13g2_fill_2 FILLER_0_46_299 ();
 sg13g2_fill_1 FILLER_0_46_301 ();
 sg13g2_fill_2 FILLER_0_46_328 ();
 sg13g2_fill_1 FILLER_0_46_330 ();
 sg13g2_decap_4 FILLER_0_46_336 ();
 sg13g2_fill_2 FILLER_0_46_340 ();
 sg13g2_fill_1 FILLER_0_46_378 ();
 sg13g2_fill_2 FILLER_0_46_389 ();
 sg13g2_fill_1 FILLER_0_46_401 ();
 sg13g2_fill_2 FILLER_0_46_406 ();
 sg13g2_fill_2 FILLER_0_46_422 ();
 sg13g2_fill_1 FILLER_0_46_424 ();
 sg13g2_fill_2 FILLER_0_46_456 ();
 sg13g2_fill_1 FILLER_0_46_484 ();
 sg13g2_decap_4 FILLER_0_46_547 ();
 sg13g2_fill_2 FILLER_0_46_551 ();
 sg13g2_decap_8 FILLER_0_46_557 ();
 sg13g2_decap_8 FILLER_0_46_564 ();
 sg13g2_decap_8 FILLER_0_46_571 ();
 sg13g2_decap_8 FILLER_0_46_578 ();
 sg13g2_decap_8 FILLER_0_46_585 ();
 sg13g2_decap_8 FILLER_0_46_592 ();
 sg13g2_fill_2 FILLER_0_46_614 ();
 sg13g2_fill_1 FILLER_0_46_616 ();
 sg13g2_decap_8 FILLER_0_46_643 ();
 sg13g2_decap_8 FILLER_0_46_650 ();
 sg13g2_fill_2 FILLER_0_46_657 ();
 sg13g2_fill_1 FILLER_0_46_664 ();
 sg13g2_fill_1 FILLER_0_46_670 ();
 sg13g2_fill_1 FILLER_0_46_723 ();
 sg13g2_fill_2 FILLER_0_46_734 ();
 sg13g2_fill_1 FILLER_0_46_736 ();
 sg13g2_decap_4 FILLER_0_46_748 ();
 sg13g2_fill_2 FILLER_0_46_752 ();
 sg13g2_decap_8 FILLER_0_46_759 ();
 sg13g2_decap_8 FILLER_0_46_766 ();
 sg13g2_fill_1 FILLER_0_46_773 ();
 sg13g2_fill_1 FILLER_0_46_779 ();
 sg13g2_fill_2 FILLER_0_46_818 ();
 sg13g2_fill_2 FILLER_0_46_824 ();
 sg13g2_decap_8 FILLER_0_46_857 ();
 sg13g2_decap_8 FILLER_0_46_864 ();
 sg13g2_decap_8 FILLER_0_46_871 ();
 sg13g2_fill_2 FILLER_0_46_878 ();
 sg13g2_decap_8 FILLER_0_46_892 ();
 sg13g2_decap_8 FILLER_0_46_899 ();
 sg13g2_decap_4 FILLER_0_46_906 ();
 sg13g2_fill_1 FILLER_0_46_910 ();
 sg13g2_decap_4 FILLER_0_46_916 ();
 sg13g2_fill_1 FILLER_0_46_920 ();
 sg13g2_decap_8 FILLER_0_46_957 ();
 sg13g2_decap_4 FILLER_0_46_964 ();
 sg13g2_fill_2 FILLER_0_46_968 ();
 sg13g2_decap_4 FILLER_0_46_998 ();
 sg13g2_fill_2 FILLER_0_46_1002 ();
 sg13g2_fill_1 FILLER_0_46_1049 ();
 sg13g2_fill_1 FILLER_0_46_1060 ();
 sg13g2_fill_1 FILLER_0_46_1071 ();
 sg13g2_fill_1 FILLER_0_46_1098 ();
 sg13g2_decap_8 FILLER_0_46_1135 ();
 sg13g2_decap_8 FILLER_0_46_1142 ();
 sg13g2_decap_8 FILLER_0_46_1149 ();
 sg13g2_decap_8 FILLER_0_46_1156 ();
 sg13g2_decap_8 FILLER_0_46_1163 ();
 sg13g2_decap_8 FILLER_0_46_1170 ();
 sg13g2_decap_8 FILLER_0_46_1177 ();
 sg13g2_decap_8 FILLER_0_46_1184 ();
 sg13g2_decap_8 FILLER_0_46_1191 ();
 sg13g2_decap_8 FILLER_0_46_1198 ();
 sg13g2_decap_8 FILLER_0_46_1205 ();
 sg13g2_decap_8 FILLER_0_46_1212 ();
 sg13g2_decap_8 FILLER_0_46_1219 ();
 sg13g2_fill_2 FILLER_0_46_1226 ();
 sg13g2_decap_8 FILLER_0_47_0 ();
 sg13g2_decap_8 FILLER_0_47_7 ();
 sg13g2_decap_8 FILLER_0_47_14 ();
 sg13g2_decap_8 FILLER_0_47_21 ();
 sg13g2_decap_8 FILLER_0_47_28 ();
 sg13g2_fill_2 FILLER_0_47_61 ();
 sg13g2_fill_1 FILLER_0_47_63 ();
 sg13g2_decap_8 FILLER_0_47_90 ();
 sg13g2_fill_2 FILLER_0_47_123 ();
 sg13g2_fill_1 FILLER_0_47_143 ();
 sg13g2_decap_8 FILLER_0_47_204 ();
 sg13g2_decap_8 FILLER_0_47_211 ();
 sg13g2_decap_8 FILLER_0_47_218 ();
 sg13g2_decap_8 FILLER_0_47_225 ();
 sg13g2_decap_8 FILLER_0_47_232 ();
 sg13g2_decap_4 FILLER_0_47_239 ();
 sg13g2_fill_1 FILLER_0_47_243 ();
 sg13g2_decap_8 FILLER_0_47_248 ();
 sg13g2_decap_4 FILLER_0_47_255 ();
 sg13g2_decap_8 FILLER_0_47_263 ();
 sg13g2_fill_2 FILLER_0_47_270 ();
 sg13g2_decap_8 FILLER_0_47_276 ();
 sg13g2_decap_8 FILLER_0_47_283 ();
 sg13g2_decap_8 FILLER_0_47_290 ();
 sg13g2_fill_1 FILLER_0_47_297 ();
 sg13g2_fill_1 FILLER_0_47_313 ();
 sg13g2_fill_1 FILLER_0_47_340 ();
 sg13g2_decap_4 FILLER_0_47_377 ();
 sg13g2_fill_2 FILLER_0_47_381 ();
 sg13g2_decap_8 FILLER_0_47_387 ();
 sg13g2_fill_1 FILLER_0_47_394 ();
 sg13g2_decap_4 FILLER_0_47_398 ();
 sg13g2_fill_2 FILLER_0_47_402 ();
 sg13g2_decap_8 FILLER_0_47_412 ();
 sg13g2_decap_8 FILLER_0_47_419 ();
 sg13g2_decap_4 FILLER_0_47_426 ();
 sg13g2_fill_2 FILLER_0_47_438 ();
 sg13g2_fill_2 FILLER_0_47_458 ();
 sg13g2_fill_1 FILLER_0_47_460 ();
 sg13g2_fill_1 FILLER_0_47_471 ();
 sg13g2_fill_1 FILLER_0_47_498 ();
 sg13g2_fill_2 FILLER_0_47_503 ();
 sg13g2_fill_1 FILLER_0_47_530 ();
 sg13g2_decap_8 FILLER_0_47_535 ();
 sg13g2_decap_4 FILLER_0_47_542 ();
 sg13g2_fill_1 FILLER_0_47_546 ();
 sg13g2_decap_8 FILLER_0_47_555 ();
 sg13g2_decap_8 FILLER_0_47_562 ();
 sg13g2_decap_8 FILLER_0_47_569 ();
 sg13g2_decap_8 FILLER_0_47_576 ();
 sg13g2_decap_8 FILLER_0_47_583 ();
 sg13g2_decap_8 FILLER_0_47_590 ();
 sg13g2_decap_8 FILLER_0_47_597 ();
 sg13g2_decap_8 FILLER_0_47_608 ();
 sg13g2_fill_1 FILLER_0_47_615 ();
 sg13g2_fill_1 FILLER_0_47_621 ();
 sg13g2_decap_8 FILLER_0_47_636 ();
 sg13g2_decap_8 FILLER_0_47_643 ();
 sg13g2_fill_2 FILLER_0_47_650 ();
 sg13g2_fill_1 FILLER_0_47_710 ();
 sg13g2_fill_2 FILLER_0_47_737 ();
 sg13g2_decap_8 FILLER_0_47_795 ();
 sg13g2_decap_8 FILLER_0_47_802 ();
 sg13g2_fill_1 FILLER_0_47_809 ();
 sg13g2_decap_8 FILLER_0_47_817 ();
 sg13g2_decap_8 FILLER_0_47_824 ();
 sg13g2_fill_2 FILLER_0_47_831 ();
 sg13g2_fill_1 FILLER_0_47_833 ();
 sg13g2_decap_8 FILLER_0_47_838 ();
 sg13g2_fill_2 FILLER_0_47_845 ();
 sg13g2_fill_2 FILLER_0_47_917 ();
 sg13g2_fill_2 FILLER_0_47_949 ();
 sg13g2_fill_1 FILLER_0_47_964 ();
 sg13g2_fill_1 FILLER_0_47_996 ();
 sg13g2_fill_2 FILLER_0_47_1052 ();
 sg13g2_fill_2 FILLER_0_47_1058 ();
 sg13g2_fill_2 FILLER_0_47_1083 ();
 sg13g2_fill_1 FILLER_0_47_1085 ();
 sg13g2_fill_2 FILLER_0_47_1090 ();
 sg13g2_fill_1 FILLER_0_47_1110 ();
 sg13g2_fill_2 FILLER_0_47_1121 ();
 sg13g2_fill_1 FILLER_0_47_1123 ();
 sg13g2_decap_8 FILLER_0_47_1128 ();
 sg13g2_decap_8 FILLER_0_47_1135 ();
 sg13g2_decap_8 FILLER_0_47_1142 ();
 sg13g2_decap_8 FILLER_0_47_1149 ();
 sg13g2_decap_8 FILLER_0_47_1156 ();
 sg13g2_decap_8 FILLER_0_47_1163 ();
 sg13g2_decap_8 FILLER_0_47_1170 ();
 sg13g2_decap_8 FILLER_0_47_1177 ();
 sg13g2_decap_8 FILLER_0_47_1184 ();
 sg13g2_decap_8 FILLER_0_47_1191 ();
 sg13g2_decap_8 FILLER_0_47_1198 ();
 sg13g2_decap_8 FILLER_0_47_1205 ();
 sg13g2_decap_8 FILLER_0_47_1212 ();
 sg13g2_decap_8 FILLER_0_47_1219 ();
 sg13g2_fill_2 FILLER_0_47_1226 ();
 sg13g2_decap_8 FILLER_0_48_0 ();
 sg13g2_decap_8 FILLER_0_48_7 ();
 sg13g2_decap_8 FILLER_0_48_14 ();
 sg13g2_fill_2 FILLER_0_48_103 ();
 sg13g2_fill_1 FILLER_0_48_105 ();
 sg13g2_decap_8 FILLER_0_48_168 ();
 sg13g2_fill_2 FILLER_0_48_175 ();
 sg13g2_decap_8 FILLER_0_48_181 ();
 sg13g2_decap_8 FILLER_0_48_188 ();
 sg13g2_decap_8 FILLER_0_48_195 ();
 sg13g2_decap_8 FILLER_0_48_202 ();
 sg13g2_decap_8 FILLER_0_48_209 ();
 sg13g2_fill_2 FILLER_0_48_216 ();
 sg13g2_decap_8 FILLER_0_48_223 ();
 sg13g2_fill_1 FILLER_0_48_230 ();
 sg13g2_decap_8 FILLER_0_48_246 ();
 sg13g2_decap_4 FILLER_0_48_253 ();
 sg13g2_fill_2 FILLER_0_48_265 ();
 sg13g2_fill_1 FILLER_0_48_267 ();
 sg13g2_decap_4 FILLER_0_48_273 ();
 sg13g2_fill_1 FILLER_0_48_277 ();
 sg13g2_decap_8 FILLER_0_48_283 ();
 sg13g2_decap_8 FILLER_0_48_290 ();
 sg13g2_fill_1 FILLER_0_48_297 ();
 sg13g2_decap_4 FILLER_0_48_357 ();
 sg13g2_decap_8 FILLER_0_48_365 ();
 sg13g2_decap_4 FILLER_0_48_372 ();
 sg13g2_decap_8 FILLER_0_48_410 ();
 sg13g2_decap_8 FILLER_0_48_417 ();
 sg13g2_decap_8 FILLER_0_48_428 ();
 sg13g2_decap_4 FILLER_0_48_435 ();
 sg13g2_decap_8 FILLER_0_48_452 ();
 sg13g2_fill_2 FILLER_0_48_459 ();
 sg13g2_fill_2 FILLER_0_48_466 ();
 sg13g2_fill_1 FILLER_0_48_468 ();
 sg13g2_decap_4 FILLER_0_48_473 ();
 sg13g2_fill_2 FILLER_0_48_477 ();
 sg13g2_decap_8 FILLER_0_48_483 ();
 sg13g2_decap_8 FILLER_0_48_490 ();
 sg13g2_decap_8 FILLER_0_48_501 ();
 sg13g2_decap_8 FILLER_0_48_508 ();
 sg13g2_decap_8 FILLER_0_48_515 ();
 sg13g2_decap_8 FILLER_0_48_522 ();
 sg13g2_decap_8 FILLER_0_48_529 ();
 sg13g2_decap_4 FILLER_0_48_536 ();
 sg13g2_fill_2 FILLER_0_48_540 ();
 sg13g2_fill_1 FILLER_0_48_582 ();
 sg13g2_decap_8 FILLER_0_48_588 ();
 sg13g2_decap_8 FILLER_0_48_605 ();
 sg13g2_decap_8 FILLER_0_48_612 ();
 sg13g2_fill_2 FILLER_0_48_619 ();
 sg13g2_fill_1 FILLER_0_48_621 ();
 sg13g2_fill_2 FILLER_0_48_631 ();
 sg13g2_fill_1 FILLER_0_48_633 ();
 sg13g2_decap_8 FILLER_0_48_691 ();
 sg13g2_fill_2 FILLER_0_48_698 ();
 sg13g2_fill_2 FILLER_0_48_704 ();
 sg13g2_fill_1 FILLER_0_48_750 ();
 sg13g2_decap_8 FILLER_0_48_785 ();
 sg13g2_decap_8 FILLER_0_48_792 ();
 sg13g2_decap_8 FILLER_0_48_799 ();
 sg13g2_decap_8 FILLER_0_48_806 ();
 sg13g2_decap_8 FILLER_0_48_813 ();
 sg13g2_decap_8 FILLER_0_48_820 ();
 sg13g2_decap_8 FILLER_0_48_827 ();
 sg13g2_decap_4 FILLER_0_48_834 ();
 sg13g2_fill_2 FILLER_0_48_838 ();
 sg13g2_fill_2 FILLER_0_48_990 ();
 sg13g2_decap_8 FILLER_0_48_1033 ();
 sg13g2_decap_8 FILLER_0_48_1040 ();
 sg13g2_decap_8 FILLER_0_48_1047 ();
 sg13g2_decap_8 FILLER_0_48_1054 ();
 sg13g2_decap_8 FILLER_0_48_1061 ();
 sg13g2_decap_8 FILLER_0_48_1068 ();
 sg13g2_fill_2 FILLER_0_48_1075 ();
 sg13g2_decap_8 FILLER_0_48_1082 ();
 sg13g2_decap_8 FILLER_0_48_1089 ();
 sg13g2_decap_4 FILLER_0_48_1096 ();
 sg13g2_decap_8 FILLER_0_48_1104 ();
 sg13g2_fill_1 FILLER_0_48_1111 ();
 sg13g2_decap_8 FILLER_0_48_1143 ();
 sg13g2_decap_8 FILLER_0_48_1150 ();
 sg13g2_decap_8 FILLER_0_48_1157 ();
 sg13g2_decap_8 FILLER_0_48_1164 ();
 sg13g2_decap_8 FILLER_0_48_1171 ();
 sg13g2_decap_8 FILLER_0_48_1178 ();
 sg13g2_decap_8 FILLER_0_48_1185 ();
 sg13g2_decap_8 FILLER_0_48_1192 ();
 sg13g2_decap_8 FILLER_0_48_1199 ();
 sg13g2_decap_8 FILLER_0_48_1206 ();
 sg13g2_decap_8 FILLER_0_48_1213 ();
 sg13g2_decap_8 FILLER_0_48_1220 ();
 sg13g2_fill_1 FILLER_0_48_1227 ();
 sg13g2_decap_8 FILLER_0_49_0 ();
 sg13g2_decap_8 FILLER_0_49_7 ();
 sg13g2_decap_8 FILLER_0_49_14 ();
 sg13g2_decap_8 FILLER_0_49_21 ();
 sg13g2_fill_1 FILLER_0_49_28 ();
 sg13g2_decap_4 FILLER_0_49_33 ();
 sg13g2_fill_2 FILLER_0_49_37 ();
 sg13g2_fill_2 FILLER_0_49_63 ();
 sg13g2_fill_1 FILLER_0_49_65 ();
 sg13g2_decap_4 FILLER_0_49_76 ();
 sg13g2_fill_1 FILLER_0_49_80 ();
 sg13g2_decap_8 FILLER_0_49_96 ();
 sg13g2_decap_8 FILLER_0_49_156 ();
 sg13g2_decap_8 FILLER_0_49_163 ();
 sg13g2_decap_4 FILLER_0_49_170 ();
 sg13g2_decap_8 FILLER_0_49_186 ();
 sg13g2_decap_8 FILLER_0_49_193 ();
 sg13g2_decap_8 FILLER_0_49_200 ();
 sg13g2_fill_1 FILLER_0_49_207 ();
 sg13g2_decap_8 FILLER_0_49_218 ();
 sg13g2_decap_4 FILLER_0_49_225 ();
 sg13g2_fill_1 FILLER_0_49_229 ();
 sg13g2_decap_4 FILLER_0_49_302 ();
 sg13g2_fill_1 FILLER_0_49_306 ();
 sg13g2_decap_8 FILLER_0_49_312 ();
 sg13g2_fill_2 FILLER_0_49_319 ();
 sg13g2_decap_8 FILLER_0_49_337 ();
 sg13g2_decap_8 FILLER_0_49_344 ();
 sg13g2_decap_8 FILLER_0_49_351 ();
 sg13g2_decap_8 FILLER_0_49_358 ();
 sg13g2_decap_8 FILLER_0_49_365 ();
 sg13g2_fill_2 FILLER_0_49_372 ();
 sg13g2_fill_1 FILLER_0_49_374 ();
 sg13g2_fill_2 FILLER_0_49_406 ();
 sg13g2_fill_1 FILLER_0_49_408 ();
 sg13g2_fill_2 FILLER_0_49_414 ();
 sg13g2_fill_1 FILLER_0_49_416 ();
 sg13g2_decap_8 FILLER_0_49_475 ();
 sg13g2_decap_8 FILLER_0_49_482 ();
 sg13g2_decap_8 FILLER_0_49_489 ();
 sg13g2_decap_8 FILLER_0_49_496 ();
 sg13g2_fill_2 FILLER_0_49_531 ();
 sg13g2_fill_1 FILLER_0_49_543 ();
 sg13g2_fill_1 FILLER_0_49_620 ();
 sg13g2_decap_8 FILLER_0_49_626 ();
 sg13g2_decap_8 FILLER_0_49_633 ();
 sg13g2_decap_8 FILLER_0_49_640 ();
 sg13g2_decap_4 FILLER_0_49_647 ();
 sg13g2_fill_2 FILLER_0_49_651 ();
 sg13g2_decap_8 FILLER_0_49_679 ();
 sg13g2_fill_2 FILLER_0_49_686 ();
 sg13g2_fill_1 FILLER_0_49_728 ();
 sg13g2_decap_8 FILLER_0_49_770 ();
 sg13g2_decap_8 FILLER_0_49_777 ();
 sg13g2_decap_8 FILLER_0_49_784 ();
 sg13g2_decap_8 FILLER_0_49_791 ();
 sg13g2_decap_4 FILLER_0_49_798 ();
 sg13g2_decap_8 FILLER_0_49_837 ();
 sg13g2_decap_4 FILLER_0_49_844 ();
 sg13g2_fill_2 FILLER_0_49_901 ();
 sg13g2_fill_1 FILLER_0_49_903 ();
 sg13g2_fill_2 FILLER_0_49_918 ();
 sg13g2_fill_1 FILLER_0_49_930 ();
 sg13g2_decap_8 FILLER_0_49_950 ();
 sg13g2_decap_4 FILLER_0_49_957 ();
 sg13g2_decap_4 FILLER_0_49_966 ();
 sg13g2_fill_1 FILLER_0_49_970 ();
 sg13g2_decap_8 FILLER_0_49_985 ();
 sg13g2_decap_4 FILLER_0_49_992 ();
 sg13g2_fill_2 FILLER_0_49_996 ();
 sg13g2_decap_8 FILLER_0_49_1039 ();
 sg13g2_decap_8 FILLER_0_49_1064 ();
 sg13g2_decap_8 FILLER_0_49_1071 ();
 sg13g2_decap_8 FILLER_0_49_1078 ();
 sg13g2_decap_8 FILLER_0_49_1085 ();
 sg13g2_decap_4 FILLER_0_49_1092 ();
 sg13g2_fill_2 FILLER_0_49_1096 ();
 sg13g2_decap_8 FILLER_0_49_1123 ();
 sg13g2_decap_8 FILLER_0_49_1130 ();
 sg13g2_decap_8 FILLER_0_49_1137 ();
 sg13g2_decap_8 FILLER_0_49_1144 ();
 sg13g2_decap_8 FILLER_0_49_1151 ();
 sg13g2_decap_8 FILLER_0_49_1158 ();
 sg13g2_decap_8 FILLER_0_49_1165 ();
 sg13g2_decap_8 FILLER_0_49_1172 ();
 sg13g2_decap_8 FILLER_0_49_1179 ();
 sg13g2_decap_8 FILLER_0_49_1186 ();
 sg13g2_decap_8 FILLER_0_49_1193 ();
 sg13g2_decap_8 FILLER_0_49_1200 ();
 sg13g2_decap_8 FILLER_0_49_1207 ();
 sg13g2_decap_8 FILLER_0_49_1214 ();
 sg13g2_decap_8 FILLER_0_49_1221 ();
 sg13g2_decap_8 FILLER_0_50_0 ();
 sg13g2_decap_8 FILLER_0_50_7 ();
 sg13g2_decap_8 FILLER_0_50_14 ();
 sg13g2_decap_8 FILLER_0_50_21 ();
 sg13g2_decap_4 FILLER_0_50_28 ();
 sg13g2_fill_1 FILLER_0_50_32 ();
 sg13g2_decap_4 FILLER_0_50_38 ();
 sg13g2_fill_1 FILLER_0_50_42 ();
 sg13g2_decap_4 FILLER_0_50_65 ();
 sg13g2_fill_2 FILLER_0_50_69 ();
 sg13g2_decap_8 FILLER_0_50_75 ();
 sg13g2_decap_8 FILLER_0_50_82 ();
 sg13g2_decap_8 FILLER_0_50_89 ();
 sg13g2_decap_4 FILLER_0_50_96 ();
 sg13g2_decap_8 FILLER_0_50_104 ();
 sg13g2_decap_8 FILLER_0_50_111 ();
 sg13g2_decap_8 FILLER_0_50_118 ();
 sg13g2_fill_2 FILLER_0_50_125 ();
 sg13g2_fill_1 FILLER_0_50_127 ();
 sg13g2_decap_8 FILLER_0_50_135 ();
 sg13g2_decap_8 FILLER_0_50_142 ();
 sg13g2_decap_8 FILLER_0_50_149 ();
 sg13g2_decap_4 FILLER_0_50_156 ();
 sg13g2_fill_1 FILLER_0_50_160 ();
 sg13g2_decap_8 FILLER_0_50_169 ();
 sg13g2_decap_8 FILLER_0_50_176 ();
 sg13g2_decap_4 FILLER_0_50_183 ();
 sg13g2_fill_1 FILLER_0_50_218 ();
 sg13g2_fill_2 FILLER_0_50_254 ();
 sg13g2_decap_8 FILLER_0_50_334 ();
 sg13g2_decap_8 FILLER_0_50_341 ();
 sg13g2_decap_8 FILLER_0_50_348 ();
 sg13g2_decap_8 FILLER_0_50_359 ();
 sg13g2_fill_1 FILLER_0_50_366 ();
 sg13g2_decap_8 FILLER_0_50_372 ();
 sg13g2_decap_8 FILLER_0_50_485 ();
 sg13g2_decap_8 FILLER_0_50_492 ();
 sg13g2_decap_4 FILLER_0_50_499 ();
 sg13g2_fill_1 FILLER_0_50_503 ();
 sg13g2_fill_2 FILLER_0_50_565 ();
 sg13g2_fill_1 FILLER_0_50_567 ();
 sg13g2_decap_8 FILLER_0_50_640 ();
 sg13g2_decap_8 FILLER_0_50_647 ();
 sg13g2_fill_2 FILLER_0_50_654 ();
 sg13g2_fill_1 FILLER_0_50_656 ();
 sg13g2_fill_2 FILLER_0_50_669 ();
 sg13g2_fill_1 FILLER_0_50_671 ();
 sg13g2_decap_4 FILLER_0_50_682 ();
 sg13g2_fill_2 FILLER_0_50_686 ();
 sg13g2_fill_2 FILLER_0_50_692 ();
 sg13g2_fill_1 FILLER_0_50_694 ();
 sg13g2_decap_4 FILLER_0_50_725 ();
 sg13g2_fill_1 FILLER_0_50_729 ();
 sg13g2_decap_4 FILLER_0_50_734 ();
 sg13g2_fill_2 FILLER_0_50_743 ();
 sg13g2_fill_1 FILLER_0_50_745 ();
 sg13g2_decap_8 FILLER_0_50_750 ();
 sg13g2_decap_8 FILLER_0_50_762 ();
 sg13g2_decap_4 FILLER_0_50_769 ();
 sg13g2_fill_2 FILLER_0_50_773 ();
 sg13g2_fill_1 FILLER_0_50_785 ();
 sg13g2_fill_2 FILLER_0_50_817 ();
 sg13g2_fill_1 FILLER_0_50_819 ();
 sg13g2_fill_2 FILLER_0_50_830 ();
 sg13g2_fill_1 FILLER_0_50_832 ();
 sg13g2_decap_8 FILLER_0_50_851 ();
 sg13g2_decap_8 FILLER_0_50_858 ();
 sg13g2_decap_8 FILLER_0_50_865 ();
 sg13g2_fill_2 FILLER_0_50_872 ();
 sg13g2_fill_1 FILLER_0_50_874 ();
 sg13g2_decap_8 FILLER_0_50_880 ();
 sg13g2_decap_8 FILLER_0_50_887 ();
 sg13g2_decap_4 FILLER_0_50_894 ();
 sg13g2_fill_1 FILLER_0_50_898 ();
 sg13g2_decap_8 FILLER_0_50_903 ();
 sg13g2_decap_8 FILLER_0_50_910 ();
 sg13g2_decap_8 FILLER_0_50_917 ();
 sg13g2_decap_4 FILLER_0_50_924 ();
 sg13g2_fill_2 FILLER_0_50_928 ();
 sg13g2_decap_8 FILLER_0_50_935 ();
 sg13g2_decap_8 FILLER_0_50_942 ();
 sg13g2_decap_8 FILLER_0_50_949 ();
 sg13g2_fill_2 FILLER_0_50_956 ();
 sg13g2_fill_1 FILLER_0_50_958 ();
 sg13g2_decap_8 FILLER_0_50_989 ();
 sg13g2_decap_8 FILLER_0_50_996 ();
 sg13g2_decap_4 FILLER_0_50_1003 ();
 sg13g2_fill_1 FILLER_0_50_1007 ();
 sg13g2_decap_8 FILLER_0_50_1069 ();
 sg13g2_fill_1 FILLER_0_50_1076 ();
 sg13g2_decap_8 FILLER_0_50_1081 ();
 sg13g2_decap_8 FILLER_0_50_1088 ();
 sg13g2_decap_8 FILLER_0_50_1129 ();
 sg13g2_decap_8 FILLER_0_50_1136 ();
 sg13g2_decap_8 FILLER_0_50_1143 ();
 sg13g2_decap_8 FILLER_0_50_1150 ();
 sg13g2_decap_8 FILLER_0_50_1157 ();
 sg13g2_decap_8 FILLER_0_50_1164 ();
 sg13g2_decap_8 FILLER_0_50_1171 ();
 sg13g2_decap_8 FILLER_0_50_1178 ();
 sg13g2_decap_8 FILLER_0_50_1185 ();
 sg13g2_decap_8 FILLER_0_50_1192 ();
 sg13g2_decap_8 FILLER_0_50_1199 ();
 sg13g2_decap_8 FILLER_0_50_1206 ();
 sg13g2_decap_8 FILLER_0_50_1213 ();
 sg13g2_decap_8 FILLER_0_50_1220 ();
 sg13g2_fill_1 FILLER_0_50_1227 ();
 sg13g2_decap_8 FILLER_0_51_0 ();
 sg13g2_decap_8 FILLER_0_51_7 ();
 sg13g2_decap_8 FILLER_0_51_14 ();
 sg13g2_fill_1 FILLER_0_51_21 ();
 sg13g2_fill_1 FILLER_0_51_58 ();
 sg13g2_decap_4 FILLER_0_51_74 ();
 sg13g2_decap_4 FILLER_0_51_96 ();
 sg13g2_fill_1 FILLER_0_51_100 ();
 sg13g2_fill_2 FILLER_0_51_106 ();
 sg13g2_decap_4 FILLER_0_51_116 ();
 sg13g2_fill_2 FILLER_0_51_120 ();
 sg13g2_decap_8 FILLER_0_51_148 ();
 sg13g2_decap_8 FILLER_0_51_155 ();
 sg13g2_decap_8 FILLER_0_51_162 ();
 sg13g2_fill_2 FILLER_0_51_169 ();
 sg13g2_fill_1 FILLER_0_51_171 ();
 sg13g2_decap_4 FILLER_0_51_176 ();
 sg13g2_fill_2 FILLER_0_51_180 ();
 sg13g2_decap_8 FILLER_0_51_191 ();
 sg13g2_fill_1 FILLER_0_51_262 ();
 sg13g2_fill_1 FILLER_0_51_297 ();
 sg13g2_fill_1 FILLER_0_51_308 ();
 sg13g2_fill_1 FILLER_0_51_319 ();
 sg13g2_fill_2 FILLER_0_51_346 ();
 sg13g2_decap_8 FILLER_0_51_374 ();
 sg13g2_decap_8 FILLER_0_51_381 ();
 sg13g2_fill_1 FILLER_0_51_392 ();
 sg13g2_fill_2 FILLER_0_51_403 ();
 sg13g2_fill_2 FILLER_0_51_409 ();
 sg13g2_decap_4 FILLER_0_51_435 ();
 sg13g2_decap_4 FILLER_0_51_491 ();
 sg13g2_fill_2 FILLER_0_51_495 ();
 sg13g2_fill_1 FILLER_0_51_559 ();
 sg13g2_decap_8 FILLER_0_51_564 ();
 sg13g2_decap_8 FILLER_0_51_571 ();
 sg13g2_decap_4 FILLER_0_51_578 ();
 sg13g2_fill_2 FILLER_0_51_582 ();
 sg13g2_fill_1 FILLER_0_51_588 ();
 sg13g2_fill_1 FILLER_0_51_593 ();
 sg13g2_fill_1 FILLER_0_51_598 ();
 sg13g2_fill_1 FILLER_0_51_604 ();
 sg13g2_fill_1 FILLER_0_51_615 ();
 sg13g2_decap_8 FILLER_0_51_642 ();
 sg13g2_decap_8 FILLER_0_51_649 ();
 sg13g2_fill_2 FILLER_0_51_656 ();
 sg13g2_fill_1 FILLER_0_51_663 ();
 sg13g2_fill_1 FILLER_0_51_690 ();
 sg13g2_fill_2 FILLER_0_51_696 ();
 sg13g2_fill_1 FILLER_0_51_708 ();
 sg13g2_decap_8 FILLER_0_51_719 ();
 sg13g2_decap_8 FILLER_0_51_726 ();
 sg13g2_decap_8 FILLER_0_51_733 ();
 sg13g2_decap_8 FILLER_0_51_740 ();
 sg13g2_decap_8 FILLER_0_51_747 ();
 sg13g2_fill_2 FILLER_0_51_754 ();
 sg13g2_decap_8 FILLER_0_51_786 ();
 sg13g2_fill_1 FILLER_0_51_811 ();
 sg13g2_fill_1 FILLER_0_51_822 ();
 sg13g2_fill_1 FILLER_0_51_867 ();
 sg13g2_decap_8 FILLER_0_51_899 ();
 sg13g2_decap_8 FILLER_0_51_906 ();
 sg13g2_decap_8 FILLER_0_51_913 ();
 sg13g2_decap_8 FILLER_0_51_920 ();
 sg13g2_decap_8 FILLER_0_51_927 ();
 sg13g2_decap_8 FILLER_0_51_934 ();
 sg13g2_decap_8 FILLER_0_51_941 ();
 sg13g2_decap_8 FILLER_0_51_948 ();
 sg13g2_decap_8 FILLER_0_51_955 ();
 sg13g2_decap_8 FILLER_0_51_962 ();
 sg13g2_fill_2 FILLER_0_51_979 ();
 sg13g2_fill_1 FILLER_0_51_981 ();
 sg13g2_decap_8 FILLER_0_51_986 ();
 sg13g2_decap_8 FILLER_0_51_993 ();
 sg13g2_decap_8 FILLER_0_51_1000 ();
 sg13g2_decap_8 FILLER_0_51_1007 ();
 sg13g2_fill_2 FILLER_0_51_1014 ();
 sg13g2_decap_8 FILLER_0_51_1025 ();
 sg13g2_decap_4 FILLER_0_51_1032 ();
 sg13g2_decap_4 FILLER_0_51_1050 ();
 sg13g2_fill_1 FILLER_0_51_1054 ();
 sg13g2_fill_2 FILLER_0_51_1085 ();
 sg13g2_fill_1 FILLER_0_51_1087 ();
 sg13g2_decap_8 FILLER_0_51_1119 ();
 sg13g2_decap_8 FILLER_0_51_1126 ();
 sg13g2_decap_8 FILLER_0_51_1133 ();
 sg13g2_decap_8 FILLER_0_51_1140 ();
 sg13g2_decap_8 FILLER_0_51_1147 ();
 sg13g2_decap_8 FILLER_0_51_1154 ();
 sg13g2_decap_8 FILLER_0_51_1161 ();
 sg13g2_decap_8 FILLER_0_51_1168 ();
 sg13g2_decap_8 FILLER_0_51_1175 ();
 sg13g2_decap_8 FILLER_0_51_1182 ();
 sg13g2_decap_8 FILLER_0_51_1189 ();
 sg13g2_decap_8 FILLER_0_51_1196 ();
 sg13g2_decap_8 FILLER_0_51_1203 ();
 sg13g2_decap_8 FILLER_0_51_1210 ();
 sg13g2_decap_8 FILLER_0_51_1217 ();
 sg13g2_decap_4 FILLER_0_51_1224 ();
 sg13g2_decap_8 FILLER_0_52_0 ();
 sg13g2_decap_8 FILLER_0_52_7 ();
 sg13g2_decap_8 FILLER_0_52_14 ();
 sg13g2_decap_4 FILLER_0_52_21 ();
 sg13g2_decap_4 FILLER_0_52_34 ();
 sg13g2_fill_1 FILLER_0_52_82 ();
 sg13g2_decap_8 FILLER_0_52_138 ();
 sg13g2_decap_8 FILLER_0_52_145 ();
 sg13g2_fill_2 FILLER_0_52_152 ();
 sg13g2_fill_1 FILLER_0_52_154 ();
 sg13g2_decap_8 FILLER_0_52_164 ();
 sg13g2_decap_8 FILLER_0_52_171 ();
 sg13g2_fill_2 FILLER_0_52_178 ();
 sg13g2_decap_8 FILLER_0_52_216 ();
 sg13g2_decap_8 FILLER_0_52_223 ();
 sg13g2_decap_8 FILLER_0_52_230 ();
 sg13g2_decap_8 FILLER_0_52_237 ();
 sg13g2_fill_2 FILLER_0_52_244 ();
 sg13g2_decap_8 FILLER_0_52_250 ();
 sg13g2_decap_8 FILLER_0_52_257 ();
 sg13g2_decap_8 FILLER_0_52_264 ();
 sg13g2_decap_4 FILLER_0_52_271 ();
 sg13g2_fill_1 FILLER_0_52_279 ();
 sg13g2_decap_4 FILLER_0_52_294 ();
 sg13g2_fill_2 FILLER_0_52_298 ();
 sg13g2_fill_1 FILLER_0_52_305 ();
 sg13g2_fill_1 FILLER_0_52_315 ();
 sg13g2_fill_1 FILLER_0_52_324 ();
 sg13g2_fill_1 FILLER_0_52_390 ();
 sg13g2_decap_8 FILLER_0_52_406 ();
 sg13g2_decap_8 FILLER_0_52_418 ();
 sg13g2_decap_8 FILLER_0_52_425 ();
 sg13g2_decap_8 FILLER_0_52_432 ();
 sg13g2_decap_8 FILLER_0_52_439 ();
 sg13g2_decap_4 FILLER_0_52_446 ();
 sg13g2_fill_2 FILLER_0_52_450 ();
 sg13g2_fill_2 FILLER_0_52_472 ();
 sg13g2_decap_8 FILLER_0_52_478 ();
 sg13g2_decap_8 FILLER_0_52_485 ();
 sg13g2_decap_4 FILLER_0_52_492 ();
 sg13g2_fill_1 FILLER_0_52_525 ();
 sg13g2_decap_8 FILLER_0_52_537 ();
 sg13g2_decap_8 FILLER_0_52_544 ();
 sg13g2_decap_8 FILLER_0_52_551 ();
 sg13g2_decap_4 FILLER_0_52_563 ();
 sg13g2_fill_1 FILLER_0_52_567 ();
 sg13g2_decap_8 FILLER_0_52_572 ();
 sg13g2_decap_8 FILLER_0_52_583 ();
 sg13g2_decap_8 FILLER_0_52_590 ();
 sg13g2_decap_4 FILLER_0_52_597 ();
 sg13g2_fill_2 FILLER_0_52_601 ();
 sg13g2_decap_8 FILLER_0_52_629 ();
 sg13g2_fill_1 FILLER_0_52_636 ();
 sg13g2_decap_4 FILLER_0_52_647 ();
 sg13g2_fill_2 FILLER_0_52_651 ();
 sg13g2_decap_8 FILLER_0_52_714 ();
 sg13g2_decap_8 FILLER_0_52_721 ();
 sg13g2_decap_8 FILLER_0_52_728 ();
 sg13g2_decap_8 FILLER_0_52_735 ();
 sg13g2_decap_8 FILLER_0_52_753 ();
 sg13g2_fill_1 FILLER_0_52_760 ();
 sg13g2_fill_1 FILLER_0_52_771 ();
 sg13g2_fill_1 FILLER_0_52_798 ();
 sg13g2_fill_1 FILLER_0_52_825 ();
 sg13g2_fill_1 FILLER_0_52_831 ();
 sg13g2_decap_8 FILLER_0_52_915 ();
 sg13g2_decap_8 FILLER_0_52_922 ();
 sg13g2_decap_8 FILLER_0_52_929 ();
 sg13g2_decap_8 FILLER_0_52_936 ();
 sg13g2_decap_8 FILLER_0_52_943 ();
 sg13g2_decap_8 FILLER_0_52_950 ();
 sg13g2_decap_8 FILLER_0_52_957 ();
 sg13g2_decap_4 FILLER_0_52_964 ();
 sg13g2_fill_2 FILLER_0_52_968 ();
 sg13g2_decap_4 FILLER_0_52_1001 ();
 sg13g2_decap_8 FILLER_0_52_1009 ();
 sg13g2_fill_2 FILLER_0_52_1016 ();
 sg13g2_decap_8 FILLER_0_52_1064 ();
 sg13g2_decap_8 FILLER_0_52_1071 ();
 sg13g2_decap_4 FILLER_0_52_1078 ();
 sg13g2_fill_1 FILLER_0_52_1082 ();
 sg13g2_decap_8 FILLER_0_52_1124 ();
 sg13g2_decap_8 FILLER_0_52_1131 ();
 sg13g2_decap_8 FILLER_0_52_1138 ();
 sg13g2_decap_8 FILLER_0_52_1145 ();
 sg13g2_decap_8 FILLER_0_52_1152 ();
 sg13g2_decap_8 FILLER_0_52_1159 ();
 sg13g2_decap_8 FILLER_0_52_1166 ();
 sg13g2_decap_8 FILLER_0_52_1173 ();
 sg13g2_decap_8 FILLER_0_52_1180 ();
 sg13g2_decap_8 FILLER_0_52_1187 ();
 sg13g2_decap_8 FILLER_0_52_1194 ();
 sg13g2_decap_8 FILLER_0_52_1201 ();
 sg13g2_decap_8 FILLER_0_52_1208 ();
 sg13g2_decap_8 FILLER_0_52_1215 ();
 sg13g2_decap_4 FILLER_0_52_1222 ();
 sg13g2_fill_2 FILLER_0_52_1226 ();
 sg13g2_decap_8 FILLER_0_53_0 ();
 sg13g2_decap_8 FILLER_0_53_7 ();
 sg13g2_decap_8 FILLER_0_53_14 ();
 sg13g2_decap_8 FILLER_0_53_21 ();
 sg13g2_decap_8 FILLER_0_53_28 ();
 sg13g2_decap_8 FILLER_0_53_35 ();
 sg13g2_decap_4 FILLER_0_53_42 ();
 sg13g2_fill_2 FILLER_0_53_76 ();
 sg13g2_fill_2 FILLER_0_53_114 ();
 sg13g2_decap_8 FILLER_0_53_178 ();
 sg13g2_decap_8 FILLER_0_53_185 ();
 sg13g2_decap_4 FILLER_0_53_192 ();
 sg13g2_fill_1 FILLER_0_53_196 ();
 sg13g2_fill_1 FILLER_0_53_202 ();
 sg13g2_decap_8 FILLER_0_53_229 ();
 sg13g2_decap_8 FILLER_0_53_236 ();
 sg13g2_decap_8 FILLER_0_53_243 ();
 sg13g2_decap_8 FILLER_0_53_250 ();
 sg13g2_decap_8 FILLER_0_53_257 ();
 sg13g2_decap_8 FILLER_0_53_264 ();
 sg13g2_decap_8 FILLER_0_53_271 ();
 sg13g2_decap_8 FILLER_0_53_278 ();
 sg13g2_decap_8 FILLER_0_53_285 ();
 sg13g2_decap_4 FILLER_0_53_292 ();
 sg13g2_fill_1 FILLER_0_53_296 ();
 sg13g2_decap_8 FILLER_0_53_305 ();
 sg13g2_fill_1 FILLER_0_53_312 ();
 sg13g2_fill_2 FILLER_0_53_317 ();
 sg13g2_fill_1 FILLER_0_53_354 ();
 sg13g2_decap_8 FILLER_0_53_417 ();
 sg13g2_decap_8 FILLER_0_53_424 ();
 sg13g2_decap_8 FILLER_0_53_431 ();
 sg13g2_decap_8 FILLER_0_53_438 ();
 sg13g2_decap_8 FILLER_0_53_445 ();
 sg13g2_decap_8 FILLER_0_53_452 ();
 sg13g2_decap_4 FILLER_0_53_459 ();
 sg13g2_fill_2 FILLER_0_53_463 ();
 sg13g2_fill_1 FILLER_0_53_470 ();
 sg13g2_decap_8 FILLER_0_53_484 ();
 sg13g2_decap_4 FILLER_0_53_491 ();
 sg13g2_fill_2 FILLER_0_53_526 ();
 sg13g2_fill_1 FILLER_0_53_528 ();
 sg13g2_decap_8 FILLER_0_53_592 ();
 sg13g2_decap_8 FILLER_0_53_599 ();
 sg13g2_decap_4 FILLER_0_53_606 ();
 sg13g2_decap_8 FILLER_0_53_636 ();
 sg13g2_decap_4 FILLER_0_53_643 ();
 sg13g2_fill_2 FILLER_0_53_647 ();
 sg13g2_fill_2 FILLER_0_53_653 ();
 sg13g2_fill_2 FILLER_0_53_673 ();
 sg13g2_fill_2 FILLER_0_53_698 ();
 sg13g2_fill_2 FILLER_0_53_714 ();
 sg13g2_decap_8 FILLER_0_53_721 ();
 sg13g2_fill_2 FILLER_0_53_728 ();
 sg13g2_decap_8 FILLER_0_53_761 ();
 sg13g2_fill_2 FILLER_0_53_773 ();
 sg13g2_fill_2 FILLER_0_53_779 ();
 sg13g2_fill_2 FILLER_0_53_789 ();
 sg13g2_fill_2 FILLER_0_53_801 ();
 sg13g2_fill_1 FILLER_0_53_803 ();
 sg13g2_fill_2 FILLER_0_53_808 ();
 sg13g2_fill_1 FILLER_0_53_810 ();
 sg13g2_decap_4 FILLER_0_53_816 ();
 sg13g2_fill_2 FILLER_0_53_820 ();
 sg13g2_fill_2 FILLER_0_53_848 ();
 sg13g2_fill_1 FILLER_0_53_854 ();
 sg13g2_fill_2 FILLER_0_53_869 ();
 sg13g2_fill_2 FILLER_0_53_895 ();
 sg13g2_decap_8 FILLER_0_53_927 ();
 sg13g2_decap_8 FILLER_0_53_934 ();
 sg13g2_decap_8 FILLER_0_53_941 ();
 sg13g2_decap_8 FILLER_0_53_948 ();
 sg13g2_decap_8 FILLER_0_53_955 ();
 sg13g2_decap_4 FILLER_0_53_962 ();
 sg13g2_fill_2 FILLER_0_53_1011 ();
 sg13g2_fill_1 FILLER_0_53_1052 ();
 sg13g2_decap_8 FILLER_0_53_1063 ();
 sg13g2_decap_8 FILLER_0_53_1070 ();
 sg13g2_decap_8 FILLER_0_53_1077 ();
 sg13g2_decap_4 FILLER_0_53_1084 ();
 sg13g2_fill_2 FILLER_0_53_1088 ();
 sg13g2_decap_8 FILLER_0_53_1117 ();
 sg13g2_decap_8 FILLER_0_53_1124 ();
 sg13g2_decap_8 FILLER_0_53_1131 ();
 sg13g2_decap_8 FILLER_0_53_1138 ();
 sg13g2_decap_8 FILLER_0_53_1145 ();
 sg13g2_decap_8 FILLER_0_53_1152 ();
 sg13g2_decap_8 FILLER_0_53_1159 ();
 sg13g2_decap_8 FILLER_0_53_1166 ();
 sg13g2_decap_8 FILLER_0_53_1173 ();
 sg13g2_decap_8 FILLER_0_53_1180 ();
 sg13g2_decap_8 FILLER_0_53_1187 ();
 sg13g2_decap_8 FILLER_0_53_1194 ();
 sg13g2_decap_8 FILLER_0_53_1201 ();
 sg13g2_decap_8 FILLER_0_53_1208 ();
 sg13g2_decap_8 FILLER_0_53_1215 ();
 sg13g2_decap_4 FILLER_0_53_1222 ();
 sg13g2_fill_2 FILLER_0_53_1226 ();
 sg13g2_decap_8 FILLER_0_54_0 ();
 sg13g2_decap_8 FILLER_0_54_7 ();
 sg13g2_decap_8 FILLER_0_54_14 ();
 sg13g2_decap_8 FILLER_0_54_21 ();
 sg13g2_decap_8 FILLER_0_54_28 ();
 sg13g2_decap_8 FILLER_0_54_35 ();
 sg13g2_decap_8 FILLER_0_54_47 ();
 sg13g2_fill_2 FILLER_0_54_54 ();
 sg13g2_fill_1 FILLER_0_54_56 ();
 sg13g2_fill_1 FILLER_0_54_101 ();
 sg13g2_fill_1 FILLER_0_54_112 ();
 sg13g2_fill_1 FILLER_0_54_149 ();
 sg13g2_fill_2 FILLER_0_54_186 ();
 sg13g2_fill_1 FILLER_0_54_188 ();
 sg13g2_fill_2 FILLER_0_54_210 ();
 sg13g2_decap_8 FILLER_0_54_216 ();
 sg13g2_decap_8 FILLER_0_54_223 ();
 sg13g2_decap_8 FILLER_0_54_230 ();
 sg13g2_decap_8 FILLER_0_54_237 ();
 sg13g2_decap_8 FILLER_0_54_244 ();
 sg13g2_decap_8 FILLER_0_54_251 ();
 sg13g2_decap_8 FILLER_0_54_258 ();
 sg13g2_decap_8 FILLER_0_54_265 ();
 sg13g2_decap_8 FILLER_0_54_272 ();
 sg13g2_decap_8 FILLER_0_54_279 ();
 sg13g2_decap_8 FILLER_0_54_286 ();
 sg13g2_decap_8 FILLER_0_54_293 ();
 sg13g2_decap_8 FILLER_0_54_300 ();
 sg13g2_decap_8 FILLER_0_54_307 ();
 sg13g2_decap_8 FILLER_0_54_314 ();
 sg13g2_decap_8 FILLER_0_54_321 ();
 sg13g2_decap_8 FILLER_0_54_328 ();
 sg13g2_decap_4 FILLER_0_54_335 ();
 sg13g2_decap_8 FILLER_0_54_343 ();
 sg13g2_decap_4 FILLER_0_54_350 ();
 sg13g2_fill_1 FILLER_0_54_354 ();
 sg13g2_decap_4 FILLER_0_54_392 ();
 sg13g2_fill_2 FILLER_0_54_396 ();
 sg13g2_decap_8 FILLER_0_54_402 ();
 sg13g2_decap_8 FILLER_0_54_409 ();
 sg13g2_fill_1 FILLER_0_54_416 ();
 sg13g2_decap_8 FILLER_0_54_443 ();
 sg13g2_decap_4 FILLER_0_54_450 ();
 sg13g2_fill_2 FILLER_0_54_454 ();
 sg13g2_decap_8 FILLER_0_54_494 ();
 sg13g2_decap_4 FILLER_0_54_501 ();
 sg13g2_fill_2 FILLER_0_54_505 ();
 sg13g2_decap_4 FILLER_0_54_511 ();
 sg13g2_fill_1 FILLER_0_54_515 ();
 sg13g2_fill_2 FILLER_0_54_542 ();
 sg13g2_decap_8 FILLER_0_54_596 ();
 sg13g2_decap_8 FILLER_0_54_603 ();
 sg13g2_decap_8 FILLER_0_54_610 ();
 sg13g2_decap_8 FILLER_0_54_617 ();
 sg13g2_decap_8 FILLER_0_54_624 ();
 sg13g2_decap_8 FILLER_0_54_631 ();
 sg13g2_fill_2 FILLER_0_54_638 ();
 sg13g2_fill_1 FILLER_0_54_640 ();
 sg13g2_decap_8 FILLER_0_54_672 ();
 sg13g2_fill_2 FILLER_0_54_679 ();
 sg13g2_fill_2 FILLER_0_54_712 ();
 sg13g2_fill_2 FILLER_0_54_766 ();
 sg13g2_fill_1 FILLER_0_54_768 ();
 sg13g2_fill_2 FILLER_0_54_804 ();
 sg13g2_decap_8 FILLER_0_54_817 ();
 sg13g2_decap_4 FILLER_0_54_824 ();
 sg13g2_fill_1 FILLER_0_54_828 ();
 sg13g2_decap_4 FILLER_0_54_833 ();
 sg13g2_fill_2 FILLER_0_54_837 ();
 sg13g2_decap_8 FILLER_0_54_843 ();
 sg13g2_decap_8 FILLER_0_54_850 ();
 sg13g2_fill_2 FILLER_0_54_857 ();
 sg13g2_decap_4 FILLER_0_54_864 ();
 sg13g2_fill_1 FILLER_0_54_868 ();
 sg13g2_fill_2 FILLER_0_54_877 ();
 sg13g2_fill_2 FILLER_0_54_893 ();
 sg13g2_fill_1 FILLER_0_54_895 ();
 sg13g2_fill_2 FILLER_0_54_906 ();
 sg13g2_decap_8 FILLER_0_54_918 ();
 sg13g2_decap_8 FILLER_0_54_925 ();
 sg13g2_decap_8 FILLER_0_54_932 ();
 sg13g2_decap_8 FILLER_0_54_939 ();
 sg13g2_fill_1 FILLER_0_54_946 ();
 sg13g2_fill_2 FILLER_0_54_964 ();
 sg13g2_fill_1 FILLER_0_54_966 ();
 sg13g2_decap_4 FILLER_0_54_986 ();
 sg13g2_decap_8 FILLER_0_54_1002 ();
 sg13g2_fill_2 FILLER_0_54_1009 ();
 sg13g2_fill_2 FILLER_0_54_1016 ();
 sg13g2_fill_1 FILLER_0_54_1018 ();
 sg13g2_fill_2 FILLER_0_54_1023 ();
 sg13g2_fill_2 FILLER_0_54_1035 ();
 sg13g2_decap_4 FILLER_0_54_1040 ();
 sg13g2_decap_8 FILLER_0_54_1048 ();
 sg13g2_decap_4 FILLER_0_54_1055 ();
 sg13g2_fill_1 FILLER_0_54_1059 ();
 sg13g2_decap_8 FILLER_0_54_1065 ();
 sg13g2_fill_1 FILLER_0_54_1072 ();
 sg13g2_decap_8 FILLER_0_54_1078 ();
 sg13g2_fill_2 FILLER_0_54_1085 ();
 sg13g2_fill_1 FILLER_0_54_1087 ();
 sg13g2_decap_8 FILLER_0_54_1118 ();
 sg13g2_decap_8 FILLER_0_54_1125 ();
 sg13g2_decap_8 FILLER_0_54_1132 ();
 sg13g2_decap_8 FILLER_0_54_1139 ();
 sg13g2_decap_8 FILLER_0_54_1146 ();
 sg13g2_decap_8 FILLER_0_54_1153 ();
 sg13g2_decap_8 FILLER_0_54_1160 ();
 sg13g2_decap_8 FILLER_0_54_1167 ();
 sg13g2_decap_8 FILLER_0_54_1174 ();
 sg13g2_decap_8 FILLER_0_54_1181 ();
 sg13g2_decap_8 FILLER_0_54_1188 ();
 sg13g2_decap_8 FILLER_0_54_1195 ();
 sg13g2_decap_8 FILLER_0_54_1202 ();
 sg13g2_decap_8 FILLER_0_54_1209 ();
 sg13g2_decap_8 FILLER_0_54_1216 ();
 sg13g2_decap_4 FILLER_0_54_1223 ();
 sg13g2_fill_1 FILLER_0_54_1227 ();
 sg13g2_decap_8 FILLER_0_55_0 ();
 sg13g2_decap_8 FILLER_0_55_7 ();
 sg13g2_decap_8 FILLER_0_55_14 ();
 sg13g2_decap_8 FILLER_0_55_21 ();
 sg13g2_decap_8 FILLER_0_55_28 ();
 sg13g2_decap_8 FILLER_0_55_35 ();
 sg13g2_decap_8 FILLER_0_55_42 ();
 sg13g2_decap_8 FILLER_0_55_49 ();
 sg13g2_decap_8 FILLER_0_55_56 ();
 sg13g2_decap_8 FILLER_0_55_63 ();
 sg13g2_decap_8 FILLER_0_55_70 ();
 sg13g2_fill_1 FILLER_0_55_77 ();
 sg13g2_decap_4 FILLER_0_55_91 ();
 sg13g2_fill_2 FILLER_0_55_103 ();
 sg13g2_fill_2 FILLER_0_55_110 ();
 sg13g2_fill_2 FILLER_0_55_117 ();
 sg13g2_fill_2 FILLER_0_55_124 ();
 sg13g2_fill_2 FILLER_0_55_130 ();
 sg13g2_fill_1 FILLER_0_55_132 ();
 sg13g2_decap_8 FILLER_0_55_137 ();
 sg13g2_fill_1 FILLER_0_55_144 ();
 sg13g2_fill_2 FILLER_0_55_157 ();
 sg13g2_fill_1 FILLER_0_55_159 ();
 sg13g2_decap_4 FILLER_0_55_191 ();
 sg13g2_fill_2 FILLER_0_55_195 ();
 sg13g2_decap_8 FILLER_0_55_228 ();
 sg13g2_decap_8 FILLER_0_55_235 ();
 sg13g2_decap_8 FILLER_0_55_242 ();
 sg13g2_decap_8 FILLER_0_55_249 ();
 sg13g2_decap_8 FILLER_0_55_256 ();
 sg13g2_decap_8 FILLER_0_55_263 ();
 sg13g2_decap_8 FILLER_0_55_270 ();
 sg13g2_decap_8 FILLER_0_55_277 ();
 sg13g2_decap_8 FILLER_0_55_284 ();
 sg13g2_decap_8 FILLER_0_55_291 ();
 sg13g2_decap_8 FILLER_0_55_298 ();
 sg13g2_decap_8 FILLER_0_55_305 ();
 sg13g2_decap_8 FILLER_0_55_312 ();
 sg13g2_decap_8 FILLER_0_55_319 ();
 sg13g2_decap_8 FILLER_0_55_326 ();
 sg13g2_decap_8 FILLER_0_55_333 ();
 sg13g2_decap_8 FILLER_0_55_340 ();
 sg13g2_decap_8 FILLER_0_55_352 ();
 sg13g2_decap_8 FILLER_0_55_359 ();
 sg13g2_decap_8 FILLER_0_55_366 ();
 sg13g2_fill_1 FILLER_0_55_373 ();
 sg13g2_decap_8 FILLER_0_55_378 ();
 sg13g2_decap_8 FILLER_0_55_385 ();
 sg13g2_decap_8 FILLER_0_55_392 ();
 sg13g2_decap_4 FILLER_0_55_399 ();
 sg13g2_fill_2 FILLER_0_55_403 ();
 sg13g2_decap_4 FILLER_0_55_409 ();
 sg13g2_fill_2 FILLER_0_55_423 ();
 sg13g2_fill_1 FILLER_0_55_425 ();
 sg13g2_decap_4 FILLER_0_55_430 ();
 sg13g2_fill_2 FILLER_0_55_524 ();
 sg13g2_fill_1 FILLER_0_55_526 ();
 sg13g2_fill_1 FILLER_0_55_531 ();
 sg13g2_decap_8 FILLER_0_55_550 ();
 sg13g2_fill_2 FILLER_0_55_557 ();
 sg13g2_fill_2 FILLER_0_55_569 ();
 sg13g2_fill_1 FILLER_0_55_571 ();
 sg13g2_fill_2 FILLER_0_55_582 ();
 sg13g2_fill_1 FILLER_0_55_584 ();
 sg13g2_decap_8 FILLER_0_55_595 ();
 sg13g2_fill_2 FILLER_0_55_602 ();
 sg13g2_decap_8 FILLER_0_55_616 ();
 sg13g2_decap_8 FILLER_0_55_623 ();
 sg13g2_decap_8 FILLER_0_55_630 ();
 sg13g2_decap_4 FILLER_0_55_637 ();
 sg13g2_decap_8 FILLER_0_55_645 ();
 sg13g2_decap_8 FILLER_0_55_652 ();
 sg13g2_decap_8 FILLER_0_55_659 ();
 sg13g2_decap_8 FILLER_0_55_666 ();
 sg13g2_decap_8 FILLER_0_55_673 ();
 sg13g2_decap_8 FILLER_0_55_680 ();
 sg13g2_decap_4 FILLER_0_55_687 ();
 sg13g2_fill_2 FILLER_0_55_691 ();
 sg13g2_fill_2 FILLER_0_55_727 ();
 sg13g2_fill_2 FILLER_0_55_749 ();
 sg13g2_fill_1 FILLER_0_55_751 ();
 sg13g2_decap_4 FILLER_0_55_756 ();
 sg13g2_decap_8 FILLER_0_55_770 ();
 sg13g2_fill_2 FILLER_0_55_777 ();
 sg13g2_decap_4 FILLER_0_55_784 ();
 sg13g2_fill_1 FILLER_0_55_788 ();
 sg13g2_fill_1 FILLER_0_55_799 ();
 sg13g2_decap_8 FILLER_0_55_805 ();
 sg13g2_decap_8 FILLER_0_55_812 ();
 sg13g2_decap_4 FILLER_0_55_823 ();
 sg13g2_fill_1 FILLER_0_55_827 ();
 sg13g2_decap_8 FILLER_0_55_833 ();
 sg13g2_decap_8 FILLER_0_55_840 ();
 sg13g2_decap_8 FILLER_0_55_847 ();
 sg13g2_fill_2 FILLER_0_55_854 ();
 sg13g2_fill_1 FILLER_0_55_856 ();
 sg13g2_fill_2 FILLER_0_55_862 ();
 sg13g2_decap_8 FILLER_0_55_868 ();
 sg13g2_fill_1 FILLER_0_55_875 ();
 sg13g2_fill_2 FILLER_0_55_881 ();
 sg13g2_decap_8 FILLER_0_55_888 ();
 sg13g2_decap_8 FILLER_0_55_895 ();
 sg13g2_fill_1 FILLER_0_55_902 ();
 sg13g2_fill_1 FILLER_0_55_907 ();
 sg13g2_decap_8 FILLER_0_55_923 ();
 sg13g2_decap_8 FILLER_0_55_930 ();
 sg13g2_decap_8 FILLER_0_55_937 ();
 sg13g2_decap_8 FILLER_0_55_944 ();
 sg13g2_decap_8 FILLER_0_55_951 ();
 sg13g2_decap_8 FILLER_0_55_984 ();
 sg13g2_decap_8 FILLER_0_55_991 ();
 sg13g2_fill_1 FILLER_0_55_998 ();
 sg13g2_fill_2 FILLER_0_55_1009 ();
 sg13g2_fill_1 FILLER_0_55_1011 ();
 sg13g2_fill_1 FILLER_0_55_1038 ();
 sg13g2_fill_1 FILLER_0_55_1044 ();
 sg13g2_fill_1 FILLER_0_55_1071 ();
 sg13g2_fill_1 FILLER_0_55_1098 ();
 sg13g2_decap_8 FILLER_0_55_1114 ();
 sg13g2_decap_8 FILLER_0_55_1121 ();
 sg13g2_decap_8 FILLER_0_55_1128 ();
 sg13g2_decap_8 FILLER_0_55_1135 ();
 sg13g2_decap_8 FILLER_0_55_1142 ();
 sg13g2_decap_8 FILLER_0_55_1149 ();
 sg13g2_decap_8 FILLER_0_55_1156 ();
 sg13g2_decap_8 FILLER_0_55_1163 ();
 sg13g2_decap_8 FILLER_0_55_1170 ();
 sg13g2_decap_8 FILLER_0_55_1177 ();
 sg13g2_decap_8 FILLER_0_55_1184 ();
 sg13g2_decap_8 FILLER_0_55_1191 ();
 sg13g2_decap_8 FILLER_0_55_1198 ();
 sg13g2_decap_8 FILLER_0_55_1205 ();
 sg13g2_decap_8 FILLER_0_55_1212 ();
 sg13g2_decap_8 FILLER_0_55_1219 ();
 sg13g2_fill_2 FILLER_0_55_1226 ();
 sg13g2_decap_8 FILLER_0_56_0 ();
 sg13g2_decap_8 FILLER_0_56_7 ();
 sg13g2_decap_8 FILLER_0_56_14 ();
 sg13g2_decap_8 FILLER_0_56_21 ();
 sg13g2_decap_8 FILLER_0_56_28 ();
 sg13g2_decap_8 FILLER_0_56_35 ();
 sg13g2_decap_8 FILLER_0_56_42 ();
 sg13g2_fill_2 FILLER_0_56_49 ();
 sg13g2_fill_1 FILLER_0_56_51 ();
 sg13g2_fill_1 FILLER_0_56_109 ();
 sg13g2_decap_8 FILLER_0_56_141 ();
 sg13g2_fill_2 FILLER_0_56_148 ();
 sg13g2_decap_4 FILLER_0_56_154 ();
 sg13g2_fill_2 FILLER_0_56_158 ();
 sg13g2_fill_1 FILLER_0_56_189 ();
 sg13g2_decap_4 FILLER_0_56_205 ();
 sg13g2_fill_1 FILLER_0_56_209 ();
 sg13g2_decap_8 FILLER_0_56_218 ();
 sg13g2_decap_8 FILLER_0_56_225 ();
 sg13g2_decap_8 FILLER_0_56_232 ();
 sg13g2_decap_8 FILLER_0_56_239 ();
 sg13g2_decap_8 FILLER_0_56_246 ();
 sg13g2_decap_8 FILLER_0_56_253 ();
 sg13g2_decap_8 FILLER_0_56_260 ();
 sg13g2_decap_8 FILLER_0_56_267 ();
 sg13g2_decap_8 FILLER_0_56_274 ();
 sg13g2_decap_8 FILLER_0_56_281 ();
 sg13g2_decap_8 FILLER_0_56_288 ();
 sg13g2_decap_8 FILLER_0_56_295 ();
 sg13g2_decap_8 FILLER_0_56_302 ();
 sg13g2_decap_8 FILLER_0_56_309 ();
 sg13g2_fill_1 FILLER_0_56_316 ();
 sg13g2_fill_1 FILLER_0_56_336 ();
 sg13g2_decap_4 FILLER_0_56_363 ();
 sg13g2_fill_1 FILLER_0_56_367 ();
 sg13g2_fill_2 FILLER_0_56_372 ();
 sg13g2_decap_4 FILLER_0_56_379 ();
 sg13g2_fill_1 FILLER_0_56_423 ();
 sg13g2_fill_2 FILLER_0_56_439 ();
 sg13g2_fill_2 FILLER_0_56_445 ();
 sg13g2_fill_1 FILLER_0_56_447 ();
 sg13g2_decap_8 FILLER_0_56_458 ();
 sg13g2_decap_8 FILLER_0_56_465 ();
 sg13g2_fill_1 FILLER_0_56_472 ();
 sg13g2_decap_8 FILLER_0_56_492 ();
 sg13g2_decap_8 FILLER_0_56_499 ();
 sg13g2_decap_8 FILLER_0_56_506 ();
 sg13g2_decap_4 FILLER_0_56_513 ();
 sg13g2_fill_1 FILLER_0_56_517 ();
 sg13g2_decap_8 FILLER_0_56_544 ();
 sg13g2_decap_8 FILLER_0_56_551 ();
 sg13g2_decap_8 FILLER_0_56_558 ();
 sg13g2_decap_4 FILLER_0_56_565 ();
 sg13g2_fill_1 FILLER_0_56_569 ();
 sg13g2_fill_2 FILLER_0_56_575 ();
 sg13g2_fill_1 FILLER_0_56_577 ();
 sg13g2_fill_1 FILLER_0_56_604 ();
 sg13g2_fill_2 FILLER_0_56_621 ();
 sg13g2_fill_1 FILLER_0_56_623 ();
 sg13g2_decap_4 FILLER_0_56_660 ();
 sg13g2_fill_1 FILLER_0_56_664 ();
 sg13g2_decap_4 FILLER_0_56_674 ();
 sg13g2_fill_2 FILLER_0_56_678 ();
 sg13g2_decap_8 FILLER_0_56_685 ();
 sg13g2_fill_2 FILLER_0_56_692 ();
 sg13g2_fill_1 FILLER_0_56_694 ();
 sg13g2_fill_1 FILLER_0_56_700 ();
 sg13g2_fill_1 FILLER_0_56_711 ();
 sg13g2_fill_2 FILLER_0_56_727 ();
 sg13g2_fill_1 FILLER_0_56_729 ();
 sg13g2_fill_1 FILLER_0_56_743 ();
 sg13g2_decap_4 FILLER_0_56_748 ();
 sg13g2_decap_4 FILLER_0_56_767 ();
 sg13g2_fill_1 FILLER_0_56_771 ();
 sg13g2_fill_1 FILLER_0_56_776 ();
 sg13g2_fill_1 FILLER_0_56_863 ();
 sg13g2_fill_1 FILLER_0_56_890 ();
 sg13g2_fill_1 FILLER_0_56_901 ();
 sg13g2_fill_1 FILLER_0_56_938 ();
 sg13g2_decap_8 FILLER_0_56_943 ();
 sg13g2_decap_8 FILLER_0_56_950 ();
 sg13g2_decap_8 FILLER_0_56_957 ();
 sg13g2_fill_2 FILLER_0_56_964 ();
 sg13g2_fill_1 FILLER_0_56_966 ();
 sg13g2_fill_2 FILLER_0_56_987 ();
 sg13g2_decap_4 FILLER_0_56_1020 ();
 sg13g2_decap_8 FILLER_0_56_1029 ();
 sg13g2_fill_1 FILLER_0_56_1036 ();
 sg13g2_fill_1 FILLER_0_56_1047 ();
 sg13g2_fill_1 FILLER_0_56_1056 ();
 sg13g2_fill_1 FILLER_0_56_1067 ();
 sg13g2_fill_1 FILLER_0_56_1078 ();
 sg13g2_decap_8 FILLER_0_56_1083 ();
 sg13g2_fill_1 FILLER_0_56_1090 ();
 sg13g2_fill_1 FILLER_0_56_1121 ();
 sg13g2_decap_8 FILLER_0_56_1132 ();
 sg13g2_decap_8 FILLER_0_56_1139 ();
 sg13g2_decap_8 FILLER_0_56_1146 ();
 sg13g2_decap_8 FILLER_0_56_1153 ();
 sg13g2_decap_8 FILLER_0_56_1160 ();
 sg13g2_decap_8 FILLER_0_56_1167 ();
 sg13g2_decap_8 FILLER_0_56_1174 ();
 sg13g2_decap_8 FILLER_0_56_1181 ();
 sg13g2_decap_8 FILLER_0_56_1188 ();
 sg13g2_decap_8 FILLER_0_56_1195 ();
 sg13g2_decap_8 FILLER_0_56_1202 ();
 sg13g2_decap_8 FILLER_0_56_1209 ();
 sg13g2_decap_8 FILLER_0_56_1216 ();
 sg13g2_decap_4 FILLER_0_56_1223 ();
 sg13g2_fill_1 FILLER_0_56_1227 ();
 sg13g2_decap_8 FILLER_0_57_0 ();
 sg13g2_decap_8 FILLER_0_57_7 ();
 sg13g2_decap_8 FILLER_0_57_14 ();
 sg13g2_decap_8 FILLER_0_57_21 ();
 sg13g2_decap_8 FILLER_0_57_28 ();
 sg13g2_decap_8 FILLER_0_57_35 ();
 sg13g2_decap_8 FILLER_0_57_42 ();
 sg13g2_decap_8 FILLER_0_57_176 ();
 sg13g2_decap_8 FILLER_0_57_183 ();
 sg13g2_decap_8 FILLER_0_57_190 ();
 sg13g2_decap_4 FILLER_0_57_197 ();
 sg13g2_fill_1 FILLER_0_57_206 ();
 sg13g2_decap_8 FILLER_0_57_233 ();
 sg13g2_decap_8 FILLER_0_57_240 ();
 sg13g2_decap_8 FILLER_0_57_247 ();
 sg13g2_decap_8 FILLER_0_57_254 ();
 sg13g2_decap_8 FILLER_0_57_261 ();
 sg13g2_decap_8 FILLER_0_57_268 ();
 sg13g2_decap_8 FILLER_0_57_275 ();
 sg13g2_decap_8 FILLER_0_57_282 ();
 sg13g2_decap_8 FILLER_0_57_289 ();
 sg13g2_decap_4 FILLER_0_57_296 ();
 sg13g2_fill_1 FILLER_0_57_300 ();
 sg13g2_fill_2 FILLER_0_57_306 ();
 sg13g2_fill_1 FILLER_0_57_308 ();
 sg13g2_fill_1 FILLER_0_57_375 ();
 sg13g2_fill_1 FILLER_0_57_402 ();
 sg13g2_fill_2 FILLER_0_57_413 ();
 sg13g2_decap_8 FILLER_0_57_469 ();
 sg13g2_decap_8 FILLER_0_57_480 ();
 sg13g2_decap_8 FILLER_0_57_487 ();
 sg13g2_decap_8 FILLER_0_57_494 ();
 sg13g2_decap_8 FILLER_0_57_501 ();
 sg13g2_decap_8 FILLER_0_57_508 ();
 sg13g2_decap_4 FILLER_0_57_515 ();
 sg13g2_decap_8 FILLER_0_57_523 ();
 sg13g2_fill_2 FILLER_0_57_530 ();
 sg13g2_fill_1 FILLER_0_57_532 ();
 sg13g2_decap_8 FILLER_0_57_543 ();
 sg13g2_decap_8 FILLER_0_57_554 ();
 sg13g2_decap_8 FILLER_0_57_561 ();
 sg13g2_decap_8 FILLER_0_57_568 ();
 sg13g2_decap_8 FILLER_0_57_575 ();
 sg13g2_fill_2 FILLER_0_57_582 ();
 sg13g2_fill_2 FILLER_0_57_589 ();
 sg13g2_fill_1 FILLER_0_57_591 ();
 sg13g2_decap_8 FILLER_0_57_602 ();
 sg13g2_fill_1 FILLER_0_57_609 ();
 sg13g2_decap_4 FILLER_0_57_698 ();
 sg13g2_fill_2 FILLER_0_57_702 ();
 sg13g2_decap_8 FILLER_0_57_708 ();
 sg13g2_decap_8 FILLER_0_57_715 ();
 sg13g2_decap_4 FILLER_0_57_722 ();
 sg13g2_fill_1 FILLER_0_57_726 ();
 sg13g2_decap_4 FILLER_0_57_732 ();
 sg13g2_fill_1 FILLER_0_57_740 ();
 sg13g2_fill_1 FILLER_0_57_745 ();
 sg13g2_fill_1 FILLER_0_57_798 ();
 sg13g2_fill_1 FILLER_0_57_825 ();
 sg13g2_fill_2 FILLER_0_57_852 ();
 sg13g2_fill_1 FILLER_0_57_880 ();
 sg13g2_fill_2 FILLER_0_57_907 ();
 sg13g2_fill_2 FILLER_0_57_918 ();
 sg13g2_fill_2 FILLER_0_57_956 ();
 sg13g2_decap_4 FILLER_0_57_984 ();
 sg13g2_decap_4 FILLER_0_57_992 ();
 sg13g2_fill_1 FILLER_0_57_996 ();
 sg13g2_fill_2 FILLER_0_57_1057 ();
 sg13g2_fill_1 FILLER_0_57_1089 ();
 sg13g2_decap_8 FILLER_0_57_1125 ();
 sg13g2_decap_8 FILLER_0_57_1132 ();
 sg13g2_decap_8 FILLER_0_57_1139 ();
 sg13g2_decap_8 FILLER_0_57_1146 ();
 sg13g2_decap_8 FILLER_0_57_1153 ();
 sg13g2_decap_8 FILLER_0_57_1160 ();
 sg13g2_decap_8 FILLER_0_57_1167 ();
 sg13g2_decap_8 FILLER_0_57_1174 ();
 sg13g2_decap_8 FILLER_0_57_1181 ();
 sg13g2_decap_8 FILLER_0_57_1188 ();
 sg13g2_decap_8 FILLER_0_57_1195 ();
 sg13g2_decap_8 FILLER_0_57_1202 ();
 sg13g2_decap_8 FILLER_0_57_1209 ();
 sg13g2_decap_8 FILLER_0_57_1216 ();
 sg13g2_decap_4 FILLER_0_57_1223 ();
 sg13g2_fill_1 FILLER_0_57_1227 ();
 sg13g2_decap_8 FILLER_0_58_0 ();
 sg13g2_decap_8 FILLER_0_58_7 ();
 sg13g2_decap_8 FILLER_0_58_14 ();
 sg13g2_decap_8 FILLER_0_58_21 ();
 sg13g2_decap_8 FILLER_0_58_28 ();
 sg13g2_decap_8 FILLER_0_58_35 ();
 sg13g2_decap_8 FILLER_0_58_42 ();
 sg13g2_decap_8 FILLER_0_58_49 ();
 sg13g2_fill_2 FILLER_0_58_56 ();
 sg13g2_fill_1 FILLER_0_58_58 ();
 sg13g2_fill_2 FILLER_0_58_69 ();
 sg13g2_fill_2 FILLER_0_58_85 ();
 sg13g2_fill_1 FILLER_0_58_87 ();
 sg13g2_fill_1 FILLER_0_58_98 ();
 sg13g2_fill_1 FILLER_0_58_113 ();
 sg13g2_fill_2 FILLER_0_58_124 ();
 sg13g2_decap_8 FILLER_0_58_146 ();
 sg13g2_decap_8 FILLER_0_58_153 ();
 sg13g2_fill_2 FILLER_0_58_160 ();
 sg13g2_decap_8 FILLER_0_58_183 ();
 sg13g2_decap_8 FILLER_0_58_190 ();
 sg13g2_decap_8 FILLER_0_58_197 ();
 sg13g2_decap_8 FILLER_0_58_204 ();
 sg13g2_decap_8 FILLER_0_58_211 ();
 sg13g2_fill_1 FILLER_0_58_218 ();
 sg13g2_fill_1 FILLER_0_58_223 ();
 sg13g2_decap_8 FILLER_0_58_227 ();
 sg13g2_fill_1 FILLER_0_58_234 ();
 sg13g2_fill_1 FILLER_0_58_245 ();
 sg13g2_decap_4 FILLER_0_58_272 ();
 sg13g2_fill_2 FILLER_0_58_276 ();
 sg13g2_fill_1 FILLER_0_58_304 ();
 sg13g2_fill_2 FILLER_0_58_331 ();
 sg13g2_fill_1 FILLER_0_58_333 ();
 sg13g2_fill_2 FILLER_0_58_349 ();
 sg13g2_fill_1 FILLER_0_58_387 ();
 sg13g2_decap_8 FILLER_0_58_414 ();
 sg13g2_decap_8 FILLER_0_58_421 ();
 sg13g2_decap_8 FILLER_0_58_428 ();
 sg13g2_decap_4 FILLER_0_58_435 ();
 sg13g2_fill_1 FILLER_0_58_439 ();
 sg13g2_fill_2 FILLER_0_58_444 ();
 sg13g2_fill_2 FILLER_0_58_450 ();
 sg13g2_fill_1 FILLER_0_58_462 ();
 sg13g2_fill_2 FILLER_0_58_504 ();
 sg13g2_fill_2 FILLER_0_58_540 ();
 sg13g2_fill_1 FILLER_0_58_542 ();
 sg13g2_decap_4 FILLER_0_58_569 ();
 sg13g2_fill_1 FILLER_0_58_603 ();
 sg13g2_fill_1 FILLER_0_58_609 ();
 sg13g2_fill_1 FILLER_0_58_634 ();
 sg13g2_fill_2 FILLER_0_58_645 ();
 sg13g2_fill_1 FILLER_0_58_647 ();
 sg13g2_decap_4 FILLER_0_58_710 ();
 sg13g2_fill_1 FILLER_0_58_714 ();
 sg13g2_fill_2 FILLER_0_58_745 ();
 sg13g2_fill_1 FILLER_0_58_789 ();
 sg13g2_fill_1 FILLER_0_58_800 ();
 sg13g2_fill_2 FILLER_0_58_840 ();
 sg13g2_fill_2 FILLER_0_58_886 ();
 sg13g2_fill_1 FILLER_0_58_888 ();
 sg13g2_fill_1 FILLER_0_58_915 ();
 sg13g2_fill_1 FILLER_0_58_926 ();
 sg13g2_fill_1 FILLER_0_58_932 ();
 sg13g2_decap_4 FILLER_0_58_968 ();
 sg13g2_decap_4 FILLER_0_58_977 ();
 sg13g2_decap_4 FILLER_0_58_985 ();
 sg13g2_decap_4 FILLER_0_58_1004 ();
 sg13g2_decap_4 FILLER_0_58_1018 ();
 sg13g2_fill_2 FILLER_0_58_1035 ();
 sg13g2_decap_4 FILLER_0_58_1047 ();
 sg13g2_fill_1 FILLER_0_58_1051 ();
 sg13g2_decap_4 FILLER_0_58_1056 ();
 sg13g2_fill_1 FILLER_0_58_1060 ();
 sg13g2_fill_2 FILLER_0_58_1066 ();
 sg13g2_fill_1 FILLER_0_58_1068 ();
 sg13g2_decap_8 FILLER_0_58_1079 ();
 sg13g2_decap_8 FILLER_0_58_1086 ();
 sg13g2_decap_8 FILLER_0_58_1093 ();
 sg13g2_decap_4 FILLER_0_58_1100 ();
 sg13g2_fill_1 FILLER_0_58_1104 ();
 sg13g2_decap_4 FILLER_0_58_1113 ();
 sg13g2_fill_2 FILLER_0_58_1117 ();
 sg13g2_decap_8 FILLER_0_58_1129 ();
 sg13g2_decap_8 FILLER_0_58_1136 ();
 sg13g2_decap_8 FILLER_0_58_1143 ();
 sg13g2_decap_8 FILLER_0_58_1150 ();
 sg13g2_decap_8 FILLER_0_58_1157 ();
 sg13g2_decap_8 FILLER_0_58_1164 ();
 sg13g2_decap_8 FILLER_0_58_1171 ();
 sg13g2_decap_8 FILLER_0_58_1178 ();
 sg13g2_decap_8 FILLER_0_58_1185 ();
 sg13g2_decap_8 FILLER_0_58_1192 ();
 sg13g2_decap_8 FILLER_0_58_1199 ();
 sg13g2_decap_8 FILLER_0_58_1206 ();
 sg13g2_decap_8 FILLER_0_58_1213 ();
 sg13g2_decap_8 FILLER_0_58_1220 ();
 sg13g2_fill_1 FILLER_0_58_1227 ();
 sg13g2_decap_8 FILLER_0_59_0 ();
 sg13g2_decap_8 FILLER_0_59_7 ();
 sg13g2_decap_8 FILLER_0_59_14 ();
 sg13g2_decap_8 FILLER_0_59_21 ();
 sg13g2_decap_8 FILLER_0_59_28 ();
 sg13g2_decap_4 FILLER_0_59_35 ();
 sg13g2_fill_1 FILLER_0_59_39 ();
 sg13g2_decap_8 FILLER_0_59_75 ();
 sg13g2_fill_1 FILLER_0_59_82 ();
 sg13g2_fill_2 FILLER_0_59_91 ();
 sg13g2_fill_1 FILLER_0_59_93 ();
 sg13g2_decap_8 FILLER_0_59_99 ();
 sg13g2_decap_4 FILLER_0_59_106 ();
 sg13g2_fill_1 FILLER_0_59_110 ();
 sg13g2_decap_8 FILLER_0_59_120 ();
 sg13g2_fill_2 FILLER_0_59_127 ();
 sg13g2_decap_8 FILLER_0_59_138 ();
 sg13g2_fill_2 FILLER_0_59_145 ();
 sg13g2_decap_4 FILLER_0_59_162 ();
 sg13g2_decap_4 FILLER_0_59_192 ();
 sg13g2_fill_1 FILLER_0_59_200 ();
 sg13g2_fill_1 FILLER_0_59_227 ();
 sg13g2_fill_1 FILLER_0_59_315 ();
 sg13g2_decap_8 FILLER_0_59_325 ();
 sg13g2_decap_4 FILLER_0_59_352 ();
 sg13g2_fill_1 FILLER_0_59_360 ();
 sg13g2_fill_1 FILLER_0_59_366 ();
 sg13g2_fill_1 FILLER_0_59_401 ();
 sg13g2_decap_8 FILLER_0_59_406 ();
 sg13g2_decap_8 FILLER_0_59_413 ();
 sg13g2_decap_8 FILLER_0_59_420 ();
 sg13g2_decap_8 FILLER_0_59_427 ();
 sg13g2_fill_1 FILLER_0_59_434 ();
 sg13g2_decap_4 FILLER_0_59_444 ();
 sg13g2_fill_1 FILLER_0_59_448 ();
 sg13g2_fill_2 FILLER_0_59_464 ();
 sg13g2_fill_1 FILLER_0_59_466 ();
 sg13g2_decap_4 FILLER_0_59_493 ();
 sg13g2_fill_2 FILLER_0_59_497 ();
 sg13g2_fill_2 FILLER_0_59_549 ();
 sg13g2_fill_1 FILLER_0_59_551 ();
 sg13g2_decap_4 FILLER_0_59_578 ();
 sg13g2_fill_1 FILLER_0_59_587 ();
 sg13g2_fill_1 FILLER_0_59_592 ();
 sg13g2_fill_1 FILLER_0_59_607 ();
 sg13g2_decap_8 FILLER_0_59_634 ();
 sg13g2_fill_1 FILLER_0_59_641 ();
 sg13g2_fill_2 FILLER_0_59_647 ();
 sg13g2_fill_1 FILLER_0_59_649 ();
 sg13g2_fill_2 FILLER_0_59_672 ();
 sg13g2_fill_1 FILLER_0_59_674 ();
 sg13g2_decap_4 FILLER_0_59_685 ();
 sg13g2_fill_2 FILLER_0_59_689 ();
 sg13g2_fill_1 FILLER_0_59_695 ();
 sg13g2_fill_1 FILLER_0_59_763 ();
 sg13g2_decap_8 FILLER_0_59_768 ();
 sg13g2_decap_4 FILLER_0_59_775 ();
 sg13g2_fill_1 FILLER_0_59_783 ();
 sg13g2_decap_8 FILLER_0_59_793 ();
 sg13g2_decap_8 FILLER_0_59_800 ();
 sg13g2_decap_8 FILLER_0_59_807 ();
 sg13g2_decap_8 FILLER_0_59_814 ();
 sg13g2_decap_8 FILLER_0_59_821 ();
 sg13g2_decap_8 FILLER_0_59_828 ();
 sg13g2_decap_8 FILLER_0_59_835 ();
 sg13g2_decap_4 FILLER_0_59_842 ();
 sg13g2_fill_1 FILLER_0_59_846 ();
 sg13g2_decap_4 FILLER_0_59_851 ();
 sg13g2_fill_1 FILLER_0_59_855 ();
 sg13g2_decap_8 FILLER_0_59_860 ();
 sg13g2_decap_8 FILLER_0_59_867 ();
 sg13g2_fill_1 FILLER_0_59_874 ();
 sg13g2_decap_4 FILLER_0_59_880 ();
 sg13g2_fill_2 FILLER_0_59_884 ();
 sg13g2_fill_1 FILLER_0_59_901 ();
 sg13g2_decap_8 FILLER_0_59_948 ();
 sg13g2_decap_8 FILLER_0_59_955 ();
 sg13g2_decap_8 FILLER_0_59_962 ();
 sg13g2_decap_4 FILLER_0_59_969 ();
 sg13g2_fill_1 FILLER_0_59_973 ();
 sg13g2_decap_8 FILLER_0_59_1000 ();
 sg13g2_decap_8 FILLER_0_59_1007 ();
 sg13g2_decap_8 FILLER_0_59_1014 ();
 sg13g2_decap_8 FILLER_0_59_1047 ();
 sg13g2_fill_1 FILLER_0_59_1054 ();
 sg13g2_fill_2 FILLER_0_59_1093 ();
 sg13g2_fill_1 FILLER_0_59_1095 ();
 sg13g2_decap_8 FILLER_0_59_1127 ();
 sg13g2_decap_8 FILLER_0_59_1134 ();
 sg13g2_decap_8 FILLER_0_59_1141 ();
 sg13g2_decap_8 FILLER_0_59_1148 ();
 sg13g2_decap_8 FILLER_0_59_1155 ();
 sg13g2_decap_8 FILLER_0_59_1162 ();
 sg13g2_decap_8 FILLER_0_59_1169 ();
 sg13g2_decap_8 FILLER_0_59_1176 ();
 sg13g2_decap_8 FILLER_0_59_1183 ();
 sg13g2_decap_8 FILLER_0_59_1190 ();
 sg13g2_decap_8 FILLER_0_59_1197 ();
 sg13g2_decap_8 FILLER_0_59_1204 ();
 sg13g2_decap_8 FILLER_0_59_1211 ();
 sg13g2_decap_8 FILLER_0_59_1218 ();
 sg13g2_fill_2 FILLER_0_59_1225 ();
 sg13g2_fill_1 FILLER_0_59_1227 ();
 sg13g2_decap_8 FILLER_0_60_0 ();
 sg13g2_decap_8 FILLER_0_60_7 ();
 sg13g2_decap_8 FILLER_0_60_14 ();
 sg13g2_decap_8 FILLER_0_60_21 ();
 sg13g2_decap_8 FILLER_0_60_28 ();
 sg13g2_decap_8 FILLER_0_60_35 ();
 sg13g2_decap_8 FILLER_0_60_42 ();
 sg13g2_decap_4 FILLER_0_60_49 ();
 sg13g2_decap_8 FILLER_0_60_57 ();
 sg13g2_decap_8 FILLER_0_60_69 ();
 sg13g2_decap_8 FILLER_0_60_76 ();
 sg13g2_decap_8 FILLER_0_60_83 ();
 sg13g2_decap_8 FILLER_0_60_90 ();
 sg13g2_decap_8 FILLER_0_60_97 ();
 sg13g2_decap_8 FILLER_0_60_104 ();
 sg13g2_decap_8 FILLER_0_60_111 ();
 sg13g2_decap_8 FILLER_0_60_118 ();
 sg13g2_decap_8 FILLER_0_60_125 ();
 sg13g2_decap_8 FILLER_0_60_132 ();
 sg13g2_decap_8 FILLER_0_60_139 ();
 sg13g2_fill_2 FILLER_0_60_146 ();
 sg13g2_fill_1 FILLER_0_60_148 ();
 sg13g2_decap_8 FILLER_0_60_185 ();
 sg13g2_fill_2 FILLER_0_60_245 ();
 sg13g2_fill_1 FILLER_0_60_247 ();
 sg13g2_fill_1 FILLER_0_60_253 ();
 sg13g2_fill_1 FILLER_0_60_264 ();
 sg13g2_decap_8 FILLER_0_60_308 ();
 sg13g2_decap_8 FILLER_0_60_315 ();
 sg13g2_decap_8 FILLER_0_60_322 ();
 sg13g2_fill_1 FILLER_0_60_329 ();
 sg13g2_decap_8 FILLER_0_60_334 ();
 sg13g2_decap_8 FILLER_0_60_341 ();
 sg13g2_decap_8 FILLER_0_60_348 ();
 sg13g2_decap_8 FILLER_0_60_355 ();
 sg13g2_decap_8 FILLER_0_60_362 ();
 sg13g2_decap_8 FILLER_0_60_369 ();
 sg13g2_decap_8 FILLER_0_60_376 ();
 sg13g2_decap_8 FILLER_0_60_394 ();
 sg13g2_decap_8 FILLER_0_60_401 ();
 sg13g2_decap_8 FILLER_0_60_408 ();
 sg13g2_decap_8 FILLER_0_60_415 ();
 sg13g2_decap_4 FILLER_0_60_422 ();
 sg13g2_decap_4 FILLER_0_60_460 ();
 sg13g2_decap_4 FILLER_0_60_541 ();
 sg13g2_decap_8 FILLER_0_60_564 ();
 sg13g2_decap_8 FILLER_0_60_571 ();
 sg13g2_fill_2 FILLER_0_60_578 ();
 sg13g2_decap_8 FILLER_0_60_606 ();
 sg13g2_fill_2 FILLER_0_60_613 ();
 sg13g2_decap_8 FILLER_0_60_639 ();
 sg13g2_decap_8 FILLER_0_60_646 ();
 sg13g2_decap_4 FILLER_0_60_653 ();
 sg13g2_fill_1 FILLER_0_60_666 ();
 sg13g2_fill_2 FILLER_0_60_680 ();
 sg13g2_fill_1 FILLER_0_60_697 ();
 sg13g2_fill_1 FILLER_0_60_708 ();
 sg13g2_decap_8 FILLER_0_60_742 ();
 sg13g2_decap_8 FILLER_0_60_753 ();
 sg13g2_decap_8 FILLER_0_60_760 ();
 sg13g2_decap_8 FILLER_0_60_767 ();
 sg13g2_decap_8 FILLER_0_60_774 ();
 sg13g2_decap_8 FILLER_0_60_781 ();
 sg13g2_decap_8 FILLER_0_60_788 ();
 sg13g2_fill_2 FILLER_0_60_795 ();
 sg13g2_fill_1 FILLER_0_60_797 ();
 sg13g2_fill_2 FILLER_0_60_834 ();
 sg13g2_fill_1 FILLER_0_60_836 ();
 sg13g2_fill_1 FILLER_0_60_876 ();
 sg13g2_fill_2 FILLER_0_60_881 ();
 sg13g2_fill_2 FILLER_0_60_888 ();
 sg13g2_fill_1 FILLER_0_60_890 ();
 sg13g2_fill_1 FILLER_0_60_901 ();
 sg13g2_decap_8 FILLER_0_60_905 ();
 sg13g2_decap_8 FILLER_0_60_912 ();
 sg13g2_fill_2 FILLER_0_60_919 ();
 sg13g2_fill_1 FILLER_0_60_921 ();
 sg13g2_decap_8 FILLER_0_60_937 ();
 sg13g2_decap_8 FILLER_0_60_944 ();
 sg13g2_decap_8 FILLER_0_60_951 ();
 sg13g2_fill_2 FILLER_0_60_958 ();
 sg13g2_decap_8 FILLER_0_60_971 ();
 sg13g2_fill_1 FILLER_0_60_978 ();
 sg13g2_decap_8 FILLER_0_60_984 ();
 sg13g2_decap_4 FILLER_0_60_991 ();
 sg13g2_fill_2 FILLER_0_60_999 ();
 sg13g2_fill_2 FILLER_0_60_1006 ();
 sg13g2_fill_2 FILLER_0_60_1029 ();
 sg13g2_fill_1 FILLER_0_60_1031 ();
 sg13g2_decap_8 FILLER_0_60_1046 ();
 sg13g2_decap_8 FILLER_0_60_1053 ();
 sg13g2_fill_2 FILLER_0_60_1060 ();
 sg13g2_fill_1 FILLER_0_60_1062 ();
 sg13g2_decap_8 FILLER_0_60_1078 ();
 sg13g2_decap_8 FILLER_0_60_1085 ();
 sg13g2_decap_8 FILLER_0_60_1092 ();
 sg13g2_decap_8 FILLER_0_60_1099 ();
 sg13g2_decap_4 FILLER_0_60_1106 ();
 sg13g2_decap_8 FILLER_0_60_1120 ();
 sg13g2_decap_8 FILLER_0_60_1127 ();
 sg13g2_decap_8 FILLER_0_60_1134 ();
 sg13g2_decap_8 FILLER_0_60_1141 ();
 sg13g2_decap_8 FILLER_0_60_1148 ();
 sg13g2_decap_8 FILLER_0_60_1155 ();
 sg13g2_decap_8 FILLER_0_60_1162 ();
 sg13g2_decap_8 FILLER_0_60_1169 ();
 sg13g2_decap_8 FILLER_0_60_1176 ();
 sg13g2_decap_8 FILLER_0_60_1183 ();
 sg13g2_decap_8 FILLER_0_60_1190 ();
 sg13g2_decap_8 FILLER_0_60_1197 ();
 sg13g2_decap_8 FILLER_0_60_1204 ();
 sg13g2_decap_8 FILLER_0_60_1211 ();
 sg13g2_decap_8 FILLER_0_60_1218 ();
 sg13g2_fill_2 FILLER_0_60_1225 ();
 sg13g2_fill_1 FILLER_0_60_1227 ();
 sg13g2_decap_8 FILLER_0_61_0 ();
 sg13g2_decap_8 FILLER_0_61_7 ();
 sg13g2_decap_8 FILLER_0_61_14 ();
 sg13g2_decap_8 FILLER_0_61_21 ();
 sg13g2_decap_8 FILLER_0_61_28 ();
 sg13g2_decap_4 FILLER_0_61_35 ();
 sg13g2_fill_1 FILLER_0_61_39 ();
 sg13g2_decap_8 FILLER_0_61_70 ();
 sg13g2_decap_8 FILLER_0_61_77 ();
 sg13g2_decap_8 FILLER_0_61_84 ();
 sg13g2_decap_8 FILLER_0_61_91 ();
 sg13g2_decap_8 FILLER_0_61_98 ();
 sg13g2_decap_8 FILLER_0_61_105 ();
 sg13g2_decap_8 FILLER_0_61_112 ();
 sg13g2_decap_8 FILLER_0_61_119 ();
 sg13g2_decap_4 FILLER_0_61_126 ();
 sg13g2_fill_2 FILLER_0_61_149 ();
 sg13g2_decap_4 FILLER_0_61_194 ();
 sg13g2_fill_1 FILLER_0_61_198 ();
 sg13g2_fill_1 FILLER_0_61_240 ();
 sg13g2_decap_4 FILLER_0_61_251 ();
 sg13g2_fill_2 FILLER_0_61_255 ();
 sg13g2_decap_8 FILLER_0_61_261 ();
 sg13g2_decap_4 FILLER_0_61_268 ();
 sg13g2_decap_4 FILLER_0_61_281 ();
 sg13g2_decap_8 FILLER_0_61_301 ();
 sg13g2_decap_8 FILLER_0_61_308 ();
 sg13g2_decap_8 FILLER_0_61_315 ();
 sg13g2_decap_8 FILLER_0_61_322 ();
 sg13g2_decap_8 FILLER_0_61_329 ();
 sg13g2_decap_8 FILLER_0_61_336 ();
 sg13g2_decap_8 FILLER_0_61_343 ();
 sg13g2_decap_8 FILLER_0_61_350 ();
 sg13g2_decap_8 FILLER_0_61_357 ();
 sg13g2_decap_8 FILLER_0_61_364 ();
 sg13g2_decap_4 FILLER_0_61_371 ();
 sg13g2_fill_2 FILLER_0_61_375 ();
 sg13g2_decap_8 FILLER_0_61_392 ();
 sg13g2_decap_8 FILLER_0_61_399 ();
 sg13g2_decap_8 FILLER_0_61_406 ();
 sg13g2_decap_8 FILLER_0_61_413 ();
 sg13g2_decap_4 FILLER_0_61_420 ();
 sg13g2_fill_2 FILLER_0_61_464 ();
 sg13g2_fill_1 FILLER_0_61_471 ();
 sg13g2_decap_8 FILLER_0_61_480 ();
 sg13g2_decap_4 FILLER_0_61_487 ();
 sg13g2_fill_1 FILLER_0_61_491 ();
 sg13g2_decap_8 FILLER_0_61_502 ();
 sg13g2_fill_1 FILLER_0_61_509 ();
 sg13g2_decap_4 FILLER_0_61_533 ();
 sg13g2_decap_4 FILLER_0_61_644 ();
 sg13g2_fill_1 FILLER_0_61_648 ();
 sg13g2_decap_4 FILLER_0_61_675 ();
 sg13g2_decap_8 FILLER_0_61_689 ();
 sg13g2_decap_8 FILLER_0_61_696 ();
 sg13g2_decap_8 FILLER_0_61_703 ();
 sg13g2_decap_8 FILLER_0_61_710 ();
 sg13g2_decap_8 FILLER_0_61_717 ();
 sg13g2_decap_8 FILLER_0_61_724 ();
 sg13g2_decap_8 FILLER_0_61_731 ();
 sg13g2_fill_2 FILLER_0_61_738 ();
 sg13g2_decap_8 FILLER_0_61_757 ();
 sg13g2_decap_8 FILLER_0_61_764 ();
 sg13g2_decap_8 FILLER_0_61_771 ();
 sg13g2_decap_8 FILLER_0_61_778 ();
 sg13g2_decap_8 FILLER_0_61_785 ();
 sg13g2_decap_8 FILLER_0_61_792 ();
 sg13g2_fill_1 FILLER_0_61_799 ();
 sg13g2_fill_2 FILLER_0_61_814 ();
 sg13g2_decap_8 FILLER_0_61_866 ();
 sg13g2_decap_8 FILLER_0_61_873 ();
 sg13g2_fill_1 FILLER_0_61_880 ();
 sg13g2_decap_8 FILLER_0_61_911 ();
 sg13g2_decap_4 FILLER_0_61_918 ();
 sg13g2_decap_8 FILLER_0_61_926 ();
 sg13g2_fill_2 FILLER_0_61_933 ();
 sg13g2_fill_1 FILLER_0_61_935 ();
 sg13g2_decap_8 FILLER_0_61_946 ();
 sg13g2_decap_8 FILLER_0_61_953 ();
 sg13g2_decap_8 FILLER_0_61_960 ();
 sg13g2_decap_8 FILLER_0_61_967 ();
 sg13g2_decap_8 FILLER_0_61_974 ();
 sg13g2_decap_4 FILLER_0_61_981 ();
 sg13g2_fill_2 FILLER_0_61_985 ();
 sg13g2_fill_2 FILLER_0_61_1013 ();
 sg13g2_decap_4 FILLER_0_61_1020 ();
 sg13g2_decap_4 FILLER_0_61_1050 ();
 sg13g2_fill_2 FILLER_0_61_1080 ();
 sg13g2_fill_1 FILLER_0_61_1082 ();
 sg13g2_decap_4 FILLER_0_61_1093 ();
 sg13g2_fill_1 FILLER_0_61_1097 ();
 sg13g2_decap_8 FILLER_0_61_1129 ();
 sg13g2_decap_8 FILLER_0_61_1136 ();
 sg13g2_decap_8 FILLER_0_61_1143 ();
 sg13g2_decap_8 FILLER_0_61_1150 ();
 sg13g2_decap_8 FILLER_0_61_1157 ();
 sg13g2_decap_8 FILLER_0_61_1164 ();
 sg13g2_decap_8 FILLER_0_61_1171 ();
 sg13g2_decap_8 FILLER_0_61_1178 ();
 sg13g2_decap_8 FILLER_0_61_1185 ();
 sg13g2_decap_8 FILLER_0_61_1192 ();
 sg13g2_decap_8 FILLER_0_61_1199 ();
 sg13g2_decap_8 FILLER_0_61_1206 ();
 sg13g2_decap_8 FILLER_0_61_1213 ();
 sg13g2_decap_8 FILLER_0_61_1220 ();
 sg13g2_fill_1 FILLER_0_61_1227 ();
 sg13g2_decap_8 FILLER_0_62_0 ();
 sg13g2_decap_8 FILLER_0_62_7 ();
 sg13g2_decap_8 FILLER_0_62_14 ();
 sg13g2_decap_8 FILLER_0_62_21 ();
 sg13g2_decap_8 FILLER_0_62_28 ();
 sg13g2_decap_8 FILLER_0_62_35 ();
 sg13g2_decap_8 FILLER_0_62_42 ();
 sg13g2_decap_8 FILLER_0_62_49 ();
 sg13g2_decap_8 FILLER_0_62_56 ();
 sg13g2_fill_2 FILLER_0_62_63 ();
 sg13g2_decap_8 FILLER_0_62_75 ();
 sg13g2_decap_8 FILLER_0_62_82 ();
 sg13g2_decap_8 FILLER_0_62_89 ();
 sg13g2_decap_8 FILLER_0_62_96 ();
 sg13g2_decap_8 FILLER_0_62_103 ();
 sg13g2_decap_8 FILLER_0_62_110 ();
 sg13g2_fill_2 FILLER_0_62_117 ();
 sg13g2_decap_8 FILLER_0_62_149 ();
 sg13g2_fill_2 FILLER_0_62_156 ();
 sg13g2_decap_8 FILLER_0_62_163 ();
 sg13g2_fill_2 FILLER_0_62_170 ();
 sg13g2_decap_4 FILLER_0_62_199 ();
 sg13g2_decap_8 FILLER_0_62_207 ();
 sg13g2_decap_8 FILLER_0_62_218 ();
 sg13g2_decap_8 FILLER_0_62_225 ();
 sg13g2_decap_8 FILLER_0_62_232 ();
 sg13g2_decap_4 FILLER_0_62_244 ();
 sg13g2_fill_2 FILLER_0_62_248 ();
 sg13g2_decap_4 FILLER_0_62_260 ();
 sg13g2_decap_8 FILLER_0_62_295 ();
 sg13g2_decap_8 FILLER_0_62_302 ();
 sg13g2_decap_8 FILLER_0_62_309 ();
 sg13g2_decap_8 FILLER_0_62_316 ();
 sg13g2_decap_8 FILLER_0_62_323 ();
 sg13g2_decap_8 FILLER_0_62_330 ();
 sg13g2_decap_8 FILLER_0_62_337 ();
 sg13g2_decap_8 FILLER_0_62_344 ();
 sg13g2_decap_8 FILLER_0_62_351 ();
 sg13g2_decap_4 FILLER_0_62_358 ();
 sg13g2_fill_1 FILLER_0_62_419 ();
 sg13g2_decap_8 FILLER_0_62_424 ();
 sg13g2_decap_8 FILLER_0_62_466 ();
 sg13g2_decap_8 FILLER_0_62_473 ();
 sg13g2_decap_8 FILLER_0_62_480 ();
 sg13g2_decap_8 FILLER_0_62_487 ();
 sg13g2_decap_8 FILLER_0_62_494 ();
 sg13g2_decap_8 FILLER_0_62_501 ();
 sg13g2_decap_8 FILLER_0_62_508 ();
 sg13g2_decap_8 FILLER_0_62_515 ();
 sg13g2_decap_8 FILLER_0_62_522 ();
 sg13g2_fill_1 FILLER_0_62_529 ();
 sg13g2_decap_4 FILLER_0_62_535 ();
 sg13g2_fill_2 FILLER_0_62_539 ();
 sg13g2_decap_8 FILLER_0_62_561 ();
 sg13g2_decap_8 FILLER_0_62_568 ();
 sg13g2_decap_4 FILLER_0_62_575 ();
 sg13g2_fill_2 FILLER_0_62_579 ();
 sg13g2_decap_8 FILLER_0_62_585 ();
 sg13g2_fill_2 FILLER_0_62_597 ();
 sg13g2_decap_8 FILLER_0_62_609 ();
 sg13g2_fill_2 FILLER_0_62_616 ();
 sg13g2_decap_8 FILLER_0_62_648 ();
 sg13g2_decap_8 FILLER_0_62_655 ();
 sg13g2_fill_1 FILLER_0_62_677 ();
 sg13g2_fill_2 FILLER_0_62_720 ();
 sg13g2_decap_8 FILLER_0_62_768 ();
 sg13g2_decap_8 FILLER_0_62_775 ();
 sg13g2_decap_8 FILLER_0_62_782 ();
 sg13g2_decap_8 FILLER_0_62_789 ();
 sg13g2_decap_8 FILLER_0_62_796 ();
 sg13g2_fill_1 FILLER_0_62_803 ();
 sg13g2_decap_4 FILLER_0_62_809 ();
 sg13g2_fill_1 FILLER_0_62_813 ();
 sg13g2_decap_8 FILLER_0_62_828 ();
 sg13g2_fill_1 FILLER_0_62_835 ();
 sg13g2_decap_8 FILLER_0_62_902 ();
 sg13g2_decap_4 FILLER_0_62_909 ();
 sg13g2_fill_2 FILLER_0_62_913 ();
 sg13g2_decap_8 FILLER_0_62_946 ();
 sg13g2_decap_8 FILLER_0_62_953 ();
 sg13g2_decap_4 FILLER_0_62_960 ();
 sg13g2_fill_1 FILLER_0_62_964 ();
 sg13g2_decap_8 FILLER_0_62_1022 ();
 sg13g2_fill_2 FILLER_0_62_1029 ();
 sg13g2_fill_1 FILLER_0_62_1031 ();
 sg13g2_decap_4 FILLER_0_62_1036 ();
 sg13g2_fill_2 FILLER_0_62_1040 ();
 sg13g2_decap_8 FILLER_0_62_1046 ();
 sg13g2_fill_2 FILLER_0_62_1053 ();
 sg13g2_fill_1 FILLER_0_62_1059 ();
 sg13g2_decap_8 FILLER_0_62_1101 ();
 sg13g2_fill_2 FILLER_0_62_1108 ();
 sg13g2_decap_8 FILLER_0_62_1114 ();
 sg13g2_fill_2 FILLER_0_62_1121 ();
 sg13g2_decap_8 FILLER_0_62_1127 ();
 sg13g2_decap_8 FILLER_0_62_1134 ();
 sg13g2_decap_8 FILLER_0_62_1141 ();
 sg13g2_decap_8 FILLER_0_62_1148 ();
 sg13g2_decap_8 FILLER_0_62_1155 ();
 sg13g2_decap_8 FILLER_0_62_1162 ();
 sg13g2_decap_8 FILLER_0_62_1169 ();
 sg13g2_decap_8 FILLER_0_62_1176 ();
 sg13g2_decap_8 FILLER_0_62_1183 ();
 sg13g2_decap_8 FILLER_0_62_1190 ();
 sg13g2_decap_8 FILLER_0_62_1197 ();
 sg13g2_decap_8 FILLER_0_62_1204 ();
 sg13g2_decap_8 FILLER_0_62_1211 ();
 sg13g2_decap_8 FILLER_0_62_1218 ();
 sg13g2_fill_2 FILLER_0_62_1225 ();
 sg13g2_fill_1 FILLER_0_62_1227 ();
 sg13g2_decap_8 FILLER_0_63_0 ();
 sg13g2_decap_8 FILLER_0_63_7 ();
 sg13g2_decap_8 FILLER_0_63_14 ();
 sg13g2_decap_8 FILLER_0_63_21 ();
 sg13g2_decap_8 FILLER_0_63_28 ();
 sg13g2_decap_4 FILLER_0_63_35 ();
 sg13g2_fill_2 FILLER_0_63_39 ();
 sg13g2_decap_8 FILLER_0_63_76 ();
 sg13g2_decap_8 FILLER_0_63_83 ();
 sg13g2_decap_8 FILLER_0_63_90 ();
 sg13g2_decap_8 FILLER_0_63_97 ();
 sg13g2_decap_8 FILLER_0_63_104 ();
 sg13g2_decap_4 FILLER_0_63_111 ();
 sg13g2_decap_8 FILLER_0_63_149 ();
 sg13g2_decap_8 FILLER_0_63_156 ();
 sg13g2_decap_4 FILLER_0_63_163 ();
 sg13g2_fill_1 FILLER_0_63_167 ();
 sg13g2_fill_2 FILLER_0_63_176 ();
 sg13g2_fill_1 FILLER_0_63_178 ();
 sg13g2_decap_8 FILLER_0_63_184 ();
 sg13g2_decap_4 FILLER_0_63_191 ();
 sg13g2_fill_2 FILLER_0_63_195 ();
 sg13g2_decap_8 FILLER_0_63_228 ();
 sg13g2_decap_8 FILLER_0_63_310 ();
 sg13g2_decap_8 FILLER_0_63_317 ();
 sg13g2_fill_2 FILLER_0_63_339 ();
 sg13g2_fill_1 FILLER_0_63_341 ();
 sg13g2_decap_4 FILLER_0_63_346 ();
 sg13g2_fill_1 FILLER_0_63_350 ();
 sg13g2_fill_2 FILLER_0_63_377 ();
 sg13g2_decap_4 FILLER_0_63_389 ();
 sg13g2_fill_1 FILLER_0_63_393 ();
 sg13g2_fill_2 FILLER_0_63_399 ();
 sg13g2_fill_1 FILLER_0_63_401 ();
 sg13g2_decap_8 FILLER_0_63_417 ();
 sg13g2_decap_8 FILLER_0_63_424 ();
 sg13g2_fill_2 FILLER_0_63_431 ();
 sg13g2_fill_2 FILLER_0_63_445 ();
 sg13g2_fill_1 FILLER_0_63_447 ();
 sg13g2_decap_8 FILLER_0_63_489 ();
 sg13g2_decap_4 FILLER_0_63_505 ();
 sg13g2_decap_8 FILLER_0_63_519 ();
 sg13g2_decap_8 FILLER_0_63_526 ();
 sg13g2_decap_8 FILLER_0_63_533 ();
 sg13g2_fill_2 FILLER_0_63_540 ();
 sg13g2_fill_1 FILLER_0_63_607 ();
 sg13g2_fill_1 FILLER_0_63_618 ();
 sg13g2_fill_1 FILLER_0_63_624 ();
 sg13g2_decap_8 FILLER_0_63_635 ();
 sg13g2_fill_1 FILLER_0_63_642 ();
 sg13g2_fill_2 FILLER_0_63_673 ();
 sg13g2_fill_2 FILLER_0_63_701 ();
 sg13g2_fill_1 FILLER_0_63_738 ();
 sg13g2_decap_4 FILLER_0_63_752 ();
 sg13g2_decap_4 FILLER_0_63_787 ();
 sg13g2_fill_2 FILLER_0_63_799 ();
 sg13g2_fill_1 FILLER_0_63_801 ();
 sg13g2_fill_2 FILLER_0_63_828 ();
 sg13g2_fill_1 FILLER_0_63_830 ();
 sg13g2_fill_2 FILLER_0_63_872 ();
 sg13g2_fill_1 FILLER_0_63_874 ();
 sg13g2_fill_2 FILLER_0_63_982 ();
 sg13g2_fill_1 FILLER_0_63_984 ();
 sg13g2_fill_2 FILLER_0_63_995 ();
 sg13g2_fill_1 FILLER_0_63_997 ();
 sg13g2_fill_1 FILLER_0_63_1059 ();
 sg13g2_fill_2 FILLER_0_63_1105 ();
 sg13g2_decap_8 FILLER_0_63_1143 ();
 sg13g2_decap_8 FILLER_0_63_1150 ();
 sg13g2_decap_8 FILLER_0_63_1157 ();
 sg13g2_decap_8 FILLER_0_63_1164 ();
 sg13g2_decap_8 FILLER_0_63_1171 ();
 sg13g2_decap_8 FILLER_0_63_1178 ();
 sg13g2_decap_8 FILLER_0_63_1185 ();
 sg13g2_decap_8 FILLER_0_63_1192 ();
 sg13g2_decap_8 FILLER_0_63_1199 ();
 sg13g2_decap_8 FILLER_0_63_1206 ();
 sg13g2_decap_8 FILLER_0_63_1213 ();
 sg13g2_decap_8 FILLER_0_63_1220 ();
 sg13g2_fill_1 FILLER_0_63_1227 ();
 sg13g2_decap_8 FILLER_0_64_0 ();
 sg13g2_decap_8 FILLER_0_64_7 ();
 sg13g2_decap_8 FILLER_0_64_14 ();
 sg13g2_decap_8 FILLER_0_64_21 ();
 sg13g2_decap_8 FILLER_0_64_28 ();
 sg13g2_decap_8 FILLER_0_64_35 ();
 sg13g2_decap_4 FILLER_0_64_47 ();
 sg13g2_fill_1 FILLER_0_64_51 ();
 sg13g2_decap_8 FILLER_0_64_72 ();
 sg13g2_decap_8 FILLER_0_64_79 ();
 sg13g2_decap_8 FILLER_0_64_86 ();
 sg13g2_decap_8 FILLER_0_64_93 ();
 sg13g2_decap_8 FILLER_0_64_100 ();
 sg13g2_decap_8 FILLER_0_64_107 ();
 sg13g2_decap_8 FILLER_0_64_114 ();
 sg13g2_fill_1 FILLER_0_64_121 ();
 sg13g2_fill_1 FILLER_0_64_140 ();
 sg13g2_fill_2 FILLER_0_64_151 ();
 sg13g2_fill_2 FILLER_0_64_157 ();
 sg13g2_fill_2 FILLER_0_64_185 ();
 sg13g2_fill_1 FILLER_0_64_197 ();
 sg13g2_fill_1 FILLER_0_64_208 ();
 sg13g2_decap_8 FILLER_0_64_213 ();
 sg13g2_fill_2 FILLER_0_64_220 ();
 sg13g2_fill_1 FILLER_0_64_222 ();
 sg13g2_fill_1 FILLER_0_64_267 ();
 sg13g2_fill_2 FILLER_0_64_277 ();
 sg13g2_decap_8 FILLER_0_64_345 ();
 sg13g2_decap_4 FILLER_0_64_352 ();
 sg13g2_fill_1 FILLER_0_64_356 ();
 sg13g2_decap_4 FILLER_0_64_361 ();
 sg13g2_fill_1 FILLER_0_64_365 ();
 sg13g2_fill_1 FILLER_0_64_429 ();
 sg13g2_fill_2 FILLER_0_64_435 ();
 sg13g2_fill_2 FILLER_0_64_447 ();
 sg13g2_fill_1 FILLER_0_64_449 ();
 sg13g2_fill_1 FILLER_0_64_465 ();
 sg13g2_fill_1 FILLER_0_64_492 ();
 sg13g2_fill_1 FILLER_0_64_524 ();
 sg13g2_decap_8 FILLER_0_64_529 ();
 sg13g2_fill_2 FILLER_0_64_536 ();
 sg13g2_fill_1 FILLER_0_64_538 ();
 sg13g2_decap_8 FILLER_0_64_565 ();
 sg13g2_decap_8 FILLER_0_64_572 ();
 sg13g2_decap_4 FILLER_0_64_579 ();
 sg13g2_fill_1 FILLER_0_64_583 ();
 sg13g2_fill_2 FILLER_0_64_610 ();
 sg13g2_decap_4 FILLER_0_64_638 ();
 sg13g2_decap_4 FILLER_0_64_647 ();
 sg13g2_decap_4 FILLER_0_64_665 ();
 sg13g2_fill_2 FILLER_0_64_679 ();
 sg13g2_fill_1 FILLER_0_64_681 ();
 sg13g2_fill_1 FILLER_0_64_748 ();
 sg13g2_decap_8 FILLER_0_64_759 ();
 sg13g2_fill_1 FILLER_0_64_766 ();
 sg13g2_decap_8 FILLER_0_64_771 ();
 sg13g2_decap_8 FILLER_0_64_778 ();
 sg13g2_decap_8 FILLER_0_64_785 ();
 sg13g2_decap_8 FILLER_0_64_792 ();
 sg13g2_decap_8 FILLER_0_64_799 ();
 sg13g2_fill_2 FILLER_0_64_806 ();
 sg13g2_decap_4 FILLER_0_64_812 ();
 sg13g2_decap_8 FILLER_0_64_826 ();
 sg13g2_decap_4 FILLER_0_64_833 ();
 sg13g2_fill_2 FILLER_0_64_837 ();
 sg13g2_decap_8 FILLER_0_64_843 ();
 sg13g2_fill_2 FILLER_0_64_850 ();
 sg13g2_fill_1 FILLER_0_64_852 ();
 sg13g2_fill_1 FILLER_0_64_858 ();
 sg13g2_decap_8 FILLER_0_64_869 ();
 sg13g2_fill_2 FILLER_0_64_913 ();
 sg13g2_decap_8 FILLER_0_64_939 ();
 sg13g2_decap_8 FILLER_0_64_946 ();
 sg13g2_decap_8 FILLER_0_64_953 ();
 sg13g2_decap_8 FILLER_0_64_964 ();
 sg13g2_fill_2 FILLER_0_64_971 ();
 sg13g2_fill_1 FILLER_0_64_973 ();
 sg13g2_decap_8 FILLER_0_64_988 ();
 sg13g2_decap_8 FILLER_0_64_995 ();
 sg13g2_decap_4 FILLER_0_64_1006 ();
 sg13g2_fill_1 FILLER_0_64_1010 ();
 sg13g2_decap_8 FILLER_0_64_1019 ();
 sg13g2_decap_8 FILLER_0_64_1026 ();
 sg13g2_decap_8 FILLER_0_64_1033 ();
 sg13g2_decap_8 FILLER_0_64_1040 ();
 sg13g2_decap_8 FILLER_0_64_1047 ();
 sg13g2_decap_8 FILLER_0_64_1054 ();
 sg13g2_decap_8 FILLER_0_64_1061 ();
 sg13g2_decap_8 FILLER_0_64_1068 ();
 sg13g2_fill_1 FILLER_0_64_1075 ();
 sg13g2_fill_2 FILLER_0_64_1084 ();
 sg13g2_fill_1 FILLER_0_64_1086 ();
 sg13g2_fill_2 FILLER_0_64_1104 ();
 sg13g2_decap_8 FILLER_0_64_1111 ();
 sg13g2_decap_8 FILLER_0_64_1118 ();
 sg13g2_decap_8 FILLER_0_64_1125 ();
 sg13g2_decap_8 FILLER_0_64_1132 ();
 sg13g2_decap_8 FILLER_0_64_1139 ();
 sg13g2_decap_8 FILLER_0_64_1146 ();
 sg13g2_decap_8 FILLER_0_64_1153 ();
 sg13g2_decap_8 FILLER_0_64_1160 ();
 sg13g2_decap_8 FILLER_0_64_1167 ();
 sg13g2_decap_8 FILLER_0_64_1174 ();
 sg13g2_decap_8 FILLER_0_64_1181 ();
 sg13g2_decap_8 FILLER_0_64_1188 ();
 sg13g2_decap_8 FILLER_0_64_1195 ();
 sg13g2_decap_8 FILLER_0_64_1202 ();
 sg13g2_decap_8 FILLER_0_64_1209 ();
 sg13g2_decap_8 FILLER_0_64_1216 ();
 sg13g2_decap_4 FILLER_0_64_1223 ();
 sg13g2_fill_1 FILLER_0_64_1227 ();
 sg13g2_decap_8 FILLER_0_65_0 ();
 sg13g2_decap_8 FILLER_0_65_7 ();
 sg13g2_decap_8 FILLER_0_65_14 ();
 sg13g2_decap_8 FILLER_0_65_21 ();
 sg13g2_decap_8 FILLER_0_65_28 ();
 sg13g2_fill_2 FILLER_0_65_35 ();
 sg13g2_fill_1 FILLER_0_65_37 ();
 sg13g2_fill_2 FILLER_0_65_68 ();
 sg13g2_fill_1 FILLER_0_65_70 ();
 sg13g2_fill_2 FILLER_0_65_112 ();
 sg13g2_fill_2 FILLER_0_65_118 ();
 sg13g2_fill_1 FILLER_0_65_120 ();
 sg13g2_fill_1 FILLER_0_65_188 ();
 sg13g2_decap_8 FILLER_0_65_220 ();
 sg13g2_decap_8 FILLER_0_65_227 ();
 sg13g2_decap_4 FILLER_0_65_234 ();
 sg13g2_fill_2 FILLER_0_65_243 ();
 sg13g2_fill_1 FILLER_0_65_245 ();
 sg13g2_decap_8 FILLER_0_65_268 ();
 sg13g2_decap_4 FILLER_0_65_275 ();
 sg13g2_fill_2 FILLER_0_65_279 ();
 sg13g2_decap_8 FILLER_0_65_291 ();
 sg13g2_fill_1 FILLER_0_65_308 ();
 sg13g2_fill_1 FILLER_0_65_340 ();
 sg13g2_fill_2 FILLER_0_65_367 ();
 sg13g2_fill_2 FILLER_0_65_395 ();
 sg13g2_fill_1 FILLER_0_65_397 ();
 sg13g2_fill_1 FILLER_0_65_501 ();
 sg13g2_fill_2 FILLER_0_65_506 ();
 sg13g2_decap_4 FILLER_0_65_534 ();
 sg13g2_decap_4 FILLER_0_65_543 ();
 sg13g2_decap_4 FILLER_0_65_551 ();
 sg13g2_decap_8 FILLER_0_65_565 ();
 sg13g2_fill_2 FILLER_0_65_572 ();
 sg13g2_fill_1 FILLER_0_65_574 ();
 sg13g2_fill_1 FILLER_0_65_606 ();
 sg13g2_fill_1 FILLER_0_65_620 ();
 sg13g2_decap_8 FILLER_0_65_625 ();
 sg13g2_decap_8 FILLER_0_65_632 ();
 sg13g2_decap_4 FILLER_0_65_639 ();
 sg13g2_fill_1 FILLER_0_65_643 ();
 sg13g2_fill_2 FILLER_0_65_670 ();
 sg13g2_decap_8 FILLER_0_65_680 ();
 sg13g2_decap_8 FILLER_0_65_687 ();
 sg13g2_decap_8 FILLER_0_65_694 ();
 sg13g2_decap_8 FILLER_0_65_701 ();
 sg13g2_decap_8 FILLER_0_65_708 ();
 sg13g2_decap_8 FILLER_0_65_715 ();
 sg13g2_decap_8 FILLER_0_65_722 ();
 sg13g2_decap_8 FILLER_0_65_729 ();
 sg13g2_decap_8 FILLER_0_65_736 ();
 sg13g2_fill_2 FILLER_0_65_743 ();
 sg13g2_fill_1 FILLER_0_65_745 ();
 sg13g2_fill_2 FILLER_0_65_750 ();
 sg13g2_decap_8 FILLER_0_65_762 ();
 sg13g2_fill_2 FILLER_0_65_769 ();
 sg13g2_decap_8 FILLER_0_65_797 ();
 sg13g2_fill_1 FILLER_0_65_804 ();
 sg13g2_decap_8 FILLER_0_65_836 ();
 sg13g2_fill_2 FILLER_0_65_843 ();
 sg13g2_decap_8 FILLER_0_65_849 ();
 sg13g2_decap_8 FILLER_0_65_856 ();
 sg13g2_fill_1 FILLER_0_65_863 ();
 sg13g2_decap_4 FILLER_0_65_874 ();
 sg13g2_fill_2 FILLER_0_65_878 ();
 sg13g2_fill_2 FILLER_0_65_885 ();
 sg13g2_decap_8 FILLER_0_65_901 ();
 sg13g2_decap_4 FILLER_0_65_908 ();
 sg13g2_fill_1 FILLER_0_65_912 ();
 sg13g2_decap_8 FILLER_0_65_954 ();
 sg13g2_decap_8 FILLER_0_65_961 ();
 sg13g2_decap_8 FILLER_0_65_1009 ();
 sg13g2_decap_8 FILLER_0_65_1016 ();
 sg13g2_decap_8 FILLER_0_65_1023 ();
 sg13g2_decap_8 FILLER_0_65_1030 ();
 sg13g2_decap_8 FILLER_0_65_1037 ();
 sg13g2_decap_8 FILLER_0_65_1044 ();
 sg13g2_decap_8 FILLER_0_65_1051 ();
 sg13g2_decap_8 FILLER_0_65_1058 ();
 sg13g2_decap_8 FILLER_0_65_1065 ();
 sg13g2_decap_8 FILLER_0_65_1072 ();
 sg13g2_decap_8 FILLER_0_65_1079 ();
 sg13g2_decap_4 FILLER_0_65_1086 ();
 sg13g2_fill_1 FILLER_0_65_1090 ();
 sg13g2_decap_8 FILLER_0_65_1104 ();
 sg13g2_decap_8 FILLER_0_65_1111 ();
 sg13g2_decap_8 FILLER_0_65_1118 ();
 sg13g2_decap_8 FILLER_0_65_1125 ();
 sg13g2_decap_8 FILLER_0_65_1132 ();
 sg13g2_decap_8 FILLER_0_65_1139 ();
 sg13g2_decap_8 FILLER_0_65_1146 ();
 sg13g2_decap_8 FILLER_0_65_1153 ();
 sg13g2_decap_8 FILLER_0_65_1160 ();
 sg13g2_decap_8 FILLER_0_65_1167 ();
 sg13g2_decap_8 FILLER_0_65_1174 ();
 sg13g2_decap_8 FILLER_0_65_1181 ();
 sg13g2_decap_8 FILLER_0_65_1188 ();
 sg13g2_decap_8 FILLER_0_65_1195 ();
 sg13g2_decap_8 FILLER_0_65_1202 ();
 sg13g2_decap_8 FILLER_0_65_1209 ();
 sg13g2_decap_8 FILLER_0_65_1216 ();
 sg13g2_decap_4 FILLER_0_65_1223 ();
 sg13g2_fill_1 FILLER_0_65_1227 ();
 sg13g2_decap_8 FILLER_0_66_0 ();
 sg13g2_decap_8 FILLER_0_66_7 ();
 sg13g2_decap_8 FILLER_0_66_14 ();
 sg13g2_decap_8 FILLER_0_66_21 ();
 sg13g2_decap_8 FILLER_0_66_28 ();
 sg13g2_fill_2 FILLER_0_66_35 ();
 sg13g2_fill_1 FILLER_0_66_37 ();
 sg13g2_decap_8 FILLER_0_66_68 ();
 sg13g2_decap_4 FILLER_0_66_75 ();
 sg13g2_fill_1 FILLER_0_66_79 ();
 sg13g2_fill_2 FILLER_0_66_150 ();
 sg13g2_decap_8 FILLER_0_66_185 ();
 sg13g2_decap_8 FILLER_0_66_192 ();
 sg13g2_decap_4 FILLER_0_66_199 ();
 sg13g2_decap_8 FILLER_0_66_207 ();
 sg13g2_decap_8 FILLER_0_66_214 ();
 sg13g2_decap_8 FILLER_0_66_221 ();
 sg13g2_decap_8 FILLER_0_66_228 ();
 sg13g2_decap_8 FILLER_0_66_235 ();
 sg13g2_decap_8 FILLER_0_66_242 ();
 sg13g2_decap_4 FILLER_0_66_249 ();
 sg13g2_fill_2 FILLER_0_66_253 ();
 sg13g2_fill_2 FILLER_0_66_259 ();
 sg13g2_decap_8 FILLER_0_66_291 ();
 sg13g2_decap_8 FILLER_0_66_298 ();
 sg13g2_decap_4 FILLER_0_66_305 ();
 sg13g2_fill_1 FILLER_0_66_309 ();
 sg13g2_decap_4 FILLER_0_66_344 ();
 sg13g2_fill_1 FILLER_0_66_352 ();
 sg13g2_decap_8 FILLER_0_66_392 ();
 sg13g2_fill_2 FILLER_0_66_399 ();
 sg13g2_fill_1 FILLER_0_66_401 ();
 sg13g2_fill_1 FILLER_0_66_407 ();
 sg13g2_decap_4 FILLER_0_66_456 ();
 sg13g2_fill_2 FILLER_0_66_460 ();
 sg13g2_fill_1 FILLER_0_66_478 ();
 sg13g2_fill_1 FILLER_0_66_483 ();
 sg13g2_fill_1 FILLER_0_66_504 ();
 sg13g2_decap_8 FILLER_0_66_535 ();
 sg13g2_decap_8 FILLER_0_66_542 ();
 sg13g2_decap_8 FILLER_0_66_549 ();
 sg13g2_decap_4 FILLER_0_66_556 ();
 sg13g2_fill_1 FILLER_0_66_560 ();
 sg13g2_decap_8 FILLER_0_66_602 ();
 sg13g2_decap_8 FILLER_0_66_609 ();
 sg13g2_decap_8 FILLER_0_66_616 ();
 sg13g2_decap_8 FILLER_0_66_623 ();
 sg13g2_decap_8 FILLER_0_66_630 ();
 sg13g2_decap_8 FILLER_0_66_637 ();
 sg13g2_decap_4 FILLER_0_66_644 ();
 sg13g2_fill_1 FILLER_0_66_648 ();
 sg13g2_decap_8 FILLER_0_66_663 ();
 sg13g2_decap_8 FILLER_0_66_670 ();
 sg13g2_decap_8 FILLER_0_66_677 ();
 sg13g2_fill_2 FILLER_0_66_684 ();
 sg13g2_decap_8 FILLER_0_66_703 ();
 sg13g2_decap_8 FILLER_0_66_710 ();
 sg13g2_fill_1 FILLER_0_66_717 ();
 sg13g2_decap_8 FILLER_0_66_723 ();
 sg13g2_fill_2 FILLER_0_66_730 ();
 sg13g2_fill_2 FILLER_0_66_773 ();
 sg13g2_fill_1 FILLER_0_66_775 ();
 sg13g2_decap_8 FILLER_0_66_802 ();
 sg13g2_fill_1 FILLER_0_66_809 ();
 sg13g2_fill_2 FILLER_0_66_840 ();
 sg13g2_decap_8 FILLER_0_66_904 ();
 sg13g2_decap_8 FILLER_0_66_911 ();
 sg13g2_decap_8 FILLER_0_66_918 ();
 sg13g2_fill_2 FILLER_0_66_961 ();
 sg13g2_fill_1 FILLER_0_66_963 ();
 sg13g2_fill_1 FILLER_0_66_988 ();
 sg13g2_decap_8 FILLER_0_66_993 ();
 sg13g2_decap_8 FILLER_0_66_1000 ();
 sg13g2_decap_8 FILLER_0_66_1007 ();
 sg13g2_decap_8 FILLER_0_66_1014 ();
 sg13g2_decap_8 FILLER_0_66_1021 ();
 sg13g2_decap_8 FILLER_0_66_1028 ();
 sg13g2_decap_8 FILLER_0_66_1035 ();
 sg13g2_decap_8 FILLER_0_66_1042 ();
 sg13g2_decap_8 FILLER_0_66_1049 ();
 sg13g2_decap_8 FILLER_0_66_1056 ();
 sg13g2_decap_8 FILLER_0_66_1063 ();
 sg13g2_decap_8 FILLER_0_66_1070 ();
 sg13g2_decap_8 FILLER_0_66_1077 ();
 sg13g2_decap_8 FILLER_0_66_1084 ();
 sg13g2_decap_8 FILLER_0_66_1091 ();
 sg13g2_decap_8 FILLER_0_66_1098 ();
 sg13g2_decap_8 FILLER_0_66_1105 ();
 sg13g2_decap_8 FILLER_0_66_1112 ();
 sg13g2_decap_8 FILLER_0_66_1119 ();
 sg13g2_decap_8 FILLER_0_66_1126 ();
 sg13g2_decap_8 FILLER_0_66_1133 ();
 sg13g2_decap_8 FILLER_0_66_1140 ();
 sg13g2_decap_8 FILLER_0_66_1147 ();
 sg13g2_decap_8 FILLER_0_66_1154 ();
 sg13g2_decap_8 FILLER_0_66_1161 ();
 sg13g2_decap_8 FILLER_0_66_1168 ();
 sg13g2_decap_8 FILLER_0_66_1175 ();
 sg13g2_decap_8 FILLER_0_66_1182 ();
 sg13g2_decap_8 FILLER_0_66_1189 ();
 sg13g2_decap_8 FILLER_0_66_1196 ();
 sg13g2_decap_8 FILLER_0_66_1203 ();
 sg13g2_decap_8 FILLER_0_66_1210 ();
 sg13g2_decap_8 FILLER_0_66_1217 ();
 sg13g2_decap_4 FILLER_0_66_1224 ();
 sg13g2_decap_8 FILLER_0_67_0 ();
 sg13g2_decap_8 FILLER_0_67_7 ();
 sg13g2_decap_8 FILLER_0_67_14 ();
 sg13g2_decap_8 FILLER_0_67_21 ();
 sg13g2_decap_8 FILLER_0_67_28 ();
 sg13g2_fill_1 FILLER_0_67_35 ();
 sg13g2_fill_2 FILLER_0_67_73 ();
 sg13g2_fill_1 FILLER_0_67_75 ();
 sg13g2_fill_2 FILLER_0_67_120 ();
 sg13g2_decap_8 FILLER_0_67_136 ();
 sg13g2_decap_8 FILLER_0_67_143 ();
 sg13g2_fill_2 FILLER_0_67_150 ();
 sg13g2_fill_1 FILLER_0_67_152 ();
 sg13g2_decap_8 FILLER_0_67_184 ();
 sg13g2_decap_8 FILLER_0_67_191 ();
 sg13g2_fill_2 FILLER_0_67_198 ();
 sg13g2_decap_4 FILLER_0_67_215 ();
 sg13g2_fill_1 FILLER_0_67_219 ();
 sg13g2_decap_8 FILLER_0_67_265 ();
 sg13g2_decap_8 FILLER_0_67_272 ();
 sg13g2_decap_8 FILLER_0_67_279 ();
 sg13g2_decap_8 FILLER_0_67_286 ();
 sg13g2_decap_8 FILLER_0_67_293 ();
 sg13g2_decap_8 FILLER_0_67_300 ();
 sg13g2_decap_8 FILLER_0_67_307 ();
 sg13g2_fill_2 FILLER_0_67_314 ();
 sg13g2_fill_1 FILLER_0_67_316 ();
 sg13g2_fill_1 FILLER_0_67_322 ();
 sg13g2_fill_2 FILLER_0_67_344 ();
 sg13g2_fill_2 FILLER_0_67_351 ();
 sg13g2_fill_1 FILLER_0_67_353 ();
 sg13g2_fill_2 FILLER_0_67_364 ();
 sg13g2_decap_8 FILLER_0_67_376 ();
 sg13g2_decap_8 FILLER_0_67_383 ();
 sg13g2_decap_8 FILLER_0_67_390 ();
 sg13g2_decap_8 FILLER_0_67_397 ();
 sg13g2_decap_8 FILLER_0_67_404 ();
 sg13g2_decap_8 FILLER_0_67_415 ();
 sg13g2_decap_8 FILLER_0_67_422 ();
 sg13g2_decap_4 FILLER_0_67_429 ();
 sg13g2_fill_2 FILLER_0_67_433 ();
 sg13g2_decap_8 FILLER_0_67_450 ();
 sg13g2_decap_8 FILLER_0_67_457 ();
 sg13g2_fill_2 FILLER_0_67_464 ();
 sg13g2_decap_8 FILLER_0_67_492 ();
 sg13g2_decap_8 FILLER_0_67_499 ();
 sg13g2_fill_2 FILLER_0_67_506 ();
 sg13g2_fill_1 FILLER_0_67_508 ();
 sg13g2_fill_1 FILLER_0_67_524 ();
 sg13g2_decap_8 FILLER_0_67_530 ();
 sg13g2_decap_8 FILLER_0_67_537 ();
 sg13g2_fill_2 FILLER_0_67_544 ();
 sg13g2_fill_1 FILLER_0_67_546 ();
 sg13g2_decap_4 FILLER_0_67_550 ();
 sg13g2_fill_2 FILLER_0_67_554 ();
 sg13g2_decap_8 FILLER_0_67_592 ();
 sg13g2_decap_8 FILLER_0_67_599 ();
 sg13g2_fill_2 FILLER_0_67_606 ();
 sg13g2_fill_1 FILLER_0_67_608 ();
 sg13g2_decap_4 FILLER_0_67_623 ();
 sg13g2_fill_2 FILLER_0_67_627 ();
 sg13g2_fill_2 FILLER_0_67_686 ();
 sg13g2_fill_1 FILLER_0_67_688 ();
 sg13g2_fill_2 FILLER_0_67_723 ();
 sg13g2_fill_1 FILLER_0_67_725 ();
 sg13g2_decap_4 FILLER_0_67_736 ();
 sg13g2_fill_1 FILLER_0_67_740 ();
 sg13g2_fill_2 FILLER_0_67_745 ();
 sg13g2_fill_1 FILLER_0_67_788 ();
 sg13g2_decap_8 FILLER_0_67_804 ();
 sg13g2_decap_8 FILLER_0_67_830 ();
 sg13g2_decap_4 FILLER_0_67_837 ();
 sg13g2_fill_1 FILLER_0_67_841 ();
 sg13g2_decap_8 FILLER_0_67_868 ();
 sg13g2_decap_4 FILLER_0_67_875 ();
 sg13g2_fill_2 FILLER_0_67_879 ();
 sg13g2_fill_2 FILLER_0_67_900 ();
 sg13g2_fill_2 FILLER_0_67_959 ();
 sg13g2_decap_8 FILLER_0_67_992 ();
 sg13g2_decap_8 FILLER_0_67_999 ();
 sg13g2_decap_8 FILLER_0_67_1006 ();
 sg13g2_decap_8 FILLER_0_67_1013 ();
 sg13g2_decap_8 FILLER_0_67_1020 ();
 sg13g2_decap_8 FILLER_0_67_1027 ();
 sg13g2_decap_8 FILLER_0_67_1034 ();
 sg13g2_decap_8 FILLER_0_67_1041 ();
 sg13g2_decap_8 FILLER_0_67_1048 ();
 sg13g2_decap_8 FILLER_0_67_1055 ();
 sg13g2_decap_8 FILLER_0_67_1062 ();
 sg13g2_decap_8 FILLER_0_67_1069 ();
 sg13g2_decap_8 FILLER_0_67_1076 ();
 sg13g2_decap_8 FILLER_0_67_1083 ();
 sg13g2_decap_8 FILLER_0_67_1090 ();
 sg13g2_decap_8 FILLER_0_67_1097 ();
 sg13g2_decap_8 FILLER_0_67_1104 ();
 sg13g2_decap_8 FILLER_0_67_1111 ();
 sg13g2_decap_8 FILLER_0_67_1118 ();
 sg13g2_decap_8 FILLER_0_67_1125 ();
 sg13g2_decap_8 FILLER_0_67_1132 ();
 sg13g2_decap_8 FILLER_0_67_1139 ();
 sg13g2_decap_8 FILLER_0_67_1146 ();
 sg13g2_decap_8 FILLER_0_67_1153 ();
 sg13g2_decap_8 FILLER_0_67_1160 ();
 sg13g2_decap_8 FILLER_0_67_1167 ();
 sg13g2_decap_8 FILLER_0_67_1174 ();
 sg13g2_decap_8 FILLER_0_67_1181 ();
 sg13g2_decap_8 FILLER_0_67_1188 ();
 sg13g2_decap_8 FILLER_0_67_1195 ();
 sg13g2_decap_8 FILLER_0_67_1202 ();
 sg13g2_decap_8 FILLER_0_67_1209 ();
 sg13g2_decap_8 FILLER_0_67_1216 ();
 sg13g2_decap_4 FILLER_0_67_1223 ();
 sg13g2_fill_1 FILLER_0_67_1227 ();
 sg13g2_decap_8 FILLER_0_68_0 ();
 sg13g2_decap_8 FILLER_0_68_7 ();
 sg13g2_decap_8 FILLER_0_68_14 ();
 sg13g2_decap_8 FILLER_0_68_21 ();
 sg13g2_decap_8 FILLER_0_68_28 ();
 sg13g2_decap_8 FILLER_0_68_35 ();
 sg13g2_fill_1 FILLER_0_68_42 ();
 sg13g2_decap_8 FILLER_0_68_74 ();
 sg13g2_decap_4 FILLER_0_68_81 ();
 sg13g2_fill_1 FILLER_0_68_85 ();
 sg13g2_decap_8 FILLER_0_68_101 ();
 sg13g2_decap_8 FILLER_0_68_108 ();
 sg13g2_decap_8 FILLER_0_68_115 ();
 sg13g2_decap_8 FILLER_0_68_122 ();
 sg13g2_decap_8 FILLER_0_68_129 ();
 sg13g2_decap_8 FILLER_0_68_136 ();
 sg13g2_decap_8 FILLER_0_68_143 ();
 sg13g2_decap_8 FILLER_0_68_150 ();
 sg13g2_fill_2 FILLER_0_68_157 ();
 sg13g2_fill_2 FILLER_0_68_163 ();
 sg13g2_fill_1 FILLER_0_68_165 ();
 sg13g2_decap_4 FILLER_0_68_171 ();
 sg13g2_fill_1 FILLER_0_68_175 ();
 sg13g2_decap_8 FILLER_0_68_186 ();
 sg13g2_decap_4 FILLER_0_68_234 ();
 sg13g2_fill_1 FILLER_0_68_238 ();
 sg13g2_decap_8 FILLER_0_68_254 ();
 sg13g2_decap_8 FILLER_0_68_261 ();
 sg13g2_decap_8 FILLER_0_68_268 ();
 sg13g2_decap_8 FILLER_0_68_275 ();
 sg13g2_decap_8 FILLER_0_68_282 ();
 sg13g2_decap_8 FILLER_0_68_289 ();
 sg13g2_decap_8 FILLER_0_68_296 ();
 sg13g2_decap_8 FILLER_0_68_303 ();
 sg13g2_decap_8 FILLER_0_68_310 ();
 sg13g2_fill_2 FILLER_0_68_317 ();
 sg13g2_decap_8 FILLER_0_68_332 ();
 sg13g2_decap_8 FILLER_0_68_339 ();
 sg13g2_decap_8 FILLER_0_68_346 ();
 sg13g2_decap_8 FILLER_0_68_353 ();
 sg13g2_decap_8 FILLER_0_68_360 ();
 sg13g2_decap_8 FILLER_0_68_367 ();
 sg13g2_decap_8 FILLER_0_68_374 ();
 sg13g2_decap_8 FILLER_0_68_381 ();
 sg13g2_decap_8 FILLER_0_68_388 ();
 sg13g2_decap_8 FILLER_0_68_395 ();
 sg13g2_decap_8 FILLER_0_68_402 ();
 sg13g2_decap_8 FILLER_0_68_409 ();
 sg13g2_decap_8 FILLER_0_68_416 ();
 sg13g2_decap_8 FILLER_0_68_423 ();
 sg13g2_decap_8 FILLER_0_68_430 ();
 sg13g2_fill_2 FILLER_0_68_437 ();
 sg13g2_fill_1 FILLER_0_68_439 ();
 sg13g2_decap_8 FILLER_0_68_455 ();
 sg13g2_decap_4 FILLER_0_68_467 ();
 sg13g2_decap_8 FILLER_0_68_485 ();
 sg13g2_decap_8 FILLER_0_68_492 ();
 sg13g2_decap_8 FILLER_0_68_499 ();
 sg13g2_fill_1 FILLER_0_68_526 ();
 sg13g2_fill_2 FILLER_0_68_561 ();
 sg13g2_fill_1 FILLER_0_68_563 ();
 sg13g2_fill_1 FILLER_0_68_574 ();
 sg13g2_decap_8 FILLER_0_68_579 ();
 sg13g2_fill_1 FILLER_0_68_586 ();
 sg13g2_decap_4 FILLER_0_68_592 ();
 sg13g2_fill_1 FILLER_0_68_596 ();
 sg13g2_decap_8 FILLER_0_68_659 ();
 sg13g2_fill_1 FILLER_0_68_666 ();
 sg13g2_fill_1 FILLER_0_68_671 ();
 sg13g2_fill_2 FILLER_0_68_698 ();
 sg13g2_fill_2 FILLER_0_68_731 ();
 sg13g2_fill_1 FILLER_0_68_733 ();
 sg13g2_fill_1 FILLER_0_68_754 ();
 sg13g2_fill_2 FILLER_0_68_759 ();
 sg13g2_decap_4 FILLER_0_68_766 ();
 sg13g2_decap_4 FILLER_0_68_774 ();
 sg13g2_fill_1 FILLER_0_68_778 ();
 sg13g2_fill_1 FILLER_0_68_783 ();
 sg13g2_decap_8 FILLER_0_68_824 ();
 sg13g2_fill_2 FILLER_0_68_831 ();
 sg13g2_fill_1 FILLER_0_68_833 ();
 sg13g2_decap_4 FILLER_0_68_845 ();
 sg13g2_fill_2 FILLER_0_68_849 ();
 sg13g2_decap_8 FILLER_0_68_870 ();
 sg13g2_decap_8 FILLER_0_68_877 ();
 sg13g2_fill_1 FILLER_0_68_943 ();
 sg13g2_fill_1 FILLER_0_68_954 ();
 sg13g2_decap_8 FILLER_0_68_986 ();
 sg13g2_decap_4 FILLER_0_68_993 ();
 sg13g2_fill_2 FILLER_0_68_997 ();
 sg13g2_fill_2 FILLER_0_68_1010 ();
 sg13g2_decap_8 FILLER_0_68_1020 ();
 sg13g2_decap_8 FILLER_0_68_1027 ();
 sg13g2_decap_8 FILLER_0_68_1034 ();
 sg13g2_decap_8 FILLER_0_68_1041 ();
 sg13g2_decap_8 FILLER_0_68_1048 ();
 sg13g2_decap_8 FILLER_0_68_1055 ();
 sg13g2_decap_8 FILLER_0_68_1062 ();
 sg13g2_decap_8 FILLER_0_68_1069 ();
 sg13g2_decap_8 FILLER_0_68_1076 ();
 sg13g2_decap_8 FILLER_0_68_1083 ();
 sg13g2_decap_8 FILLER_0_68_1090 ();
 sg13g2_decap_8 FILLER_0_68_1097 ();
 sg13g2_decap_8 FILLER_0_68_1104 ();
 sg13g2_decap_8 FILLER_0_68_1111 ();
 sg13g2_decap_8 FILLER_0_68_1118 ();
 sg13g2_decap_8 FILLER_0_68_1125 ();
 sg13g2_decap_8 FILLER_0_68_1132 ();
 sg13g2_decap_8 FILLER_0_68_1139 ();
 sg13g2_decap_8 FILLER_0_68_1146 ();
 sg13g2_decap_8 FILLER_0_68_1153 ();
 sg13g2_decap_8 FILLER_0_68_1160 ();
 sg13g2_decap_8 FILLER_0_68_1167 ();
 sg13g2_decap_8 FILLER_0_68_1174 ();
 sg13g2_decap_8 FILLER_0_68_1181 ();
 sg13g2_decap_8 FILLER_0_68_1188 ();
 sg13g2_decap_8 FILLER_0_68_1195 ();
 sg13g2_decap_8 FILLER_0_68_1202 ();
 sg13g2_decap_8 FILLER_0_68_1209 ();
 sg13g2_decap_8 FILLER_0_68_1216 ();
 sg13g2_decap_4 FILLER_0_68_1223 ();
 sg13g2_fill_1 FILLER_0_68_1227 ();
 sg13g2_decap_8 FILLER_0_69_0 ();
 sg13g2_decap_8 FILLER_0_69_7 ();
 sg13g2_decap_8 FILLER_0_69_14 ();
 sg13g2_decap_8 FILLER_0_69_21 ();
 sg13g2_decap_8 FILLER_0_69_28 ();
 sg13g2_decap_8 FILLER_0_69_35 ();
 sg13g2_decap_4 FILLER_0_69_42 ();
 sg13g2_fill_2 FILLER_0_69_46 ();
 sg13g2_decap_4 FILLER_0_69_57 ();
 sg13g2_fill_1 FILLER_0_69_61 ();
 sg13g2_fill_2 FILLER_0_69_72 ();
 sg13g2_fill_1 FILLER_0_69_74 ();
 sg13g2_fill_2 FILLER_0_69_83 ();
 sg13g2_fill_1 FILLER_0_69_85 ();
 sg13g2_decap_8 FILLER_0_69_101 ();
 sg13g2_decap_8 FILLER_0_69_108 ();
 sg13g2_decap_8 FILLER_0_69_115 ();
 sg13g2_decap_8 FILLER_0_69_122 ();
 sg13g2_decap_8 FILLER_0_69_129 ();
 sg13g2_fill_2 FILLER_0_69_136 ();
 sg13g2_decap_8 FILLER_0_69_143 ();
 sg13g2_decap_4 FILLER_0_69_150 ();
 sg13g2_fill_1 FILLER_0_69_154 ();
 sg13g2_fill_2 FILLER_0_69_196 ();
 sg13g2_decap_8 FILLER_0_69_228 ();
 sg13g2_decap_8 FILLER_0_69_235 ();
 sg13g2_decap_8 FILLER_0_69_242 ();
 sg13g2_decap_8 FILLER_0_69_249 ();
 sg13g2_decap_8 FILLER_0_69_256 ();
 sg13g2_decap_8 FILLER_0_69_263 ();
 sg13g2_decap_8 FILLER_0_69_270 ();
 sg13g2_decap_8 FILLER_0_69_277 ();
 sg13g2_decap_8 FILLER_0_69_284 ();
 sg13g2_decap_8 FILLER_0_69_291 ();
 sg13g2_decap_8 FILLER_0_69_298 ();
 sg13g2_fill_1 FILLER_0_69_305 ();
 sg13g2_fill_2 FILLER_0_69_315 ();
 sg13g2_fill_1 FILLER_0_69_343 ();
 sg13g2_decap_4 FILLER_0_69_353 ();
 sg13g2_decap_8 FILLER_0_69_367 ();
 sg13g2_decap_8 FILLER_0_69_374 ();
 sg13g2_decap_8 FILLER_0_69_381 ();
 sg13g2_decap_8 FILLER_0_69_388 ();
 sg13g2_decap_8 FILLER_0_69_395 ();
 sg13g2_decap_8 FILLER_0_69_402 ();
 sg13g2_decap_8 FILLER_0_69_409 ();
 sg13g2_decap_8 FILLER_0_69_416 ();
 sg13g2_decap_8 FILLER_0_69_423 ();
 sg13g2_fill_1 FILLER_0_69_430 ();
 sg13g2_fill_1 FILLER_0_69_457 ();
 sg13g2_fill_2 FILLER_0_69_489 ();
 sg13g2_fill_1 FILLER_0_69_491 ();
 sg13g2_decap_8 FILLER_0_69_581 ();
 sg13g2_fill_1 FILLER_0_69_647 ();
 sg13g2_decap_4 FILLER_0_69_658 ();
 sg13g2_fill_2 FILLER_0_69_662 ();
 sg13g2_decap_4 FILLER_0_69_675 ();
 sg13g2_fill_2 FILLER_0_69_679 ();
 sg13g2_fill_1 FILLER_0_69_685 ();
 sg13g2_fill_2 FILLER_0_69_696 ();
 sg13g2_fill_2 FILLER_0_69_708 ();
 sg13g2_fill_2 FILLER_0_69_740 ();
 sg13g2_fill_2 FILLER_0_69_747 ();
 sg13g2_decap_4 FILLER_0_69_754 ();
 sg13g2_fill_1 FILLER_0_69_758 ();
 sg13g2_decap_8 FILLER_0_69_764 ();
 sg13g2_decap_8 FILLER_0_69_771 ();
 sg13g2_decap_8 FILLER_0_69_778 ();
 sg13g2_fill_2 FILLER_0_69_785 ();
 sg13g2_fill_1 FILLER_0_69_795 ();
 sg13g2_decap_4 FILLER_0_69_801 ();
 sg13g2_decap_8 FILLER_0_69_809 ();
 sg13g2_decap_8 FILLER_0_69_816 ();
 sg13g2_decap_8 FILLER_0_69_823 ();
 sg13g2_decap_8 FILLER_0_69_830 ();
 sg13g2_decap_4 FILLER_0_69_837 ();
 sg13g2_decap_4 FILLER_0_69_867 ();
 sg13g2_fill_2 FILLER_0_69_871 ();
 sg13g2_fill_2 FILLER_0_69_883 ();
 sg13g2_decap_4 FILLER_0_69_890 ();
 sg13g2_fill_2 FILLER_0_69_894 ();
 sg13g2_decap_8 FILLER_0_69_918 ();
 sg13g2_decap_8 FILLER_0_69_925 ();
 sg13g2_fill_2 FILLER_0_69_932 ();
 sg13g2_decap_4 FILLER_0_69_938 ();
 sg13g2_fill_2 FILLER_0_69_942 ();
 sg13g2_decap_8 FILLER_0_69_952 ();
 sg13g2_fill_2 FILLER_0_69_959 ();
 sg13g2_fill_1 FILLER_0_69_961 ();
 sg13g2_fill_1 FILLER_0_69_966 ();
 sg13g2_decap_4 FILLER_0_69_1002 ();
 sg13g2_decap_8 FILLER_0_69_1042 ();
 sg13g2_decap_8 FILLER_0_69_1049 ();
 sg13g2_decap_8 FILLER_0_69_1056 ();
 sg13g2_decap_8 FILLER_0_69_1063 ();
 sg13g2_decap_8 FILLER_0_69_1070 ();
 sg13g2_decap_8 FILLER_0_69_1077 ();
 sg13g2_decap_8 FILLER_0_69_1084 ();
 sg13g2_decap_8 FILLER_0_69_1091 ();
 sg13g2_decap_8 FILLER_0_69_1098 ();
 sg13g2_decap_8 FILLER_0_69_1105 ();
 sg13g2_decap_8 FILLER_0_69_1112 ();
 sg13g2_decap_8 FILLER_0_69_1119 ();
 sg13g2_decap_8 FILLER_0_69_1126 ();
 sg13g2_decap_8 FILLER_0_69_1133 ();
 sg13g2_decap_8 FILLER_0_69_1140 ();
 sg13g2_decap_8 FILLER_0_69_1147 ();
 sg13g2_decap_8 FILLER_0_69_1154 ();
 sg13g2_decap_8 FILLER_0_69_1161 ();
 sg13g2_decap_8 FILLER_0_69_1168 ();
 sg13g2_decap_8 FILLER_0_69_1175 ();
 sg13g2_decap_8 FILLER_0_69_1182 ();
 sg13g2_decap_8 FILLER_0_69_1189 ();
 sg13g2_decap_8 FILLER_0_69_1196 ();
 sg13g2_decap_8 FILLER_0_69_1203 ();
 sg13g2_decap_8 FILLER_0_69_1210 ();
 sg13g2_decap_8 FILLER_0_69_1217 ();
 sg13g2_decap_4 FILLER_0_69_1224 ();
 sg13g2_decap_8 FILLER_0_70_0 ();
 sg13g2_decap_8 FILLER_0_70_7 ();
 sg13g2_decap_8 FILLER_0_70_14 ();
 sg13g2_decap_8 FILLER_0_70_21 ();
 sg13g2_decap_8 FILLER_0_70_28 ();
 sg13g2_decap_8 FILLER_0_70_35 ();
 sg13g2_decap_8 FILLER_0_70_68 ();
 sg13g2_decap_4 FILLER_0_70_75 ();
 sg13g2_fill_2 FILLER_0_70_105 ();
 sg13g2_decap_8 FILLER_0_70_143 ();
 sg13g2_decap_4 FILLER_0_70_150 ();
 sg13g2_fill_1 FILLER_0_70_154 ();
 sg13g2_fill_2 FILLER_0_70_216 ();
 sg13g2_fill_1 FILLER_0_70_218 ();
 sg13g2_decap_8 FILLER_0_70_224 ();
 sg13g2_decap_8 FILLER_0_70_231 ();
 sg13g2_decap_8 FILLER_0_70_238 ();
 sg13g2_decap_8 FILLER_0_70_245 ();
 sg13g2_decap_8 FILLER_0_70_252 ();
 sg13g2_decap_8 FILLER_0_70_259 ();
 sg13g2_decap_8 FILLER_0_70_266 ();
 sg13g2_decap_8 FILLER_0_70_273 ();
 sg13g2_decap_8 FILLER_0_70_280 ();
 sg13g2_decap_8 FILLER_0_70_287 ();
 sg13g2_decap_8 FILLER_0_70_294 ();
 sg13g2_fill_2 FILLER_0_70_301 ();
 sg13g2_decap_8 FILLER_0_70_360 ();
 sg13g2_decap_8 FILLER_0_70_367 ();
 sg13g2_decap_8 FILLER_0_70_374 ();
 sg13g2_decap_8 FILLER_0_70_381 ();
 sg13g2_decap_8 FILLER_0_70_388 ();
 sg13g2_decap_8 FILLER_0_70_395 ();
 sg13g2_decap_8 FILLER_0_70_402 ();
 sg13g2_decap_8 FILLER_0_70_409 ();
 sg13g2_decap_8 FILLER_0_70_416 ();
 sg13g2_decap_8 FILLER_0_70_423 ();
 sg13g2_decap_4 FILLER_0_70_430 ();
 sg13g2_fill_1 FILLER_0_70_434 ();
 sg13g2_decap_8 FILLER_0_70_439 ();
 sg13g2_decap_8 FILLER_0_70_446 ();
 sg13g2_decap_4 FILLER_0_70_453 ();
 sg13g2_decap_8 FILLER_0_70_493 ();
 sg13g2_decap_8 FILLER_0_70_500 ();
 sg13g2_fill_2 FILLER_0_70_507 ();
 sg13g2_fill_1 FILLER_0_70_528 ();
 sg13g2_fill_1 FILLER_0_70_539 ();
 sg13g2_fill_1 FILLER_0_70_544 ();
 sg13g2_fill_1 FILLER_0_70_553 ();
 sg13g2_fill_2 FILLER_0_70_564 ();
 sg13g2_decap_8 FILLER_0_70_570 ();
 sg13g2_decap_8 FILLER_0_70_577 ();
 sg13g2_decap_8 FILLER_0_70_584 ();
 sg13g2_fill_1 FILLER_0_70_591 ();
 sg13g2_decap_8 FILLER_0_70_640 ();
 sg13g2_decap_8 FILLER_0_70_647 ();
 sg13g2_decap_8 FILLER_0_70_654 ();
 sg13g2_fill_1 FILLER_0_70_661 ();
 sg13g2_fill_1 FILLER_0_70_682 ();
 sg13g2_decap_8 FILLER_0_70_693 ();
 sg13g2_decap_8 FILLER_0_70_700 ();
 sg13g2_decap_8 FILLER_0_70_776 ();
 sg13g2_decap_8 FILLER_0_70_783 ();
 sg13g2_decap_8 FILLER_0_70_790 ();
 sg13g2_decap_8 FILLER_0_70_797 ();
 sg13g2_decap_8 FILLER_0_70_804 ();
 sg13g2_decap_4 FILLER_0_70_811 ();
 sg13g2_decap_8 FILLER_0_70_830 ();
 sg13g2_decap_8 FILLER_0_70_837 ();
 sg13g2_decap_4 FILLER_0_70_844 ();
 sg13g2_fill_2 FILLER_0_70_848 ();
 sg13g2_decap_8 FILLER_0_70_854 ();
 sg13g2_decap_4 FILLER_0_70_866 ();
 sg13g2_fill_1 FILLER_0_70_870 ();
 sg13g2_decap_8 FILLER_0_70_881 ();
 sg13g2_fill_1 FILLER_0_70_888 ();
 sg13g2_decap_8 FILLER_0_70_914 ();
 sg13g2_decap_8 FILLER_0_70_921 ();
 sg13g2_decap_8 FILLER_0_70_928 ();
 sg13g2_decap_8 FILLER_0_70_935 ();
 sg13g2_decap_8 FILLER_0_70_942 ();
 sg13g2_decap_8 FILLER_0_70_949 ();
 sg13g2_decap_8 FILLER_0_70_956 ();
 sg13g2_decap_8 FILLER_0_70_963 ();
 sg13g2_decap_8 FILLER_0_70_970 ();
 sg13g2_decap_8 FILLER_0_70_977 ();
 sg13g2_decap_4 FILLER_0_70_984 ();
 sg13g2_fill_2 FILLER_0_70_988 ();
 sg13g2_decap_8 FILLER_0_70_1040 ();
 sg13g2_decap_8 FILLER_0_70_1047 ();
 sg13g2_decap_8 FILLER_0_70_1054 ();
 sg13g2_decap_8 FILLER_0_70_1061 ();
 sg13g2_decap_8 FILLER_0_70_1068 ();
 sg13g2_decap_8 FILLER_0_70_1075 ();
 sg13g2_decap_8 FILLER_0_70_1082 ();
 sg13g2_decap_8 FILLER_0_70_1089 ();
 sg13g2_decap_8 FILLER_0_70_1096 ();
 sg13g2_decap_8 FILLER_0_70_1103 ();
 sg13g2_decap_8 FILLER_0_70_1110 ();
 sg13g2_decap_8 FILLER_0_70_1117 ();
 sg13g2_decap_8 FILLER_0_70_1124 ();
 sg13g2_decap_8 FILLER_0_70_1131 ();
 sg13g2_decap_8 FILLER_0_70_1138 ();
 sg13g2_decap_8 FILLER_0_70_1145 ();
 sg13g2_decap_8 FILLER_0_70_1152 ();
 sg13g2_decap_8 FILLER_0_70_1159 ();
 sg13g2_decap_8 FILLER_0_70_1166 ();
 sg13g2_decap_8 FILLER_0_70_1173 ();
 sg13g2_decap_8 FILLER_0_70_1180 ();
 sg13g2_decap_8 FILLER_0_70_1187 ();
 sg13g2_decap_8 FILLER_0_70_1194 ();
 sg13g2_decap_8 FILLER_0_70_1201 ();
 sg13g2_decap_8 FILLER_0_70_1208 ();
 sg13g2_decap_8 FILLER_0_70_1215 ();
 sg13g2_decap_4 FILLER_0_70_1222 ();
 sg13g2_fill_2 FILLER_0_70_1226 ();
 sg13g2_decap_8 FILLER_0_71_0 ();
 sg13g2_decap_8 FILLER_0_71_7 ();
 sg13g2_decap_8 FILLER_0_71_14 ();
 sg13g2_decap_8 FILLER_0_71_21 ();
 sg13g2_decap_8 FILLER_0_71_28 ();
 sg13g2_fill_2 FILLER_0_71_35 ();
 sg13g2_fill_1 FILLER_0_71_37 ();
 sg13g2_decap_4 FILLER_0_71_68 ();
 sg13g2_fill_1 FILLER_0_71_72 ();
 sg13g2_fill_1 FILLER_0_71_78 ();
 sg13g2_fill_1 FILLER_0_71_126 ();
 sg13g2_decap_8 FILLER_0_71_158 ();
 sg13g2_fill_2 FILLER_0_71_165 ();
 sg13g2_fill_1 FILLER_0_71_167 ();
 sg13g2_fill_2 FILLER_0_71_172 ();
 sg13g2_fill_1 FILLER_0_71_174 ();
 sg13g2_fill_2 FILLER_0_71_180 ();
 sg13g2_fill_2 FILLER_0_71_198 ();
 sg13g2_decap_8 FILLER_0_71_221 ();
 sg13g2_decap_8 FILLER_0_71_228 ();
 sg13g2_decap_8 FILLER_0_71_235 ();
 sg13g2_decap_8 FILLER_0_71_242 ();
 sg13g2_decap_8 FILLER_0_71_249 ();
 sg13g2_decap_8 FILLER_0_71_256 ();
 sg13g2_decap_8 FILLER_0_71_263 ();
 sg13g2_decap_8 FILLER_0_71_270 ();
 sg13g2_decap_8 FILLER_0_71_277 ();
 sg13g2_decap_8 FILLER_0_71_284 ();
 sg13g2_decap_8 FILLER_0_71_291 ();
 sg13g2_fill_2 FILLER_0_71_298 ();
 sg13g2_fill_1 FILLER_0_71_300 ();
 sg13g2_fill_1 FILLER_0_71_306 ();
 sg13g2_fill_1 FILLER_0_71_312 ();
 sg13g2_fill_1 FILLER_0_71_333 ();
 sg13g2_decap_8 FILLER_0_71_374 ();
 sg13g2_fill_2 FILLER_0_71_381 ();
 sg13g2_decap_8 FILLER_0_71_386 ();
 sg13g2_decap_8 FILLER_0_71_393 ();
 sg13g2_decap_8 FILLER_0_71_400 ();
 sg13g2_decap_8 FILLER_0_71_420 ();
 sg13g2_decap_8 FILLER_0_71_427 ();
 sg13g2_decap_8 FILLER_0_71_434 ();
 sg13g2_decap_8 FILLER_0_71_441 ();
 sg13g2_fill_2 FILLER_0_71_448 ();
 sg13g2_fill_1 FILLER_0_71_463 ();
 sg13g2_decap_8 FILLER_0_71_509 ();
 sg13g2_decap_8 FILLER_0_71_516 ();
 sg13g2_decap_8 FILLER_0_71_523 ();
 sg13g2_decap_4 FILLER_0_71_530 ();
 sg13g2_fill_1 FILLER_0_71_534 ();
 sg13g2_decap_8 FILLER_0_71_539 ();
 sg13g2_decap_8 FILLER_0_71_546 ();
 sg13g2_decap_8 FILLER_0_71_553 ();
 sg13g2_decap_8 FILLER_0_71_560 ();
 sg13g2_decap_8 FILLER_0_71_567 ();
 sg13g2_decap_8 FILLER_0_71_574 ();
 sg13g2_decap_8 FILLER_0_71_581 ();
 sg13g2_decap_8 FILLER_0_71_588 ();
 sg13g2_fill_1 FILLER_0_71_595 ();
 sg13g2_decap_8 FILLER_0_71_634 ();
 sg13g2_fill_1 FILLER_0_71_646 ();
 sg13g2_fill_2 FILLER_0_71_652 ();
 sg13g2_decap_4 FILLER_0_71_690 ();
 sg13g2_fill_1 FILLER_0_71_694 ();
 sg13g2_decap_8 FILLER_0_71_700 ();
 sg13g2_fill_2 FILLER_0_71_707 ();
 sg13g2_fill_1 FILLER_0_71_709 ();
 sg13g2_decap_8 FILLER_0_71_725 ();
 sg13g2_fill_1 FILLER_0_71_732 ();
 sg13g2_decap_8 FILLER_0_71_737 ();
 sg13g2_fill_1 FILLER_0_71_744 ();
 sg13g2_fill_2 FILLER_0_71_759 ();
 sg13g2_fill_2 FILLER_0_71_787 ();
 sg13g2_fill_2 FILLER_0_71_794 ();
 sg13g2_fill_1 FILLER_0_71_796 ();
 sg13g2_fill_2 FILLER_0_71_828 ();
 sg13g2_fill_1 FILLER_0_71_830 ();
 sg13g2_decap_8 FILLER_0_71_887 ();
 sg13g2_decap_4 FILLER_0_71_894 ();
 sg13g2_decap_8 FILLER_0_71_929 ();
 sg13g2_decap_8 FILLER_0_71_936 ();
 sg13g2_decap_8 FILLER_0_71_943 ();
 sg13g2_decap_8 FILLER_0_71_950 ();
 sg13g2_decap_8 FILLER_0_71_957 ();
 sg13g2_decap_8 FILLER_0_71_1010 ();
 sg13g2_decap_8 FILLER_0_71_1017 ();
 sg13g2_fill_1 FILLER_0_71_1024 ();
 sg13g2_decap_8 FILLER_0_71_1035 ();
 sg13g2_decap_8 FILLER_0_71_1042 ();
 sg13g2_decap_8 FILLER_0_71_1049 ();
 sg13g2_decap_8 FILLER_0_71_1056 ();
 sg13g2_decap_8 FILLER_0_71_1063 ();
 sg13g2_decap_8 FILLER_0_71_1070 ();
 sg13g2_decap_8 FILLER_0_71_1077 ();
 sg13g2_decap_8 FILLER_0_71_1084 ();
 sg13g2_decap_8 FILLER_0_71_1091 ();
 sg13g2_decap_8 FILLER_0_71_1098 ();
 sg13g2_decap_8 FILLER_0_71_1105 ();
 sg13g2_decap_8 FILLER_0_71_1112 ();
 sg13g2_decap_8 FILLER_0_71_1119 ();
 sg13g2_decap_8 FILLER_0_71_1126 ();
 sg13g2_decap_8 FILLER_0_71_1133 ();
 sg13g2_decap_8 FILLER_0_71_1140 ();
 sg13g2_decap_8 FILLER_0_71_1147 ();
 sg13g2_decap_8 FILLER_0_71_1154 ();
 sg13g2_decap_8 FILLER_0_71_1161 ();
 sg13g2_decap_8 FILLER_0_71_1168 ();
 sg13g2_decap_8 FILLER_0_71_1175 ();
 sg13g2_decap_8 FILLER_0_71_1182 ();
 sg13g2_decap_8 FILLER_0_71_1189 ();
 sg13g2_decap_8 FILLER_0_71_1196 ();
 sg13g2_decap_8 FILLER_0_71_1203 ();
 sg13g2_decap_8 FILLER_0_71_1210 ();
 sg13g2_decap_8 FILLER_0_71_1217 ();
 sg13g2_decap_4 FILLER_0_71_1224 ();
 sg13g2_decap_8 FILLER_0_72_0 ();
 sg13g2_decap_8 FILLER_0_72_7 ();
 sg13g2_decap_8 FILLER_0_72_14 ();
 sg13g2_decap_8 FILLER_0_72_21 ();
 sg13g2_decap_8 FILLER_0_72_28 ();
 sg13g2_decap_8 FILLER_0_72_35 ();
 sg13g2_fill_2 FILLER_0_72_82 ();
 sg13g2_fill_1 FILLER_0_72_84 ();
 sg13g2_decap_4 FILLER_0_72_98 ();
 sg13g2_fill_1 FILLER_0_72_128 ();
 sg13g2_decap_8 FILLER_0_72_170 ();
 sg13g2_decap_4 FILLER_0_72_177 ();
 sg13g2_decap_8 FILLER_0_72_215 ();
 sg13g2_decap_8 FILLER_0_72_222 ();
 sg13g2_decap_8 FILLER_0_72_229 ();
 sg13g2_decap_8 FILLER_0_72_236 ();
 sg13g2_decap_8 FILLER_0_72_243 ();
 sg13g2_decap_8 FILLER_0_72_250 ();
 sg13g2_decap_8 FILLER_0_72_257 ();
 sg13g2_decap_8 FILLER_0_72_264 ();
 sg13g2_decap_8 FILLER_0_72_271 ();
 sg13g2_decap_8 FILLER_0_72_278 ();
 sg13g2_decap_8 FILLER_0_72_285 ();
 sg13g2_decap_8 FILLER_0_72_292 ();
 sg13g2_fill_2 FILLER_0_72_299 ();
 sg13g2_fill_2 FILLER_0_72_342 ();
 sg13g2_fill_1 FILLER_0_72_344 ();
 sg13g2_decap_8 FILLER_0_72_363 ();
 sg13g2_decap_4 FILLER_0_72_370 ();
 sg13g2_fill_2 FILLER_0_72_374 ();
 sg13g2_fill_2 FILLER_0_72_385 ();
 sg13g2_decap_8 FILLER_0_72_413 ();
 sg13g2_decap_8 FILLER_0_72_420 ();
 sg13g2_decap_8 FILLER_0_72_427 ();
 sg13g2_decap_8 FILLER_0_72_434 ();
 sg13g2_decap_8 FILLER_0_72_441 ();
 sg13g2_decap_8 FILLER_0_72_448 ();
 sg13g2_decap_4 FILLER_0_72_455 ();
 sg13g2_fill_1 FILLER_0_72_459 ();
 sg13g2_fill_1 FILLER_0_72_470 ();
 sg13g2_fill_2 FILLER_0_72_475 ();
 sg13g2_fill_1 FILLER_0_72_477 ();
 sg13g2_decap_8 FILLER_0_72_497 ();
 sg13g2_fill_1 FILLER_0_72_504 ();
 sg13g2_fill_2 FILLER_0_72_520 ();
 sg13g2_fill_1 FILLER_0_72_527 ();
 sg13g2_decap_8 FILLER_0_72_532 ();
 sg13g2_decap_8 FILLER_0_72_539 ();
 sg13g2_decap_4 FILLER_0_72_546 ();
 sg13g2_fill_1 FILLER_0_72_550 ();
 sg13g2_decap_8 FILLER_0_72_581 ();
 sg13g2_decap_8 FILLER_0_72_588 ();
 sg13g2_decap_8 FILLER_0_72_595 ();
 sg13g2_decap_4 FILLER_0_72_602 ();
 sg13g2_fill_1 FILLER_0_72_606 ();
 sg13g2_fill_1 FILLER_0_72_612 ();
 sg13g2_fill_1 FILLER_0_72_623 ();
 sg13g2_fill_1 FILLER_0_72_650 ();
 sg13g2_fill_1 FILLER_0_72_677 ();
 sg13g2_decap_8 FILLER_0_72_682 ();
 sg13g2_decap_4 FILLER_0_72_719 ();
 sg13g2_decap_4 FILLER_0_72_749 ();
 sg13g2_decap_8 FILLER_0_72_828 ();
 sg13g2_fill_2 FILLER_0_72_835 ();
 sg13g2_fill_2 FILLER_0_72_847 ();
 sg13g2_fill_1 FILLER_0_72_849 ();
 sg13g2_decap_8 FILLER_0_72_854 ();
 sg13g2_fill_2 FILLER_0_72_876 ();
 sg13g2_fill_1 FILLER_0_72_904 ();
 sg13g2_decap_8 FILLER_0_72_920 ();
 sg13g2_decap_8 FILLER_0_72_927 ();
 sg13g2_fill_1 FILLER_0_72_934 ();
 sg13g2_decap_4 FILLER_0_72_939 ();
 sg13g2_fill_2 FILLER_0_72_943 ();
 sg13g2_decap_8 FILLER_0_72_950 ();
 sg13g2_decap_8 FILLER_0_72_957 ();
 sg13g2_decap_8 FILLER_0_72_964 ();
 sg13g2_decap_8 FILLER_0_72_971 ();
 sg13g2_decap_8 FILLER_0_72_992 ();
 sg13g2_decap_8 FILLER_0_72_999 ();
 sg13g2_fill_2 FILLER_0_72_1006 ();
 sg13g2_fill_1 FILLER_0_72_1008 ();
 sg13g2_decap_4 FILLER_0_72_1013 ();
 sg13g2_fill_1 FILLER_0_72_1017 ();
 sg13g2_fill_1 FILLER_0_72_1022 ();
 sg13g2_decap_8 FILLER_0_72_1054 ();
 sg13g2_decap_8 FILLER_0_72_1061 ();
 sg13g2_decap_8 FILLER_0_72_1068 ();
 sg13g2_decap_8 FILLER_0_72_1075 ();
 sg13g2_decap_8 FILLER_0_72_1082 ();
 sg13g2_decap_8 FILLER_0_72_1089 ();
 sg13g2_decap_8 FILLER_0_72_1096 ();
 sg13g2_decap_8 FILLER_0_72_1103 ();
 sg13g2_decap_8 FILLER_0_72_1110 ();
 sg13g2_decap_8 FILLER_0_72_1117 ();
 sg13g2_decap_8 FILLER_0_72_1124 ();
 sg13g2_decap_8 FILLER_0_72_1131 ();
 sg13g2_decap_8 FILLER_0_72_1138 ();
 sg13g2_decap_8 FILLER_0_72_1145 ();
 sg13g2_decap_8 FILLER_0_72_1152 ();
 sg13g2_decap_8 FILLER_0_72_1159 ();
 sg13g2_decap_8 FILLER_0_72_1166 ();
 sg13g2_decap_8 FILLER_0_72_1173 ();
 sg13g2_decap_8 FILLER_0_72_1180 ();
 sg13g2_decap_8 FILLER_0_72_1187 ();
 sg13g2_decap_8 FILLER_0_72_1194 ();
 sg13g2_decap_8 FILLER_0_72_1201 ();
 sg13g2_decap_8 FILLER_0_72_1208 ();
 sg13g2_decap_8 FILLER_0_72_1215 ();
 sg13g2_decap_4 FILLER_0_72_1222 ();
 sg13g2_fill_2 FILLER_0_72_1226 ();
 sg13g2_decap_8 FILLER_0_73_0 ();
 sg13g2_decap_8 FILLER_0_73_7 ();
 sg13g2_decap_8 FILLER_0_73_14 ();
 sg13g2_decap_8 FILLER_0_73_21 ();
 sg13g2_decap_8 FILLER_0_73_28 ();
 sg13g2_decap_8 FILLER_0_73_35 ();
 sg13g2_decap_4 FILLER_0_73_42 ();
 sg13g2_fill_1 FILLER_0_73_55 ();
 sg13g2_decap_8 FILLER_0_73_74 ();
 sg13g2_decap_8 FILLER_0_73_81 ();
 sg13g2_decap_8 FILLER_0_73_88 ();
 sg13g2_decap_4 FILLER_0_73_95 ();
 sg13g2_fill_1 FILLER_0_73_99 ();
 sg13g2_fill_1 FILLER_0_73_105 ();
 sg13g2_fill_1 FILLER_0_73_110 ();
 sg13g2_fill_1 FILLER_0_73_121 ();
 sg13g2_fill_1 FILLER_0_73_132 ();
 sg13g2_decap_4 FILLER_0_73_142 ();
 sg13g2_decap_4 FILLER_0_73_150 ();
 sg13g2_fill_1 FILLER_0_73_154 ();
 sg13g2_fill_1 FILLER_0_73_181 ();
 sg13g2_decap_8 FILLER_0_73_227 ();
 sg13g2_decap_8 FILLER_0_73_234 ();
 sg13g2_decap_8 FILLER_0_73_241 ();
 sg13g2_decap_8 FILLER_0_73_248 ();
 sg13g2_decap_8 FILLER_0_73_255 ();
 sg13g2_decap_8 FILLER_0_73_262 ();
 sg13g2_decap_8 FILLER_0_73_269 ();
 sg13g2_decap_8 FILLER_0_73_276 ();
 sg13g2_decap_8 FILLER_0_73_283 ();
 sg13g2_decap_8 FILLER_0_73_290 ();
 sg13g2_decap_8 FILLER_0_73_297 ();
 sg13g2_decap_4 FILLER_0_73_304 ();
 sg13g2_fill_2 FILLER_0_73_368 ();
 sg13g2_fill_1 FILLER_0_73_396 ();
 sg13g2_fill_1 FILLER_0_73_402 ();
 sg13g2_fill_2 FILLER_0_73_429 ();
 sg13g2_fill_2 FILLER_0_73_477 ();
 sg13g2_fill_1 FILLER_0_73_520 ();
 sg13g2_decap_4 FILLER_0_73_547 ();
 sg13g2_fill_1 FILLER_0_73_551 ();
 sg13g2_decap_8 FILLER_0_73_603 ();
 sg13g2_fill_2 FILLER_0_73_610 ();
 sg13g2_fill_2 FILLER_0_73_667 ();
 sg13g2_fill_1 FILLER_0_73_669 ();
 sg13g2_fill_1 FILLER_0_73_675 ();
 sg13g2_fill_2 FILLER_0_73_711 ();
 sg13g2_decap_8 FILLER_0_73_737 ();
 sg13g2_decap_4 FILLER_0_73_744 ();
 sg13g2_fill_2 FILLER_0_73_748 ();
 sg13g2_fill_1 FILLER_0_73_760 ();
 sg13g2_fill_1 FILLER_0_73_766 ();
 sg13g2_fill_1 FILLER_0_73_771 ();
 sg13g2_fill_1 FILLER_0_73_798 ();
 sg13g2_fill_1 FILLER_0_73_803 ();
 sg13g2_decap_4 FILLER_0_73_808 ();
 sg13g2_decap_4 FILLER_0_73_822 ();
 sg13g2_fill_2 FILLER_0_73_861 ();
 sg13g2_fill_1 FILLER_0_73_863 ();
 sg13g2_fill_2 FILLER_0_73_894 ();
 sg13g2_decap_8 FILLER_0_73_953 ();
 sg13g2_decap_4 FILLER_0_73_960 ();
 sg13g2_fill_2 FILLER_0_73_964 ();
 sg13g2_decap_8 FILLER_0_73_992 ();
 sg13g2_decap_8 FILLER_0_73_999 ();
 sg13g2_fill_2 FILLER_0_73_1006 ();
 sg13g2_decap_4 FILLER_0_73_1013 ();
 sg13g2_fill_1 FILLER_0_73_1017 ();
 sg13g2_decap_8 FILLER_0_73_1028 ();
 sg13g2_decap_8 FILLER_0_73_1035 ();
 sg13g2_decap_8 FILLER_0_73_1042 ();
 sg13g2_decap_8 FILLER_0_73_1049 ();
 sg13g2_decap_8 FILLER_0_73_1056 ();
 sg13g2_decap_8 FILLER_0_73_1063 ();
 sg13g2_decap_8 FILLER_0_73_1070 ();
 sg13g2_decap_8 FILLER_0_73_1077 ();
 sg13g2_decap_8 FILLER_0_73_1084 ();
 sg13g2_decap_8 FILLER_0_73_1091 ();
 sg13g2_decap_8 FILLER_0_73_1098 ();
 sg13g2_decap_8 FILLER_0_73_1105 ();
 sg13g2_decap_8 FILLER_0_73_1112 ();
 sg13g2_decap_8 FILLER_0_73_1119 ();
 sg13g2_decap_8 FILLER_0_73_1126 ();
 sg13g2_decap_8 FILLER_0_73_1133 ();
 sg13g2_decap_8 FILLER_0_73_1140 ();
 sg13g2_decap_8 FILLER_0_73_1147 ();
 sg13g2_decap_8 FILLER_0_73_1154 ();
 sg13g2_decap_8 FILLER_0_73_1161 ();
 sg13g2_decap_8 FILLER_0_73_1168 ();
 sg13g2_decap_8 FILLER_0_73_1175 ();
 sg13g2_decap_8 FILLER_0_73_1182 ();
 sg13g2_decap_8 FILLER_0_73_1189 ();
 sg13g2_decap_8 FILLER_0_73_1196 ();
 sg13g2_decap_8 FILLER_0_73_1203 ();
 sg13g2_decap_8 FILLER_0_73_1210 ();
 sg13g2_decap_8 FILLER_0_73_1217 ();
 sg13g2_decap_4 FILLER_0_73_1224 ();
 sg13g2_decap_8 FILLER_0_74_0 ();
 sg13g2_decap_8 FILLER_0_74_7 ();
 sg13g2_decap_8 FILLER_0_74_14 ();
 sg13g2_decap_8 FILLER_0_74_21 ();
 sg13g2_decap_8 FILLER_0_74_28 ();
 sg13g2_decap_4 FILLER_0_74_35 ();
 sg13g2_fill_2 FILLER_0_74_39 ();
 sg13g2_decap_8 FILLER_0_74_45 ();
 sg13g2_fill_2 FILLER_0_74_52 ();
 sg13g2_fill_1 FILLER_0_74_54 ();
 sg13g2_decap_4 FILLER_0_74_60 ();
 sg13g2_fill_1 FILLER_0_74_64 ();
 sg13g2_decap_8 FILLER_0_74_75 ();
 sg13g2_decap_8 FILLER_0_74_82 ();
 sg13g2_decap_8 FILLER_0_74_89 ();
 sg13g2_decap_8 FILLER_0_74_96 ();
 sg13g2_decap_8 FILLER_0_74_103 ();
 sg13g2_decap_8 FILLER_0_74_110 ();
 sg13g2_fill_2 FILLER_0_74_117 ();
 sg13g2_fill_1 FILLER_0_74_131 ();
 sg13g2_fill_2 FILLER_0_74_142 ();
 sg13g2_decap_4 FILLER_0_74_149 ();
 sg13g2_fill_2 FILLER_0_74_153 ();
 sg13g2_fill_1 FILLER_0_74_169 ();
 sg13g2_fill_2 FILLER_0_74_200 ();
 sg13g2_fill_1 FILLER_0_74_202 ();
 sg13g2_fill_2 FILLER_0_74_213 ();
 sg13g2_fill_1 FILLER_0_74_225 ();
 sg13g2_decap_8 FILLER_0_74_230 ();
 sg13g2_decap_8 FILLER_0_74_237 ();
 sg13g2_decap_4 FILLER_0_74_244 ();
 sg13g2_decap_4 FILLER_0_74_274 ();
 sg13g2_fill_2 FILLER_0_74_278 ();
 sg13g2_fill_2 FILLER_0_74_342 ();
 sg13g2_fill_1 FILLER_0_74_344 ();
 sg13g2_decap_4 FILLER_0_74_349 ();
 sg13g2_fill_1 FILLER_0_74_353 ();
 sg13g2_fill_2 FILLER_0_74_380 ();
 sg13g2_fill_1 FILLER_0_74_444 ();
 sg13g2_decap_8 FILLER_0_74_471 ();
 sg13g2_decap_8 FILLER_0_74_478 ();
 sg13g2_fill_2 FILLER_0_74_485 ();
 sg13g2_fill_1 FILLER_0_74_491 ();
 sg13g2_fill_1 FILLER_0_74_518 ();
 sg13g2_decap_8 FILLER_0_74_554 ();
 sg13g2_fill_1 FILLER_0_74_561 ();
 sg13g2_decap_4 FILLER_0_74_566 ();
 sg13g2_fill_2 FILLER_0_74_570 ();
 sg13g2_decap_8 FILLER_0_74_616 ();
 sg13g2_decap_8 FILLER_0_74_623 ();
 sg13g2_fill_1 FILLER_0_74_630 ();
 sg13g2_decap_8 FILLER_0_74_635 ();
 sg13g2_fill_2 FILLER_0_74_642 ();
 sg13g2_decap_8 FILLER_0_74_658 ();
 sg13g2_fill_2 FILLER_0_74_665 ();
 sg13g2_fill_1 FILLER_0_74_667 ();
 sg13g2_decap_4 FILLER_0_74_677 ();
 sg13g2_decap_4 FILLER_0_74_686 ();
 sg13g2_fill_2 FILLER_0_74_690 ();
 sg13g2_fill_1 FILLER_0_74_702 ();
 sg13g2_decap_4 FILLER_0_74_747 ();
 sg13g2_decap_8 FILLER_0_74_756 ();
 sg13g2_decap_8 FILLER_0_74_763 ();
 sg13g2_fill_1 FILLER_0_74_770 ();
 sg13g2_fill_1 FILLER_0_74_790 ();
 sg13g2_fill_1 FILLER_0_74_817 ();
 sg13g2_decap_4 FILLER_0_74_822 ();
 sg13g2_fill_2 FILLER_0_74_826 ();
 sg13g2_decap_8 FILLER_0_74_847 ();
 sg13g2_decap_8 FILLER_0_74_854 ();
 sg13g2_decap_4 FILLER_0_74_861 ();
 sg13g2_fill_1 FILLER_0_74_865 ();
 sg13g2_decap_8 FILLER_0_74_881 ();
 sg13g2_decap_4 FILLER_0_74_888 ();
 sg13g2_fill_1 FILLER_0_74_892 ();
 sg13g2_fill_2 FILLER_0_74_906 ();
 sg13g2_fill_2 FILLER_0_74_922 ();
 sg13g2_fill_1 FILLER_0_74_924 ();
 sg13g2_decap_4 FILLER_0_74_930 ();
 sg13g2_fill_2 FILLER_0_74_934 ();
 sg13g2_fill_1 FILLER_0_74_948 ();
 sg13g2_decap_8 FILLER_0_74_993 ();
 sg13g2_decap_8 FILLER_0_74_1000 ();
 sg13g2_decap_8 FILLER_0_74_1033 ();
 sg13g2_decap_8 FILLER_0_74_1040 ();
 sg13g2_decap_8 FILLER_0_74_1047 ();
 sg13g2_decap_8 FILLER_0_74_1054 ();
 sg13g2_decap_8 FILLER_0_74_1061 ();
 sg13g2_decap_8 FILLER_0_74_1068 ();
 sg13g2_decap_8 FILLER_0_74_1075 ();
 sg13g2_decap_8 FILLER_0_74_1082 ();
 sg13g2_decap_8 FILLER_0_74_1089 ();
 sg13g2_decap_8 FILLER_0_74_1096 ();
 sg13g2_decap_8 FILLER_0_74_1103 ();
 sg13g2_decap_8 FILLER_0_74_1110 ();
 sg13g2_decap_8 FILLER_0_74_1117 ();
 sg13g2_decap_8 FILLER_0_74_1124 ();
 sg13g2_decap_8 FILLER_0_74_1131 ();
 sg13g2_decap_8 FILLER_0_74_1138 ();
 sg13g2_decap_8 FILLER_0_74_1145 ();
 sg13g2_decap_8 FILLER_0_74_1152 ();
 sg13g2_decap_8 FILLER_0_74_1159 ();
 sg13g2_decap_8 FILLER_0_74_1166 ();
 sg13g2_decap_8 FILLER_0_74_1173 ();
 sg13g2_decap_8 FILLER_0_74_1180 ();
 sg13g2_decap_8 FILLER_0_74_1187 ();
 sg13g2_decap_8 FILLER_0_74_1194 ();
 sg13g2_decap_8 FILLER_0_74_1201 ();
 sg13g2_decap_8 FILLER_0_74_1208 ();
 sg13g2_decap_8 FILLER_0_74_1215 ();
 sg13g2_decap_4 FILLER_0_74_1222 ();
 sg13g2_fill_2 FILLER_0_74_1226 ();
 sg13g2_decap_8 FILLER_0_75_0 ();
 sg13g2_decap_8 FILLER_0_75_7 ();
 sg13g2_decap_8 FILLER_0_75_14 ();
 sg13g2_decap_8 FILLER_0_75_21 ();
 sg13g2_decap_8 FILLER_0_75_28 ();
 sg13g2_decap_8 FILLER_0_75_35 ();
 sg13g2_decap_8 FILLER_0_75_42 ();
 sg13g2_fill_2 FILLER_0_75_49 ();
 sg13g2_fill_2 FILLER_0_75_87 ();
 sg13g2_fill_1 FILLER_0_75_89 ();
 sg13g2_decap_8 FILLER_0_75_120 ();
 sg13g2_decap_8 FILLER_0_75_127 ();
 sg13g2_decap_4 FILLER_0_75_134 ();
 sg13g2_decap_4 FILLER_0_75_142 ();
 sg13g2_decap_8 FILLER_0_75_151 ();
 sg13g2_decap_4 FILLER_0_75_158 ();
 sg13g2_fill_2 FILLER_0_75_162 ();
 sg13g2_decap_4 FILLER_0_75_183 ();
 sg13g2_fill_2 FILLER_0_75_187 ();
 sg13g2_decap_8 FILLER_0_75_193 ();
 sg13g2_fill_2 FILLER_0_75_200 ();
 sg13g2_decap_8 FILLER_0_75_237 ();
 sg13g2_decap_4 FILLER_0_75_244 ();
 sg13g2_fill_2 FILLER_0_75_248 ();
 sg13g2_fill_1 FILLER_0_75_259 ();
 sg13g2_decap_8 FILLER_0_75_326 ();
 sg13g2_decap_8 FILLER_0_75_333 ();
 sg13g2_decap_8 FILLER_0_75_340 ();
 sg13g2_decap_8 FILLER_0_75_347 ();
 sg13g2_fill_1 FILLER_0_75_359 ();
 sg13g2_fill_1 FILLER_0_75_364 ();
 sg13g2_fill_1 FILLER_0_75_375 ();
 sg13g2_decap_4 FILLER_0_75_395 ();
 sg13g2_fill_1 FILLER_0_75_399 ();
 sg13g2_fill_2 FILLER_0_75_405 ();
 sg13g2_fill_1 FILLER_0_75_412 ();
 sg13g2_fill_1 FILLER_0_75_423 ();
 sg13g2_fill_2 FILLER_0_75_428 ();
 sg13g2_fill_2 FILLER_0_75_440 ();
 sg13g2_fill_2 FILLER_0_75_446 ();
 sg13g2_fill_1 FILLER_0_75_448 ();
 sg13g2_decap_4 FILLER_0_75_492 ();
 sg13g2_fill_2 FILLER_0_75_496 ();
 sg13g2_decap_8 FILLER_0_75_502 ();
 sg13g2_decap_8 FILLER_0_75_509 ();
 sg13g2_fill_2 FILLER_0_75_516 ();
 sg13g2_fill_1 FILLER_0_75_518 ();
 sg13g2_decap_8 FILLER_0_75_550 ();
 sg13g2_decap_8 FILLER_0_75_557 ();
 sg13g2_decap_4 FILLER_0_75_564 ();
 sg13g2_fill_1 FILLER_0_75_583 ();
 sg13g2_decap_4 FILLER_0_75_589 ();
 sg13g2_fill_1 FILLER_0_75_593 ();
 sg13g2_decap_8 FILLER_0_75_608 ();
 sg13g2_decap_8 FILLER_0_75_615 ();
 sg13g2_decap_8 FILLER_0_75_622 ();
 sg13g2_decap_8 FILLER_0_75_629 ();
 sg13g2_decap_8 FILLER_0_75_636 ();
 sg13g2_decap_8 FILLER_0_75_643 ();
 sg13g2_decap_8 FILLER_0_75_650 ();
 sg13g2_decap_8 FILLER_0_75_657 ();
 sg13g2_decap_8 FILLER_0_75_669 ();
 sg13g2_fill_2 FILLER_0_75_676 ();
 sg13g2_fill_1 FILLER_0_75_678 ();
 sg13g2_decap_8 FILLER_0_75_705 ();
 sg13g2_decap_4 FILLER_0_75_712 ();
 sg13g2_fill_1 FILLER_0_75_716 ();
 sg13g2_fill_1 FILLER_0_75_758 ();
 sg13g2_decap_8 FILLER_0_75_767 ();
 sg13g2_fill_2 FILLER_0_75_774 ();
 sg13g2_fill_1 FILLER_0_75_776 ();
 sg13g2_decap_4 FILLER_0_75_782 ();
 sg13g2_fill_2 FILLER_0_75_791 ();
 sg13g2_decap_4 FILLER_0_75_807 ();
 sg13g2_fill_2 FILLER_0_75_811 ();
 sg13g2_decap_8 FILLER_0_75_857 ();
 sg13g2_fill_1 FILLER_0_75_864 ();
 sg13g2_fill_1 FILLER_0_75_870 ();
 sg13g2_decap_4 FILLER_0_75_885 ();
 sg13g2_fill_2 FILLER_0_75_889 ();
 sg13g2_decap_8 FILLER_0_75_896 ();
 sg13g2_decap_8 FILLER_0_75_903 ();
 sg13g2_decap_8 FILLER_0_75_910 ();
 sg13g2_fill_2 FILLER_0_75_917 ();
 sg13g2_decap_8 FILLER_0_75_997 ();
 sg13g2_fill_2 FILLER_0_75_1004 ();
 sg13g2_fill_1 FILLER_0_75_1006 ();
 sg13g2_decap_8 FILLER_0_75_1037 ();
 sg13g2_decap_8 FILLER_0_75_1044 ();
 sg13g2_decap_8 FILLER_0_75_1051 ();
 sg13g2_decap_8 FILLER_0_75_1058 ();
 sg13g2_decap_8 FILLER_0_75_1065 ();
 sg13g2_decap_8 FILLER_0_75_1072 ();
 sg13g2_decap_8 FILLER_0_75_1079 ();
 sg13g2_decap_8 FILLER_0_75_1086 ();
 sg13g2_decap_8 FILLER_0_75_1093 ();
 sg13g2_decap_8 FILLER_0_75_1100 ();
 sg13g2_decap_8 FILLER_0_75_1107 ();
 sg13g2_decap_8 FILLER_0_75_1114 ();
 sg13g2_decap_8 FILLER_0_75_1121 ();
 sg13g2_decap_8 FILLER_0_75_1128 ();
 sg13g2_decap_8 FILLER_0_75_1135 ();
 sg13g2_decap_8 FILLER_0_75_1142 ();
 sg13g2_decap_8 FILLER_0_75_1149 ();
 sg13g2_decap_8 FILLER_0_75_1156 ();
 sg13g2_decap_8 FILLER_0_75_1163 ();
 sg13g2_decap_8 FILLER_0_75_1170 ();
 sg13g2_decap_8 FILLER_0_75_1177 ();
 sg13g2_decap_8 FILLER_0_75_1184 ();
 sg13g2_decap_8 FILLER_0_75_1191 ();
 sg13g2_decap_8 FILLER_0_75_1198 ();
 sg13g2_decap_8 FILLER_0_75_1205 ();
 sg13g2_decap_8 FILLER_0_75_1212 ();
 sg13g2_decap_8 FILLER_0_75_1219 ();
 sg13g2_fill_2 FILLER_0_75_1226 ();
 sg13g2_decap_8 FILLER_0_76_0 ();
 sg13g2_decap_8 FILLER_0_76_7 ();
 sg13g2_decap_8 FILLER_0_76_14 ();
 sg13g2_decap_8 FILLER_0_76_21 ();
 sg13g2_decap_8 FILLER_0_76_28 ();
 sg13g2_decap_8 FILLER_0_76_35 ();
 sg13g2_decap_8 FILLER_0_76_42 ();
 sg13g2_decap_8 FILLER_0_76_49 ();
 sg13g2_fill_2 FILLER_0_76_56 ();
 sg13g2_fill_1 FILLER_0_76_62 ();
 sg13g2_fill_1 FILLER_0_76_68 ();
 sg13g2_fill_1 FILLER_0_76_95 ();
 sg13g2_fill_1 FILLER_0_76_101 ();
 sg13g2_decap_4 FILLER_0_76_128 ();
 sg13g2_decap_8 FILLER_0_76_158 ();
 sg13g2_decap_8 FILLER_0_76_165 ();
 sg13g2_fill_2 FILLER_0_76_172 ();
 sg13g2_fill_1 FILLER_0_76_179 ();
 sg13g2_decap_8 FILLER_0_76_184 ();
 sg13g2_fill_1 FILLER_0_76_191 ();
 sg13g2_decap_4 FILLER_0_76_196 ();
 sg13g2_fill_1 FILLER_0_76_200 ();
 sg13g2_decap_8 FILLER_0_76_228 ();
 sg13g2_decap_4 FILLER_0_76_235 ();
 sg13g2_fill_2 FILLER_0_76_239 ();
 sg13g2_fill_2 FILLER_0_76_267 ();
 sg13g2_fill_1 FILLER_0_76_294 ();
 sg13g2_decap_8 FILLER_0_76_303 ();
 sg13g2_decap_8 FILLER_0_76_320 ();
 sg13g2_decap_8 FILLER_0_76_327 ();
 sg13g2_decap_8 FILLER_0_76_334 ();
 sg13g2_decap_4 FILLER_0_76_341 ();
 sg13g2_fill_2 FILLER_0_76_345 ();
 sg13g2_decap_8 FILLER_0_76_358 ();
 sg13g2_decap_8 FILLER_0_76_365 ();
 sg13g2_decap_8 FILLER_0_76_372 ();
 sg13g2_decap_8 FILLER_0_76_379 ();
 sg13g2_decap_8 FILLER_0_76_386 ();
 sg13g2_decap_8 FILLER_0_76_393 ();
 sg13g2_decap_8 FILLER_0_76_400 ();
 sg13g2_decap_8 FILLER_0_76_407 ();
 sg13g2_decap_8 FILLER_0_76_414 ();
 sg13g2_decap_8 FILLER_0_76_421 ();
 sg13g2_decap_4 FILLER_0_76_428 ();
 sg13g2_fill_2 FILLER_0_76_432 ();
 sg13g2_decap_4 FILLER_0_76_439 ();
 sg13g2_fill_2 FILLER_0_76_452 ();
 sg13g2_fill_2 FILLER_0_76_459 ();
 sg13g2_fill_2 FILLER_0_76_489 ();
 sg13g2_fill_1 FILLER_0_76_491 ();
 sg13g2_decap_8 FILLER_0_76_501 ();
 sg13g2_fill_2 FILLER_0_76_508 ();
 sg13g2_decap_4 FILLER_0_76_541 ();
 sg13g2_decap_8 FILLER_0_76_576 ();
 sg13g2_fill_2 FILLER_0_76_583 ();
 sg13g2_fill_1 FILLER_0_76_585 ();
 sg13g2_decap_8 FILLER_0_76_612 ();
 sg13g2_decap_8 FILLER_0_76_619 ();
 sg13g2_decap_8 FILLER_0_76_626 ();
 sg13g2_decap_8 FILLER_0_76_633 ();
 sg13g2_decap_8 FILLER_0_76_640 ();
 sg13g2_decap_8 FILLER_0_76_647 ();
 sg13g2_decap_8 FILLER_0_76_654 ();
 sg13g2_fill_2 FILLER_0_76_661 ();
 sg13g2_fill_1 FILLER_0_76_663 ();
 sg13g2_fill_1 FILLER_0_76_675 ();
 sg13g2_decap_8 FILLER_0_76_707 ();
 sg13g2_decap_8 FILLER_0_76_714 ();
 sg13g2_fill_2 FILLER_0_76_721 ();
 sg13g2_fill_1 FILLER_0_76_723 ();
 sg13g2_decap_8 FILLER_0_76_775 ();
 sg13g2_decap_8 FILLER_0_76_782 ();
 sg13g2_decap_8 FILLER_0_76_789 ();
 sg13g2_decap_8 FILLER_0_76_796 ();
 sg13g2_decap_8 FILLER_0_76_803 ();
 sg13g2_decap_8 FILLER_0_76_810 ();
 sg13g2_fill_1 FILLER_0_76_817 ();
 sg13g2_decap_8 FILLER_0_76_849 ();
 sg13g2_decap_8 FILLER_0_76_856 ();
 sg13g2_fill_1 FILLER_0_76_863 ();
 sg13g2_fill_1 FILLER_0_76_894 ();
 sg13g2_fill_1 FILLER_0_76_926 ();
 sg13g2_fill_2 FILLER_0_76_958 ();
 sg13g2_fill_1 FILLER_0_76_960 ();
 sg13g2_decap_8 FILLER_0_76_997 ();
 sg13g2_decap_4 FILLER_0_76_1004 ();
 sg13g2_decap_8 FILLER_0_76_1027 ();
 sg13g2_decap_8 FILLER_0_76_1034 ();
 sg13g2_decap_8 FILLER_0_76_1041 ();
 sg13g2_decap_8 FILLER_0_76_1048 ();
 sg13g2_decap_8 FILLER_0_76_1055 ();
 sg13g2_decap_8 FILLER_0_76_1062 ();
 sg13g2_decap_8 FILLER_0_76_1069 ();
 sg13g2_decap_8 FILLER_0_76_1076 ();
 sg13g2_decap_8 FILLER_0_76_1083 ();
 sg13g2_decap_8 FILLER_0_76_1090 ();
 sg13g2_decap_8 FILLER_0_76_1097 ();
 sg13g2_decap_8 FILLER_0_76_1104 ();
 sg13g2_decap_8 FILLER_0_76_1111 ();
 sg13g2_decap_8 FILLER_0_76_1118 ();
 sg13g2_decap_8 FILLER_0_76_1125 ();
 sg13g2_decap_8 FILLER_0_76_1132 ();
 sg13g2_decap_8 FILLER_0_76_1139 ();
 sg13g2_decap_8 FILLER_0_76_1146 ();
 sg13g2_decap_8 FILLER_0_76_1153 ();
 sg13g2_decap_8 FILLER_0_76_1160 ();
 sg13g2_decap_8 FILLER_0_76_1167 ();
 sg13g2_decap_8 FILLER_0_76_1174 ();
 sg13g2_decap_8 FILLER_0_76_1181 ();
 sg13g2_decap_8 FILLER_0_76_1188 ();
 sg13g2_decap_8 FILLER_0_76_1195 ();
 sg13g2_decap_8 FILLER_0_76_1202 ();
 sg13g2_decap_8 FILLER_0_76_1209 ();
 sg13g2_decap_8 FILLER_0_76_1216 ();
 sg13g2_decap_4 FILLER_0_76_1223 ();
 sg13g2_fill_1 FILLER_0_76_1227 ();
 sg13g2_decap_8 FILLER_0_77_0 ();
 sg13g2_decap_8 FILLER_0_77_7 ();
 sg13g2_decap_8 FILLER_0_77_14 ();
 sg13g2_decap_8 FILLER_0_77_21 ();
 sg13g2_decap_8 FILLER_0_77_28 ();
 sg13g2_decap_8 FILLER_0_77_35 ();
 sg13g2_decap_8 FILLER_0_77_42 ();
 sg13g2_decap_8 FILLER_0_77_49 ();
 sg13g2_decap_4 FILLER_0_77_56 ();
 sg13g2_fill_2 FILLER_0_77_60 ();
 sg13g2_fill_1 FILLER_0_77_66 ();
 sg13g2_fill_2 FILLER_0_77_93 ();
 sg13g2_fill_2 FILLER_0_77_105 ();
 sg13g2_fill_1 FILLER_0_77_107 ();
 sg13g2_fill_1 FILLER_0_77_134 ();
 sg13g2_fill_2 FILLER_0_77_140 ();
 sg13g2_fill_1 FILLER_0_77_142 ();
 sg13g2_decap_4 FILLER_0_77_169 ();
 sg13g2_decap_8 FILLER_0_77_199 ();
 sg13g2_decap_4 FILLER_0_77_236 ();
 sg13g2_fill_1 FILLER_0_77_240 ();
 sg13g2_decap_8 FILLER_0_77_278 ();
 sg13g2_decap_8 FILLER_0_77_285 ();
 sg13g2_decap_8 FILLER_0_77_292 ();
 sg13g2_decap_8 FILLER_0_77_299 ();
 sg13g2_decap_8 FILLER_0_77_306 ();
 sg13g2_decap_8 FILLER_0_77_313 ();
 sg13g2_decap_8 FILLER_0_77_320 ();
 sg13g2_fill_2 FILLER_0_77_327 ();
 sg13g2_fill_1 FILLER_0_77_329 ();
 sg13g2_fill_2 FILLER_0_77_334 ();
 sg13g2_decap_8 FILLER_0_77_341 ();
 sg13g2_decap_4 FILLER_0_77_348 ();
 sg13g2_fill_2 FILLER_0_77_362 ();
 sg13g2_decap_8 FILLER_0_77_395 ();
 sg13g2_decap_8 FILLER_0_77_402 ();
 sg13g2_decap_8 FILLER_0_77_409 ();
 sg13g2_decap_8 FILLER_0_77_416 ();
 sg13g2_decap_8 FILLER_0_77_423 ();
 sg13g2_decap_8 FILLER_0_77_430 ();
 sg13g2_fill_2 FILLER_0_77_437 ();
 sg13g2_fill_1 FILLER_0_77_439 ();
 sg13g2_fill_1 FILLER_0_77_451 ();
 sg13g2_fill_2 FILLER_0_77_478 ();
 sg13g2_fill_1 FILLER_0_77_480 ();
 sg13g2_fill_2 FILLER_0_77_547 ();
 sg13g2_fill_1 FILLER_0_77_558 ();
 sg13g2_decap_8 FILLER_0_77_579 ();
 sg13g2_decap_8 FILLER_0_77_586 ();
 sg13g2_fill_1 FILLER_0_77_593 ();
 sg13g2_fill_2 FILLER_0_77_630 ();
 sg13g2_fill_1 FILLER_0_77_632 ();
 sg13g2_decap_8 FILLER_0_77_637 ();
 sg13g2_decap_8 FILLER_0_77_644 ();
 sg13g2_decap_8 FILLER_0_77_651 ();
 sg13g2_decap_8 FILLER_0_77_658 ();
 sg13g2_decap_8 FILLER_0_77_665 ();
 sg13g2_decap_8 FILLER_0_77_672 ();
 sg13g2_decap_8 FILLER_0_77_679 ();
 sg13g2_decap_8 FILLER_0_77_712 ();
 sg13g2_decap_8 FILLER_0_77_719 ();
 sg13g2_decap_8 FILLER_0_77_726 ();
 sg13g2_decap_8 FILLER_0_77_737 ();
 sg13g2_fill_2 FILLER_0_77_744 ();
 sg13g2_decap_8 FILLER_0_77_782 ();
 sg13g2_decap_8 FILLER_0_77_789 ();
 sg13g2_decap_8 FILLER_0_77_796 ();
 sg13g2_decap_8 FILLER_0_77_803 ();
 sg13g2_fill_2 FILLER_0_77_810 ();
 sg13g2_fill_1 FILLER_0_77_812 ();
 sg13g2_decap_8 FILLER_0_77_843 ();
 sg13g2_decap_4 FILLER_0_77_850 ();
 sg13g2_fill_2 FILLER_0_77_854 ();
 sg13g2_fill_1 FILLER_0_77_905 ();
 sg13g2_fill_2 FILLER_0_77_934 ();
 sg13g2_fill_1 FILLER_0_77_956 ();
 sg13g2_decap_4 FILLER_0_77_961 ();
 sg13g2_decap_8 FILLER_0_77_972 ();
 sg13g2_fill_1 FILLER_0_77_979 ();
 sg13g2_decap_8 FILLER_0_77_984 ();
 sg13g2_decap_8 FILLER_0_77_991 ();
 sg13g2_decap_8 FILLER_0_77_998 ();
 sg13g2_decap_4 FILLER_0_77_1005 ();
 sg13g2_fill_1 FILLER_0_77_1009 ();
 sg13g2_fill_1 FILLER_0_77_1023 ();
 sg13g2_decap_8 FILLER_0_77_1038 ();
 sg13g2_decap_8 FILLER_0_77_1045 ();
 sg13g2_decap_8 FILLER_0_77_1052 ();
 sg13g2_decap_8 FILLER_0_77_1059 ();
 sg13g2_decap_8 FILLER_0_77_1066 ();
 sg13g2_decap_8 FILLER_0_77_1073 ();
 sg13g2_decap_8 FILLER_0_77_1080 ();
 sg13g2_decap_8 FILLER_0_77_1087 ();
 sg13g2_decap_8 FILLER_0_77_1094 ();
 sg13g2_decap_8 FILLER_0_77_1101 ();
 sg13g2_decap_8 FILLER_0_77_1108 ();
 sg13g2_decap_8 FILLER_0_77_1115 ();
 sg13g2_decap_8 FILLER_0_77_1122 ();
 sg13g2_decap_8 FILLER_0_77_1129 ();
 sg13g2_decap_8 FILLER_0_77_1136 ();
 sg13g2_decap_8 FILLER_0_77_1143 ();
 sg13g2_decap_8 FILLER_0_77_1150 ();
 sg13g2_decap_8 FILLER_0_77_1157 ();
 sg13g2_decap_8 FILLER_0_77_1164 ();
 sg13g2_decap_8 FILLER_0_77_1171 ();
 sg13g2_decap_8 FILLER_0_77_1178 ();
 sg13g2_decap_8 FILLER_0_77_1185 ();
 sg13g2_decap_8 FILLER_0_77_1192 ();
 sg13g2_decap_8 FILLER_0_77_1199 ();
 sg13g2_decap_8 FILLER_0_77_1206 ();
 sg13g2_decap_8 FILLER_0_77_1213 ();
 sg13g2_decap_8 FILLER_0_77_1220 ();
 sg13g2_fill_1 FILLER_0_77_1227 ();
 sg13g2_decap_8 FILLER_0_78_0 ();
 sg13g2_decap_8 FILLER_0_78_7 ();
 sg13g2_decap_8 FILLER_0_78_14 ();
 sg13g2_decap_8 FILLER_0_78_21 ();
 sg13g2_decap_8 FILLER_0_78_28 ();
 sg13g2_decap_8 FILLER_0_78_35 ();
 sg13g2_decap_8 FILLER_0_78_42 ();
 sg13g2_decap_8 FILLER_0_78_49 ();
 sg13g2_decap_4 FILLER_0_78_56 ();
 sg13g2_fill_1 FILLER_0_78_60 ();
 sg13g2_fill_2 FILLER_0_78_78 ();
 sg13g2_fill_1 FILLER_0_78_80 ();
 sg13g2_fill_2 FILLER_0_78_125 ();
 sg13g2_fill_1 FILLER_0_78_127 ();
 sg13g2_fill_1 FILLER_0_78_148 ();
 sg13g2_fill_1 FILLER_0_78_175 ();
 sg13g2_fill_1 FILLER_0_78_181 ();
 sg13g2_fill_1 FILLER_0_78_208 ();
 sg13g2_fill_1 FILLER_0_78_214 ();
 sg13g2_decap_8 FILLER_0_78_229 ();
 sg13g2_decap_4 FILLER_0_78_236 ();
 sg13g2_fill_1 FILLER_0_78_240 ();
 sg13g2_decap_8 FILLER_0_78_264 ();
 sg13g2_decap_8 FILLER_0_78_271 ();
 sg13g2_decap_8 FILLER_0_78_278 ();
 sg13g2_decap_8 FILLER_0_78_285 ();
 sg13g2_decap_8 FILLER_0_78_292 ();
 sg13g2_decap_8 FILLER_0_78_299 ();
 sg13g2_decap_8 FILLER_0_78_306 ();
 sg13g2_fill_2 FILLER_0_78_313 ();
 sg13g2_fill_1 FILLER_0_78_315 ();
 sg13g2_fill_1 FILLER_0_78_320 ();
 sg13g2_fill_2 FILLER_0_78_383 ();
 sg13g2_decap_8 FILLER_0_78_389 ();
 sg13g2_decap_8 FILLER_0_78_396 ();
 sg13g2_decap_8 FILLER_0_78_403 ();
 sg13g2_decap_8 FILLER_0_78_410 ();
 sg13g2_decap_8 FILLER_0_78_417 ();
 sg13g2_fill_2 FILLER_0_78_424 ();
 sg13g2_fill_2 FILLER_0_78_457 ();
 sg13g2_fill_1 FILLER_0_78_463 ();
 sg13g2_fill_1 FILLER_0_78_520 ();
 sg13g2_fill_2 FILLER_0_78_526 ();
 sg13g2_fill_2 FILLER_0_78_532 ();
 sg13g2_decap_4 FILLER_0_78_544 ();
 sg13g2_fill_2 FILLER_0_78_548 ();
 sg13g2_decap_8 FILLER_0_78_576 ();
 sg13g2_decap_8 FILLER_0_78_583 ();
 sg13g2_fill_2 FILLER_0_78_590 ();
 sg13g2_fill_1 FILLER_0_78_592 ();
 sg13g2_decap_8 FILLER_0_78_663 ();
 sg13g2_decap_8 FILLER_0_78_670 ();
 sg13g2_decap_8 FILLER_0_78_677 ();
 sg13g2_decap_8 FILLER_0_78_715 ();
 sg13g2_decap_8 FILLER_0_78_722 ();
 sg13g2_decap_8 FILLER_0_78_729 ();
 sg13g2_decap_8 FILLER_0_78_736 ();
 sg13g2_decap_8 FILLER_0_78_743 ();
 sg13g2_fill_1 FILLER_0_78_750 ();
 sg13g2_decap_8 FILLER_0_78_795 ();
 sg13g2_decap_8 FILLER_0_78_802 ();
 sg13g2_decap_4 FILLER_0_78_809 ();
 sg13g2_fill_2 FILLER_0_78_813 ();
 sg13g2_fill_1 FILLER_0_78_824 ();
 sg13g2_decap_4 FILLER_0_78_835 ();
 sg13g2_fill_1 FILLER_0_78_839 ();
 sg13g2_decap_8 FILLER_0_78_850 ();
 sg13g2_fill_2 FILLER_0_78_857 ();
 sg13g2_decap_8 FILLER_0_78_890 ();
 sg13g2_decap_8 FILLER_0_78_897 ();
 sg13g2_decap_8 FILLER_0_78_904 ();
 sg13g2_decap_8 FILLER_0_78_911 ();
 sg13g2_decap_8 FILLER_0_78_918 ();
 sg13g2_decap_8 FILLER_0_78_930 ();
 sg13g2_decap_8 FILLER_0_78_937 ();
 sg13g2_decap_8 FILLER_0_78_944 ();
 sg13g2_decap_4 FILLER_0_78_951 ();
 sg13g2_decap_4 FILLER_0_78_978 ();
 sg13g2_fill_2 FILLER_0_78_982 ();
 sg13g2_decap_8 FILLER_0_78_988 ();
 sg13g2_decap_8 FILLER_0_78_995 ();
 sg13g2_fill_2 FILLER_0_78_1002 ();
 sg13g2_fill_2 FILLER_0_78_1012 ();
 sg13g2_decap_8 FILLER_0_78_1040 ();
 sg13g2_decap_8 FILLER_0_78_1047 ();
 sg13g2_decap_8 FILLER_0_78_1054 ();
 sg13g2_decap_8 FILLER_0_78_1061 ();
 sg13g2_decap_8 FILLER_0_78_1068 ();
 sg13g2_decap_8 FILLER_0_78_1075 ();
 sg13g2_decap_8 FILLER_0_78_1082 ();
 sg13g2_decap_8 FILLER_0_78_1089 ();
 sg13g2_decap_8 FILLER_0_78_1096 ();
 sg13g2_decap_8 FILLER_0_78_1103 ();
 sg13g2_decap_8 FILLER_0_78_1110 ();
 sg13g2_decap_8 FILLER_0_78_1117 ();
 sg13g2_decap_8 FILLER_0_78_1124 ();
 sg13g2_decap_8 FILLER_0_78_1131 ();
 sg13g2_decap_8 FILLER_0_78_1138 ();
 sg13g2_decap_8 FILLER_0_78_1145 ();
 sg13g2_decap_8 FILLER_0_78_1152 ();
 sg13g2_decap_8 FILLER_0_78_1159 ();
 sg13g2_decap_8 FILLER_0_78_1166 ();
 sg13g2_decap_8 FILLER_0_78_1173 ();
 sg13g2_decap_8 FILLER_0_78_1180 ();
 sg13g2_decap_8 FILLER_0_78_1187 ();
 sg13g2_decap_8 FILLER_0_78_1194 ();
 sg13g2_decap_8 FILLER_0_78_1201 ();
 sg13g2_decap_8 FILLER_0_78_1208 ();
 sg13g2_decap_8 FILLER_0_78_1215 ();
 sg13g2_decap_4 FILLER_0_78_1222 ();
 sg13g2_fill_2 FILLER_0_78_1226 ();
 sg13g2_decap_8 FILLER_0_79_0 ();
 sg13g2_decap_8 FILLER_0_79_7 ();
 sg13g2_fill_2 FILLER_0_79_14 ();
 sg13g2_fill_1 FILLER_0_79_16 ();
 sg13g2_fill_2 FILLER_0_79_22 ();
 sg13g2_fill_1 FILLER_0_79_75 ();
 sg13g2_decap_8 FILLER_0_79_80 ();
 sg13g2_decap_8 FILLER_0_79_87 ();
 sg13g2_decap_8 FILLER_0_79_94 ();
 sg13g2_decap_4 FILLER_0_79_101 ();
 sg13g2_fill_1 FILLER_0_79_105 ();
 sg13g2_decap_4 FILLER_0_79_111 ();
 sg13g2_fill_1 FILLER_0_79_115 ();
 sg13g2_decap_8 FILLER_0_79_125 ();
 sg13g2_decap_8 FILLER_0_79_132 ();
 sg13g2_decap_4 FILLER_0_79_139 ();
 sg13g2_fill_2 FILLER_0_79_156 ();
 sg13g2_fill_2 FILLER_0_79_196 ();
 sg13g2_decap_8 FILLER_0_79_206 ();
 sg13g2_fill_2 FILLER_0_79_213 ();
 sg13g2_fill_1 FILLER_0_79_215 ();
 sg13g2_fill_2 FILLER_0_79_242 ();
 sg13g2_decap_8 FILLER_0_79_273 ();
 sg13g2_decap_8 FILLER_0_79_280 ();
 sg13g2_decap_8 FILLER_0_79_287 ();
 sg13g2_decap_8 FILLER_0_79_294 ();
 sg13g2_decap_4 FILLER_0_79_301 ();
 sg13g2_fill_1 FILLER_0_79_336 ();
 sg13g2_decap_8 FILLER_0_79_397 ();
 sg13g2_fill_2 FILLER_0_79_409 ();
 sg13g2_decap_8 FILLER_0_79_421 ();
 sg13g2_fill_2 FILLER_0_79_428 ();
 sg13g2_decap_4 FILLER_0_79_460 ();
 sg13g2_fill_2 FILLER_0_79_464 ();
 sg13g2_fill_2 FILLER_0_79_492 ();
 sg13g2_fill_1 FILLER_0_79_494 ();
 sg13g2_fill_2 FILLER_0_79_509 ();
 sg13g2_fill_1 FILLER_0_79_511 ();
 sg13g2_decap_8 FILLER_0_79_520 ();
 sg13g2_decap_8 FILLER_0_79_527 ();
 sg13g2_decap_8 FILLER_0_79_534 ();
 sg13g2_fill_2 FILLER_0_79_541 ();
 sg13g2_fill_1 FILLER_0_79_543 ();
 sg13g2_decap_4 FILLER_0_79_549 ();
 sg13g2_fill_1 FILLER_0_79_553 ();
 sg13g2_decap_4 FILLER_0_79_562 ();
 sg13g2_fill_2 FILLER_0_79_566 ();
 sg13g2_decap_8 FILLER_0_79_578 ();
 sg13g2_decap_8 FILLER_0_79_585 ();
 sg13g2_decap_8 FILLER_0_79_592 ();
 sg13g2_fill_2 FILLER_0_79_599 ();
 sg13g2_fill_1 FILLER_0_79_605 ();
 sg13g2_fill_2 FILLER_0_79_680 ();
 sg13g2_fill_1 FILLER_0_79_682 ();
 sg13g2_fill_1 FILLER_0_79_693 ();
 sg13g2_fill_2 FILLER_0_79_704 ();
 sg13g2_decap_8 FILLER_0_79_710 ();
 sg13g2_decap_8 FILLER_0_79_729 ();
 sg13g2_decap_8 FILLER_0_79_736 ();
 sg13g2_decap_8 FILLER_0_79_743 ();
 sg13g2_decap_8 FILLER_0_79_750 ();
 sg13g2_decap_4 FILLER_0_79_757 ();
 sg13g2_decap_8 FILLER_0_79_806 ();
 sg13g2_fill_1 FILLER_0_79_817 ();
 sg13g2_decap_8 FILLER_0_79_849 ();
 sg13g2_decap_8 FILLER_0_79_856 ();
 sg13g2_decap_4 FILLER_0_79_863 ();
 sg13g2_fill_2 FILLER_0_79_871 ();
 sg13g2_fill_1 FILLER_0_79_873 ();
 sg13g2_decap_4 FILLER_0_79_877 ();
 sg13g2_fill_1 FILLER_0_79_881 ();
 sg13g2_decap_8 FILLER_0_79_892 ();
 sg13g2_decap_4 FILLER_0_79_899 ();
 sg13g2_fill_2 FILLER_0_79_903 ();
 sg13g2_decap_8 FILLER_0_79_910 ();
 sg13g2_fill_2 FILLER_0_79_917 ();
 sg13g2_fill_1 FILLER_0_79_919 ();
 sg13g2_fill_2 FILLER_0_79_964 ();
 sg13g2_fill_1 FILLER_0_79_976 ();
 sg13g2_decap_8 FILLER_0_79_1044 ();
 sg13g2_decap_8 FILLER_0_79_1051 ();
 sg13g2_decap_8 FILLER_0_79_1058 ();
 sg13g2_decap_8 FILLER_0_79_1065 ();
 sg13g2_decap_8 FILLER_0_79_1072 ();
 sg13g2_decap_8 FILLER_0_79_1079 ();
 sg13g2_decap_8 FILLER_0_79_1086 ();
 sg13g2_decap_8 FILLER_0_79_1093 ();
 sg13g2_decap_8 FILLER_0_79_1100 ();
 sg13g2_decap_8 FILLER_0_79_1107 ();
 sg13g2_decap_8 FILLER_0_79_1114 ();
 sg13g2_decap_8 FILLER_0_79_1121 ();
 sg13g2_decap_8 FILLER_0_79_1128 ();
 sg13g2_decap_8 FILLER_0_79_1135 ();
 sg13g2_decap_8 FILLER_0_79_1142 ();
 sg13g2_decap_8 FILLER_0_79_1149 ();
 sg13g2_decap_8 FILLER_0_79_1156 ();
 sg13g2_decap_8 FILLER_0_79_1163 ();
 sg13g2_decap_8 FILLER_0_79_1170 ();
 sg13g2_decap_8 FILLER_0_79_1177 ();
 sg13g2_decap_8 FILLER_0_79_1184 ();
 sg13g2_decap_8 FILLER_0_79_1191 ();
 sg13g2_decap_8 FILLER_0_79_1198 ();
 sg13g2_decap_8 FILLER_0_79_1205 ();
 sg13g2_decap_8 FILLER_0_79_1212 ();
 sg13g2_decap_8 FILLER_0_79_1219 ();
 sg13g2_fill_2 FILLER_0_79_1226 ();
 sg13g2_decap_8 FILLER_0_80_0 ();
 sg13g2_fill_2 FILLER_0_80_7 ();
 sg13g2_decap_8 FILLER_0_80_13 ();
 sg13g2_fill_2 FILLER_0_80_20 ();
 sg13g2_fill_1 FILLER_0_80_22 ();
 sg13g2_decap_8 FILLER_0_80_89 ();
 sg13g2_decap_8 FILLER_0_80_96 ();
 sg13g2_decap_8 FILLER_0_80_138 ();
 sg13g2_decap_4 FILLER_0_80_145 ();
 sg13g2_fill_2 FILLER_0_80_149 ();
 sg13g2_decap_8 FILLER_0_80_155 ();
 sg13g2_decap_8 FILLER_0_80_162 ();
 sg13g2_decap_4 FILLER_0_80_169 ();
 sg13g2_fill_2 FILLER_0_80_213 ();
 sg13g2_fill_1 FILLER_0_80_235 ();
 sg13g2_decap_8 FILLER_0_80_246 ();
 sg13g2_decap_8 FILLER_0_80_253 ();
 sg13g2_decap_8 FILLER_0_80_260 ();
 sg13g2_decap_4 FILLER_0_80_267 ();
 sg13g2_decap_8 FILLER_0_80_275 ();
 sg13g2_decap_8 FILLER_0_80_282 ();
 sg13g2_decap_8 FILLER_0_80_289 ();
 sg13g2_decap_8 FILLER_0_80_296 ();
 sg13g2_decap_4 FILLER_0_80_303 ();
 sg13g2_fill_2 FILLER_0_80_307 ();
 sg13g2_fill_1 FILLER_0_80_322 ();
 sg13g2_decap_4 FILLER_0_80_343 ();
 sg13g2_decap_8 FILLER_0_80_355 ();
 sg13g2_fill_1 FILLER_0_80_362 ();
 sg13g2_decap_8 FILLER_0_80_367 ();
 sg13g2_decap_8 FILLER_0_80_374 ();
 sg13g2_decap_8 FILLER_0_80_381 ();
 sg13g2_decap_4 FILLER_0_80_432 ();
 sg13g2_fill_1 FILLER_0_80_436 ();
 sg13g2_fill_1 FILLER_0_80_442 ();
 sg13g2_decap_4 FILLER_0_80_457 ();
 sg13g2_fill_2 FILLER_0_80_461 ();
 sg13g2_fill_2 FILLER_0_80_471 ();
 sg13g2_fill_1 FILLER_0_80_473 ();
 sg13g2_decap_4 FILLER_0_80_478 ();
 sg13g2_fill_1 FILLER_0_80_482 ();
 sg13g2_decap_8 FILLER_0_80_488 ();
 sg13g2_decap_8 FILLER_0_80_495 ();
 sg13g2_decap_8 FILLER_0_80_502 ();
 sg13g2_decap_8 FILLER_0_80_509 ();
 sg13g2_decap_8 FILLER_0_80_516 ();
 sg13g2_decap_8 FILLER_0_80_523 ();
 sg13g2_decap_4 FILLER_0_80_530 ();
 sg13g2_fill_1 FILLER_0_80_534 ();
 sg13g2_decap_8 FILLER_0_80_573 ();
 sg13g2_decap_8 FILLER_0_80_580 ();
 sg13g2_decap_8 FILLER_0_80_587 ();
 sg13g2_decap_8 FILLER_0_80_594 ();
 sg13g2_decap_8 FILLER_0_80_601 ();
 sg13g2_decap_8 FILLER_0_80_608 ();
 sg13g2_decap_8 FILLER_0_80_615 ();
 sg13g2_fill_1 FILLER_0_80_637 ();
 sg13g2_decap_8 FILLER_0_80_735 ();
 sg13g2_decap_8 FILLER_0_80_742 ();
 sg13g2_decap_8 FILLER_0_80_749 ();
 sg13g2_decap_8 FILLER_0_80_756 ();
 sg13g2_decap_8 FILLER_0_80_763 ();
 sg13g2_fill_1 FILLER_0_80_770 ();
 sg13g2_fill_2 FILLER_0_80_800 ();
 sg13g2_fill_2 FILLER_0_80_832 ();
 sg13g2_fill_1 FILLER_0_80_834 ();
 sg13g2_fill_2 FILLER_0_80_845 ();
 sg13g2_decap_8 FILLER_0_80_851 ();
 sg13g2_decap_4 FILLER_0_80_858 ();
 sg13g2_fill_1 FILLER_0_80_862 ();
 sg13g2_fill_1 FILLER_0_80_924 ();
 sg13g2_fill_2 FILLER_0_80_987 ();
 sg13g2_fill_2 FILLER_0_80_1015 ();
 sg13g2_decap_8 FILLER_0_80_1043 ();
 sg13g2_decap_8 FILLER_0_80_1050 ();
 sg13g2_decap_8 FILLER_0_80_1057 ();
 sg13g2_decap_8 FILLER_0_80_1064 ();
 sg13g2_decap_8 FILLER_0_80_1071 ();
 sg13g2_decap_8 FILLER_0_80_1078 ();
 sg13g2_decap_8 FILLER_0_80_1085 ();
 sg13g2_decap_8 FILLER_0_80_1092 ();
 sg13g2_decap_8 FILLER_0_80_1099 ();
 sg13g2_decap_8 FILLER_0_80_1106 ();
 sg13g2_decap_8 FILLER_0_80_1113 ();
 sg13g2_decap_8 FILLER_0_80_1120 ();
 sg13g2_decap_8 FILLER_0_80_1127 ();
 sg13g2_decap_8 FILLER_0_80_1134 ();
 sg13g2_decap_8 FILLER_0_80_1141 ();
 sg13g2_decap_8 FILLER_0_80_1148 ();
 sg13g2_decap_8 FILLER_0_80_1155 ();
 sg13g2_decap_8 FILLER_0_80_1162 ();
 sg13g2_decap_8 FILLER_0_80_1169 ();
 sg13g2_decap_8 FILLER_0_80_1176 ();
 sg13g2_decap_8 FILLER_0_80_1183 ();
 sg13g2_decap_8 FILLER_0_80_1190 ();
 sg13g2_decap_8 FILLER_0_80_1197 ();
 sg13g2_decap_8 FILLER_0_80_1204 ();
 sg13g2_decap_8 FILLER_0_80_1211 ();
 sg13g2_decap_8 FILLER_0_80_1218 ();
 sg13g2_fill_2 FILLER_0_80_1225 ();
 sg13g2_fill_1 FILLER_0_80_1227 ();
 sg13g2_decap_8 FILLER_0_81_0 ();
 sg13g2_fill_1 FILLER_0_81_16 ();
 sg13g2_fill_2 FILLER_0_81_27 ();
 sg13g2_fill_2 FILLER_0_81_91 ();
 sg13g2_fill_1 FILLER_0_81_93 ();
 sg13g2_decap_8 FILLER_0_81_118 ();
 sg13g2_decap_8 FILLER_0_81_125 ();
 sg13g2_decap_8 FILLER_0_81_132 ();
 sg13g2_decap_8 FILLER_0_81_139 ();
 sg13g2_decap_8 FILLER_0_81_146 ();
 sg13g2_decap_4 FILLER_0_81_153 ();
 sg13g2_fill_2 FILLER_0_81_157 ();
 sg13g2_decap_4 FILLER_0_81_163 ();
 sg13g2_fill_2 FILLER_0_81_167 ();
 sg13g2_fill_1 FILLER_0_81_257 ();
 sg13g2_fill_2 FILLER_0_81_263 ();
 sg13g2_decap_8 FILLER_0_81_291 ();
 sg13g2_decap_8 FILLER_0_81_298 ();
 sg13g2_decap_8 FILLER_0_81_342 ();
 sg13g2_decap_8 FILLER_0_81_349 ();
 sg13g2_decap_8 FILLER_0_81_356 ();
 sg13g2_fill_2 FILLER_0_81_363 ();
 sg13g2_fill_1 FILLER_0_81_365 ();
 sg13g2_fill_2 FILLER_0_81_392 ();
 sg13g2_fill_1 FILLER_0_81_394 ();
 sg13g2_fill_1 FILLER_0_81_400 ();
 sg13g2_fill_2 FILLER_0_81_411 ();
 sg13g2_fill_1 FILLER_0_81_413 ();
 sg13g2_decap_8 FILLER_0_81_418 ();
 sg13g2_decap_8 FILLER_0_81_425 ();
 sg13g2_decap_8 FILLER_0_81_432 ();
 sg13g2_decap_8 FILLER_0_81_439 ();
 sg13g2_fill_2 FILLER_0_81_446 ();
 sg13g2_decap_8 FILLER_0_81_458 ();
 sg13g2_decap_4 FILLER_0_81_465 ();
 sg13g2_fill_2 FILLER_0_81_469 ();
 sg13g2_fill_1 FILLER_0_81_502 ();
 sg13g2_decap_8 FILLER_0_81_534 ();
 sg13g2_decap_8 FILLER_0_81_541 ();
 sg13g2_fill_2 FILLER_0_81_548 ();
 sg13g2_decap_8 FILLER_0_81_569 ();
 sg13g2_decap_8 FILLER_0_81_576 ();
 sg13g2_decap_8 FILLER_0_81_583 ();
 sg13g2_fill_1 FILLER_0_81_590 ();
 sg13g2_decap_8 FILLER_0_81_595 ();
 sg13g2_decap_8 FILLER_0_81_602 ();
 sg13g2_decap_8 FILLER_0_81_609 ();
 sg13g2_fill_2 FILLER_0_81_616 ();
 sg13g2_decap_8 FILLER_0_81_623 ();
 sg13g2_decap_8 FILLER_0_81_630 ();
 sg13g2_fill_2 FILLER_0_81_637 ();
 sg13g2_fill_1 FILLER_0_81_639 ();
 sg13g2_fill_1 FILLER_0_81_644 ();
 sg13g2_fill_2 FILLER_0_81_660 ();
 sg13g2_fill_1 FILLER_0_81_662 ();
 sg13g2_fill_2 FILLER_0_81_667 ();
 sg13g2_decap_4 FILLER_0_81_679 ();
 sg13g2_fill_2 FILLER_0_81_688 ();
 sg13g2_decap_4 FILLER_0_81_694 ();
 sg13g2_fill_2 FILLER_0_81_708 ();
 sg13g2_fill_1 FILLER_0_81_710 ();
 sg13g2_decap_8 FILLER_0_81_724 ();
 sg13g2_decap_8 FILLER_0_81_735 ();
 sg13g2_decap_8 FILLER_0_81_746 ();
 sg13g2_decap_8 FILLER_0_81_753 ();
 sg13g2_decap_8 FILLER_0_81_760 ();
 sg13g2_decap_8 FILLER_0_81_767 ();
 sg13g2_decap_4 FILLER_0_81_774 ();
 sg13g2_fill_2 FILLER_0_81_778 ();
 sg13g2_decap_4 FILLER_0_81_788 ();
 sg13g2_fill_1 FILLER_0_81_792 ();
 sg13g2_decap_8 FILLER_0_81_861 ();
 sg13g2_fill_1 FILLER_0_81_868 ();
 sg13g2_decap_4 FILLER_0_81_904 ();
 sg13g2_fill_1 FILLER_0_81_934 ();
 sg13g2_fill_1 FILLER_0_81_949 ();
 sg13g2_fill_2 FILLER_0_81_981 ();
 sg13g2_fill_1 FILLER_0_81_983 ();
 sg13g2_fill_2 FILLER_0_81_999 ();
 sg13g2_fill_1 FILLER_0_81_1015 ();
 sg13g2_decap_8 FILLER_0_81_1021 ();
 sg13g2_decap_8 FILLER_0_81_1042 ();
 sg13g2_decap_8 FILLER_0_81_1049 ();
 sg13g2_decap_8 FILLER_0_81_1056 ();
 sg13g2_decap_8 FILLER_0_81_1063 ();
 sg13g2_decap_8 FILLER_0_81_1070 ();
 sg13g2_decap_8 FILLER_0_81_1077 ();
 sg13g2_decap_8 FILLER_0_81_1084 ();
 sg13g2_decap_8 FILLER_0_81_1091 ();
 sg13g2_decap_8 FILLER_0_81_1098 ();
 sg13g2_decap_8 FILLER_0_81_1105 ();
 sg13g2_decap_8 FILLER_0_81_1112 ();
 sg13g2_decap_8 FILLER_0_81_1119 ();
 sg13g2_decap_8 FILLER_0_81_1126 ();
 sg13g2_decap_8 FILLER_0_81_1133 ();
 sg13g2_decap_8 FILLER_0_81_1140 ();
 sg13g2_decap_8 FILLER_0_81_1147 ();
 sg13g2_decap_8 FILLER_0_81_1154 ();
 sg13g2_decap_8 FILLER_0_81_1161 ();
 sg13g2_decap_8 FILLER_0_81_1168 ();
 sg13g2_decap_8 FILLER_0_81_1175 ();
 sg13g2_decap_8 FILLER_0_81_1182 ();
 sg13g2_decap_8 FILLER_0_81_1189 ();
 sg13g2_decap_8 FILLER_0_81_1196 ();
 sg13g2_decap_8 FILLER_0_81_1203 ();
 sg13g2_decap_8 FILLER_0_81_1210 ();
 sg13g2_decap_8 FILLER_0_81_1217 ();
 sg13g2_decap_4 FILLER_0_81_1224 ();
 sg13g2_decap_8 FILLER_0_82_0 ();
 sg13g2_fill_1 FILLER_0_82_37 ();
 sg13g2_decap_8 FILLER_0_82_42 ();
 sg13g2_decap_8 FILLER_0_82_49 ();
 sg13g2_decap_8 FILLER_0_82_56 ();
 sg13g2_decap_8 FILLER_0_82_88 ();
 sg13g2_fill_2 FILLER_0_82_95 ();
 sg13g2_decap_8 FILLER_0_82_128 ();
 sg13g2_decap_8 FILLER_0_82_135 ();
 sg13g2_decap_4 FILLER_0_82_142 ();
 sg13g2_fill_1 FILLER_0_82_146 ();
 sg13g2_fill_2 FILLER_0_82_248 ();
 sg13g2_decap_8 FILLER_0_82_260 ();
 sg13g2_decap_8 FILLER_0_82_267 ();
 sg13g2_decap_8 FILLER_0_82_274 ();
 sg13g2_decap_8 FILLER_0_82_281 ();
 sg13g2_decap_8 FILLER_0_82_288 ();
 sg13g2_decap_8 FILLER_0_82_295 ();
 sg13g2_decap_8 FILLER_0_82_302 ();
 sg13g2_fill_2 FILLER_0_82_309 ();
 sg13g2_decap_8 FILLER_0_82_345 ();
 sg13g2_decap_8 FILLER_0_82_352 ();
 sg13g2_fill_1 FILLER_0_82_359 ();
 sg13g2_fill_2 FILLER_0_82_400 ();
 sg13g2_fill_1 FILLER_0_82_402 ();
 sg13g2_fill_2 FILLER_0_82_434 ();
 sg13g2_fill_1 FILLER_0_82_436 ();
 sg13g2_fill_1 FILLER_0_82_463 ();
 sg13g2_decap_4 FILLER_0_82_479 ();
 sg13g2_fill_2 FILLER_0_82_483 ();
 sg13g2_fill_2 FILLER_0_82_546 ();
 sg13g2_decap_4 FILLER_0_82_605 ();
 sg13g2_decap_8 FILLER_0_82_661 ();
 sg13g2_decap_8 FILLER_0_82_668 ();
 sg13g2_decap_8 FILLER_0_82_675 ();
 sg13g2_decap_8 FILLER_0_82_682 ();
 sg13g2_decap_4 FILLER_0_82_689 ();
 sg13g2_fill_1 FILLER_0_82_693 ();
 sg13g2_fill_2 FILLER_0_82_704 ();
 sg13g2_decap_4 FILLER_0_82_711 ();
 sg13g2_decap_4 FILLER_0_82_720 ();
 sg13g2_decap_4 FILLER_0_82_750 ();
 sg13g2_fill_1 FILLER_0_82_754 ();
 sg13g2_decap_8 FILLER_0_82_760 ();
 sg13g2_decap_8 FILLER_0_82_767 ();
 sg13g2_decap_8 FILLER_0_82_774 ();
 sg13g2_decap_4 FILLER_0_82_781 ();
 sg13g2_fill_1 FILLER_0_82_785 ();
 sg13g2_fill_1 FILLER_0_82_816 ();
 sg13g2_fill_2 FILLER_0_82_822 ();
 sg13g2_fill_2 FILLER_0_82_829 ();
 sg13g2_fill_2 FILLER_0_82_835 ();
 sg13g2_decap_8 FILLER_0_82_863 ();
 sg13g2_fill_2 FILLER_0_82_870 ();
 sg13g2_fill_1 FILLER_0_82_872 ();
 sg13g2_fill_2 FILLER_0_82_902 ();
 sg13g2_fill_1 FILLER_0_82_904 ();
 sg13g2_decap_4 FILLER_0_82_919 ();
 sg13g2_decap_8 FILLER_0_82_933 ();
 sg13g2_decap_8 FILLER_0_82_944 ();
 sg13g2_decap_8 FILLER_0_82_951 ();
 sg13g2_fill_2 FILLER_0_82_958 ();
 sg13g2_fill_1 FILLER_0_82_960 ();
 sg13g2_decap_4 FILLER_0_82_965 ();
 sg13g2_decap_8 FILLER_0_82_973 ();
 sg13g2_fill_2 FILLER_0_82_980 ();
 sg13g2_decap_8 FILLER_0_82_987 ();
 sg13g2_fill_2 FILLER_0_82_994 ();
 sg13g2_decap_8 FILLER_0_82_1000 ();
 sg13g2_decap_8 FILLER_0_82_1007 ();
 sg13g2_decap_8 FILLER_0_82_1014 ();
 sg13g2_decap_8 FILLER_0_82_1021 ();
 sg13g2_decap_8 FILLER_0_82_1028 ();
 sg13g2_decap_8 FILLER_0_82_1035 ();
 sg13g2_decap_8 FILLER_0_82_1042 ();
 sg13g2_decap_8 FILLER_0_82_1049 ();
 sg13g2_decap_8 FILLER_0_82_1056 ();
 sg13g2_decap_8 FILLER_0_82_1063 ();
 sg13g2_decap_8 FILLER_0_82_1070 ();
 sg13g2_decap_8 FILLER_0_82_1077 ();
 sg13g2_decap_8 FILLER_0_82_1084 ();
 sg13g2_decap_8 FILLER_0_82_1091 ();
 sg13g2_decap_8 FILLER_0_82_1098 ();
 sg13g2_decap_8 FILLER_0_82_1105 ();
 sg13g2_decap_8 FILLER_0_82_1112 ();
 sg13g2_decap_8 FILLER_0_82_1119 ();
 sg13g2_decap_8 FILLER_0_82_1126 ();
 sg13g2_decap_8 FILLER_0_82_1133 ();
 sg13g2_decap_8 FILLER_0_82_1140 ();
 sg13g2_decap_8 FILLER_0_82_1147 ();
 sg13g2_decap_8 FILLER_0_82_1154 ();
 sg13g2_decap_8 FILLER_0_82_1161 ();
 sg13g2_decap_8 FILLER_0_82_1168 ();
 sg13g2_decap_8 FILLER_0_82_1175 ();
 sg13g2_decap_8 FILLER_0_82_1182 ();
 sg13g2_decap_8 FILLER_0_82_1189 ();
 sg13g2_decap_8 FILLER_0_82_1196 ();
 sg13g2_decap_8 FILLER_0_82_1203 ();
 sg13g2_decap_8 FILLER_0_82_1210 ();
 sg13g2_decap_8 FILLER_0_82_1217 ();
 sg13g2_decap_4 FILLER_0_82_1224 ();
 sg13g2_decap_8 FILLER_0_83_40 ();
 sg13g2_decap_8 FILLER_0_83_47 ();
 sg13g2_decap_8 FILLER_0_83_54 ();
 sg13g2_decap_8 FILLER_0_83_61 ();
 sg13g2_decap_4 FILLER_0_83_68 ();
 sg13g2_decap_8 FILLER_0_83_76 ();
 sg13g2_decap_8 FILLER_0_83_83 ();
 sg13g2_decap_4 FILLER_0_83_90 ();
 sg13g2_fill_1 FILLER_0_83_94 ();
 sg13g2_decap_4 FILLER_0_83_126 ();
 sg13g2_fill_1 FILLER_0_83_130 ();
 sg13g2_decap_4 FILLER_0_83_162 ();
 sg13g2_decap_8 FILLER_0_83_201 ();
 sg13g2_decap_8 FILLER_0_83_208 ();
 sg13g2_fill_2 FILLER_0_83_215 ();
 sg13g2_fill_1 FILLER_0_83_217 ();
 sg13g2_decap_8 FILLER_0_83_222 ();
 sg13g2_decap_8 FILLER_0_83_229 ();
 sg13g2_fill_1 FILLER_0_83_236 ();
 sg13g2_decap_8 FILLER_0_83_241 ();
 sg13g2_decap_8 FILLER_0_83_248 ();
 sg13g2_decap_8 FILLER_0_83_267 ();
 sg13g2_fill_2 FILLER_0_83_274 ();
 sg13g2_fill_1 FILLER_0_83_276 ();
 sg13g2_fill_1 FILLER_0_83_282 ();
 sg13g2_decap_8 FILLER_0_83_287 ();
 sg13g2_decap_8 FILLER_0_83_294 ();
 sg13g2_decap_8 FILLER_0_83_301 ();
 sg13g2_decap_8 FILLER_0_83_308 ();
 sg13g2_decap_4 FILLER_0_83_315 ();
 sg13g2_fill_2 FILLER_0_83_319 ();
 sg13g2_fill_2 FILLER_0_83_326 ();
 sg13g2_decap_8 FILLER_0_83_348 ();
 sg13g2_decap_8 FILLER_0_83_355 ();
 sg13g2_fill_2 FILLER_0_83_362 ();
 sg13g2_fill_1 FILLER_0_83_377 ();
 sg13g2_fill_1 FILLER_0_83_404 ();
 sg13g2_fill_1 FILLER_0_83_431 ();
 sg13g2_fill_2 FILLER_0_83_436 ();
 sg13g2_decap_4 FILLER_0_83_510 ();
 sg13g2_decap_4 FILLER_0_83_528 ();
 sg13g2_decap_4 FILLER_0_83_542 ();
 sg13g2_fill_2 FILLER_0_83_572 ();
 sg13g2_fill_1 FILLER_0_83_574 ();
 sg13g2_fill_1 FILLER_0_83_611 ();
 sg13g2_fill_2 FILLER_0_83_616 ();
 sg13g2_decap_4 FILLER_0_83_638 ();
 sg13g2_decap_8 FILLER_0_83_646 ();
 sg13g2_decap_8 FILLER_0_83_653 ();
 sg13g2_decap_4 FILLER_0_83_660 ();
 sg13g2_fill_1 FILLER_0_83_664 ();
 sg13g2_fill_1 FILLER_0_83_670 ();
 sg13g2_decap_8 FILLER_0_83_722 ();
 sg13g2_fill_2 FILLER_0_83_729 ();
 sg13g2_decap_4 FILLER_0_83_735 ();
 sg13g2_decap_8 FILLER_0_83_770 ();
 sg13g2_decap_8 FILLER_0_83_777 ();
 sg13g2_decap_8 FILLER_0_83_784 ();
 sg13g2_fill_1 FILLER_0_83_791 ();
 sg13g2_decap_8 FILLER_0_83_822 ();
 sg13g2_decap_8 FILLER_0_83_829 ();
 sg13g2_decap_4 FILLER_0_83_841 ();
 sg13g2_fill_1 FILLER_0_83_845 ();
 sg13g2_decap_8 FILLER_0_83_865 ();
 sg13g2_decap_8 FILLER_0_83_872 ();
 sg13g2_decap_4 FILLER_0_83_879 ();
 sg13g2_fill_1 FILLER_0_83_883 ();
 sg13g2_decap_8 FILLER_0_83_904 ();
 sg13g2_decap_8 FILLER_0_83_911 ();
 sg13g2_decap_8 FILLER_0_83_918 ();
 sg13g2_decap_8 FILLER_0_83_925 ();
 sg13g2_decap_8 FILLER_0_83_932 ();
 sg13g2_decap_8 FILLER_0_83_939 ();
 sg13g2_decap_8 FILLER_0_83_946 ();
 sg13g2_decap_8 FILLER_0_83_953 ();
 sg13g2_decap_8 FILLER_0_83_960 ();
 sg13g2_decap_8 FILLER_0_83_967 ();
 sg13g2_decap_8 FILLER_0_83_974 ();
 sg13g2_decap_8 FILLER_0_83_981 ();
 sg13g2_decap_8 FILLER_0_83_988 ();
 sg13g2_decap_8 FILLER_0_83_995 ();
 sg13g2_decap_8 FILLER_0_83_1002 ();
 sg13g2_decap_8 FILLER_0_83_1009 ();
 sg13g2_decap_8 FILLER_0_83_1016 ();
 sg13g2_decap_8 FILLER_0_83_1023 ();
 sg13g2_decap_8 FILLER_0_83_1030 ();
 sg13g2_decap_8 FILLER_0_83_1037 ();
 sg13g2_decap_8 FILLER_0_83_1044 ();
 sg13g2_decap_8 FILLER_0_83_1051 ();
 sg13g2_decap_8 FILLER_0_83_1058 ();
 sg13g2_decap_8 FILLER_0_83_1065 ();
 sg13g2_decap_8 FILLER_0_83_1072 ();
 sg13g2_decap_8 FILLER_0_83_1079 ();
 sg13g2_decap_8 FILLER_0_83_1086 ();
 sg13g2_decap_8 FILLER_0_83_1093 ();
 sg13g2_decap_8 FILLER_0_83_1100 ();
 sg13g2_decap_8 FILLER_0_83_1107 ();
 sg13g2_decap_8 FILLER_0_83_1114 ();
 sg13g2_decap_8 FILLER_0_83_1121 ();
 sg13g2_decap_8 FILLER_0_83_1128 ();
 sg13g2_decap_8 FILLER_0_83_1135 ();
 sg13g2_decap_8 FILLER_0_83_1142 ();
 sg13g2_decap_8 FILLER_0_83_1149 ();
 sg13g2_decap_8 FILLER_0_83_1156 ();
 sg13g2_decap_8 FILLER_0_83_1163 ();
 sg13g2_decap_8 FILLER_0_83_1170 ();
 sg13g2_decap_8 FILLER_0_83_1177 ();
 sg13g2_decap_8 FILLER_0_83_1184 ();
 sg13g2_decap_8 FILLER_0_83_1191 ();
 sg13g2_decap_8 FILLER_0_83_1198 ();
 sg13g2_decap_8 FILLER_0_83_1205 ();
 sg13g2_decap_8 FILLER_0_83_1212 ();
 sg13g2_decap_8 FILLER_0_83_1219 ();
 sg13g2_fill_2 FILLER_0_83_1226 ();
 sg13g2_decap_4 FILLER_0_84_0 ();
 sg13g2_fill_1 FILLER_0_84_4 ();
 sg13g2_decap_4 FILLER_0_84_27 ();
 sg13g2_decap_8 FILLER_0_84_41 ();
 sg13g2_decap_8 FILLER_0_84_48 ();
 sg13g2_decap_8 FILLER_0_84_55 ();
 sg13g2_decap_8 FILLER_0_84_62 ();
 sg13g2_decap_8 FILLER_0_84_69 ();
 sg13g2_decap_8 FILLER_0_84_76 ();
 sg13g2_fill_2 FILLER_0_84_83 ();
 sg13g2_decap_4 FILLER_0_84_121 ();
 sg13g2_decap_8 FILLER_0_84_135 ();
 sg13g2_fill_1 FILLER_0_84_142 ();
 sg13g2_decap_8 FILLER_0_84_147 ();
 sg13g2_fill_1 FILLER_0_84_154 ();
 sg13g2_fill_1 FILLER_0_84_165 ();
 sg13g2_decap_8 FILLER_0_84_181 ();
 sg13g2_decap_8 FILLER_0_84_188 ();
 sg13g2_decap_8 FILLER_0_84_195 ();
 sg13g2_decap_8 FILLER_0_84_202 ();
 sg13g2_decap_8 FILLER_0_84_209 ();
 sg13g2_decap_8 FILLER_0_84_216 ();
 sg13g2_decap_8 FILLER_0_84_223 ();
 sg13g2_decap_8 FILLER_0_84_230 ();
 sg13g2_decap_4 FILLER_0_84_237 ();
 sg13g2_fill_1 FILLER_0_84_241 ();
 sg13g2_fill_2 FILLER_0_84_257 ();
 sg13g2_fill_1 FILLER_0_84_259 ();
 sg13g2_fill_2 FILLER_0_84_264 ();
 sg13g2_decap_8 FILLER_0_84_302 ();
 sg13g2_decap_8 FILLER_0_84_309 ();
 sg13g2_fill_2 FILLER_0_84_321 ();
 sg13g2_fill_1 FILLER_0_84_323 ();
 sg13g2_decap_8 FILLER_0_84_355 ();
 sg13g2_decap_4 FILLER_0_84_362 ();
 sg13g2_fill_2 FILLER_0_84_366 ();
 sg13g2_decap_8 FILLER_0_84_373 ();
 sg13g2_fill_1 FILLER_0_84_399 ();
 sg13g2_decap_4 FILLER_0_84_436 ();
 sg13g2_fill_1 FILLER_0_84_444 ();
 sg13g2_fill_1 FILLER_0_84_450 ();
 sg13g2_fill_1 FILLER_0_84_471 ();
 sg13g2_fill_2 FILLER_0_84_477 ();
 sg13g2_fill_2 FILLER_0_84_483 ();
 sg13g2_fill_2 FILLER_0_84_489 ();
 sg13g2_fill_1 FILLER_0_84_491 ();
 sg13g2_decap_8 FILLER_0_84_496 ();
 sg13g2_decap_4 FILLER_0_84_503 ();
 sg13g2_fill_2 FILLER_0_84_507 ();
 sg13g2_decap_8 FILLER_0_84_514 ();
 sg13g2_decap_4 FILLER_0_84_521 ();
 sg13g2_decap_4 FILLER_0_84_544 ();
 sg13g2_decap_4 FILLER_0_84_557 ();
 sg13g2_fill_2 FILLER_0_84_561 ();
 sg13g2_fill_1 FILLER_0_84_573 ();
 sg13g2_fill_1 FILLER_0_84_582 ();
 sg13g2_decap_8 FILLER_0_84_587 ();
 sg13g2_decap_4 FILLER_0_84_599 ();
 sg13g2_decap_4 FILLER_0_84_613 ();
 sg13g2_fill_2 FILLER_0_84_617 ();
 sg13g2_fill_1 FILLER_0_84_624 ();
 sg13g2_fill_1 FILLER_0_84_635 ();
 sg13g2_decap_8 FILLER_0_84_641 ();
 sg13g2_fill_2 FILLER_0_84_648 ();
 sg13g2_fill_1 FILLER_0_84_650 ();
 sg13g2_decap_4 FILLER_0_84_716 ();
 sg13g2_decap_8 FILLER_0_84_787 ();
 sg13g2_fill_1 FILLER_0_84_794 ();
 sg13g2_decap_8 FILLER_0_84_800 ();
 sg13g2_decap_8 FILLER_0_84_825 ();
 sg13g2_decap_8 FILLER_0_84_832 ();
 sg13g2_fill_1 FILLER_0_84_839 ();
 sg13g2_decap_8 FILLER_0_84_881 ();
 sg13g2_fill_2 FILLER_0_84_888 ();
 sg13g2_decap_8 FILLER_0_84_894 ();
 sg13g2_decap_8 FILLER_0_84_901 ();
 sg13g2_decap_8 FILLER_0_84_908 ();
 sg13g2_decap_8 FILLER_0_84_915 ();
 sg13g2_decap_8 FILLER_0_84_922 ();
 sg13g2_decap_8 FILLER_0_84_929 ();
 sg13g2_decap_8 FILLER_0_84_936 ();
 sg13g2_decap_8 FILLER_0_84_943 ();
 sg13g2_decap_8 FILLER_0_84_950 ();
 sg13g2_decap_8 FILLER_0_84_957 ();
 sg13g2_decap_8 FILLER_0_84_964 ();
 sg13g2_decap_8 FILLER_0_84_971 ();
 sg13g2_decap_8 FILLER_0_84_978 ();
 sg13g2_decap_8 FILLER_0_84_985 ();
 sg13g2_decap_8 FILLER_0_84_992 ();
 sg13g2_decap_8 FILLER_0_84_999 ();
 sg13g2_decap_8 FILLER_0_84_1006 ();
 sg13g2_decap_8 FILLER_0_84_1013 ();
 sg13g2_decap_8 FILLER_0_84_1020 ();
 sg13g2_decap_8 FILLER_0_84_1027 ();
 sg13g2_decap_8 FILLER_0_84_1034 ();
 sg13g2_decap_8 FILLER_0_84_1041 ();
 sg13g2_decap_8 FILLER_0_84_1048 ();
 sg13g2_decap_8 FILLER_0_84_1055 ();
 sg13g2_decap_8 FILLER_0_84_1062 ();
 sg13g2_decap_8 FILLER_0_84_1069 ();
 sg13g2_decap_8 FILLER_0_84_1076 ();
 sg13g2_decap_8 FILLER_0_84_1083 ();
 sg13g2_decap_8 FILLER_0_84_1090 ();
 sg13g2_decap_8 FILLER_0_84_1097 ();
 sg13g2_decap_8 FILLER_0_84_1104 ();
 sg13g2_decap_8 FILLER_0_84_1111 ();
 sg13g2_decap_8 FILLER_0_84_1118 ();
 sg13g2_decap_8 FILLER_0_84_1125 ();
 sg13g2_decap_8 FILLER_0_84_1132 ();
 sg13g2_decap_8 FILLER_0_84_1139 ();
 sg13g2_decap_8 FILLER_0_84_1146 ();
 sg13g2_decap_8 FILLER_0_84_1153 ();
 sg13g2_decap_8 FILLER_0_84_1160 ();
 sg13g2_decap_8 FILLER_0_84_1167 ();
 sg13g2_decap_8 FILLER_0_84_1174 ();
 sg13g2_decap_8 FILLER_0_84_1181 ();
 sg13g2_decap_8 FILLER_0_84_1188 ();
 sg13g2_decap_8 FILLER_0_84_1195 ();
 sg13g2_decap_8 FILLER_0_84_1202 ();
 sg13g2_decap_8 FILLER_0_84_1209 ();
 sg13g2_decap_8 FILLER_0_84_1216 ();
 sg13g2_decap_4 FILLER_0_84_1223 ();
 sg13g2_fill_1 FILLER_0_84_1227 ();
 sg13g2_decap_8 FILLER_0_85_0 ();
 sg13g2_fill_1 FILLER_0_85_7 ();
 sg13g2_decap_8 FILLER_0_85_39 ();
 sg13g2_decap_8 FILLER_0_85_46 ();
 sg13g2_decap_8 FILLER_0_85_53 ();
 sg13g2_decap_8 FILLER_0_85_60 ();
 sg13g2_decap_4 FILLER_0_85_67 ();
 sg13g2_fill_1 FILLER_0_85_71 ();
 sg13g2_fill_2 FILLER_0_85_106 ();
 sg13g2_decap_8 FILLER_0_85_112 ();
 sg13g2_fill_2 FILLER_0_85_119 ();
 sg13g2_fill_1 FILLER_0_85_121 ();
 sg13g2_decap_8 FILLER_0_85_164 ();
 sg13g2_decap_8 FILLER_0_85_171 ();
 sg13g2_decap_8 FILLER_0_85_178 ();
 sg13g2_fill_2 FILLER_0_85_185 ();
 sg13g2_decap_8 FILLER_0_85_191 ();
 sg13g2_fill_1 FILLER_0_85_198 ();
 sg13g2_decap_8 FILLER_0_85_209 ();
 sg13g2_fill_2 FILLER_0_85_216 ();
 sg13g2_fill_2 FILLER_0_85_280 ();
 sg13g2_decap_4 FILLER_0_85_344 ();
 sg13g2_decap_8 FILLER_0_85_382 ();
 sg13g2_fill_2 FILLER_0_85_389 ();
 sg13g2_fill_1 FILLER_0_85_391 ();
 sg13g2_fill_2 FILLER_0_85_402 ();
 sg13g2_fill_2 FILLER_0_85_421 ();
 sg13g2_decap_8 FILLER_0_85_427 ();
 sg13g2_decap_8 FILLER_0_85_434 ();
 sg13g2_fill_2 FILLER_0_85_441 ();
 sg13g2_fill_1 FILLER_0_85_443 ();
 sg13g2_decap_4 FILLER_0_85_448 ();
 sg13g2_decap_8 FILLER_0_85_463 ();
 sg13g2_decap_4 FILLER_0_85_470 ();
 sg13g2_decap_4 FILLER_0_85_479 ();
 sg13g2_fill_2 FILLER_0_85_488 ();
 sg13g2_decap_8 FILLER_0_85_501 ();
 sg13g2_fill_2 FILLER_0_85_508 ();
 sg13g2_fill_2 FILLER_0_85_518 ();
 sg13g2_decap_8 FILLER_0_85_556 ();
 sg13g2_decap_8 FILLER_0_85_563 ();
 sg13g2_decap_4 FILLER_0_85_570 ();
 sg13g2_fill_2 FILLER_0_85_577 ();
 sg13g2_fill_2 FILLER_0_85_584 ();
 sg13g2_fill_1 FILLER_0_85_586 ();
 sg13g2_decap_8 FILLER_0_85_592 ();
 sg13g2_decap_8 FILLER_0_85_599 ();
 sg13g2_decap_8 FILLER_0_85_606 ();
 sg13g2_decap_8 FILLER_0_85_613 ();
 sg13g2_fill_1 FILLER_0_85_620 ();
 sg13g2_fill_1 FILLER_0_85_652 ();
 sg13g2_fill_1 FILLER_0_85_666 ();
 sg13g2_decap_4 FILLER_0_85_677 ();
 sg13g2_fill_2 FILLER_0_85_681 ();
 sg13g2_fill_2 FILLER_0_85_687 ();
 sg13g2_fill_1 FILLER_0_85_689 ();
 sg13g2_decap_8 FILLER_0_85_707 ();
 sg13g2_decap_8 FILLER_0_85_714 ();
 sg13g2_decap_8 FILLER_0_85_721 ();
 sg13g2_fill_2 FILLER_0_85_728 ();
 sg13g2_fill_1 FILLER_0_85_730 ();
 sg13g2_fill_1 FILLER_0_85_754 ();
 sg13g2_fill_1 FILLER_0_85_765 ();
 sg13g2_decap_8 FILLER_0_85_792 ();
 sg13g2_fill_2 FILLER_0_85_799 ();
 sg13g2_fill_1 FILLER_0_85_801 ();
 sg13g2_fill_2 FILLER_0_85_833 ();
 sg13g2_fill_1 FILLER_0_85_835 ();
 sg13g2_decap_8 FILLER_0_85_841 ();
 sg13g2_fill_1 FILLER_0_85_848 ();
 sg13g2_fill_2 FILLER_0_85_859 ();
 sg13g2_decap_8 FILLER_0_85_891 ();
 sg13g2_decap_8 FILLER_0_85_898 ();
 sg13g2_decap_8 FILLER_0_85_905 ();
 sg13g2_decap_8 FILLER_0_85_912 ();
 sg13g2_decap_8 FILLER_0_85_919 ();
 sg13g2_decap_8 FILLER_0_85_926 ();
 sg13g2_decap_8 FILLER_0_85_933 ();
 sg13g2_decap_8 FILLER_0_85_940 ();
 sg13g2_decap_8 FILLER_0_85_947 ();
 sg13g2_decap_8 FILLER_0_85_954 ();
 sg13g2_decap_8 FILLER_0_85_961 ();
 sg13g2_decap_8 FILLER_0_85_968 ();
 sg13g2_decap_8 FILLER_0_85_975 ();
 sg13g2_decap_8 FILLER_0_85_982 ();
 sg13g2_decap_8 FILLER_0_85_989 ();
 sg13g2_decap_8 FILLER_0_85_996 ();
 sg13g2_decap_8 FILLER_0_85_1003 ();
 sg13g2_decap_8 FILLER_0_85_1010 ();
 sg13g2_decap_8 FILLER_0_85_1017 ();
 sg13g2_decap_8 FILLER_0_85_1024 ();
 sg13g2_decap_8 FILLER_0_85_1031 ();
 sg13g2_decap_8 FILLER_0_85_1038 ();
 sg13g2_decap_8 FILLER_0_85_1045 ();
 sg13g2_decap_8 FILLER_0_85_1052 ();
 sg13g2_decap_8 FILLER_0_85_1059 ();
 sg13g2_decap_8 FILLER_0_85_1066 ();
 sg13g2_decap_8 FILLER_0_85_1073 ();
 sg13g2_decap_8 FILLER_0_85_1080 ();
 sg13g2_decap_8 FILLER_0_85_1087 ();
 sg13g2_decap_8 FILLER_0_85_1094 ();
 sg13g2_decap_8 FILLER_0_85_1101 ();
 sg13g2_decap_8 FILLER_0_85_1108 ();
 sg13g2_decap_8 FILLER_0_85_1115 ();
 sg13g2_decap_8 FILLER_0_85_1122 ();
 sg13g2_decap_8 FILLER_0_85_1129 ();
 sg13g2_decap_8 FILLER_0_85_1136 ();
 sg13g2_decap_8 FILLER_0_85_1143 ();
 sg13g2_decap_8 FILLER_0_85_1150 ();
 sg13g2_decap_8 FILLER_0_85_1157 ();
 sg13g2_decap_8 FILLER_0_85_1164 ();
 sg13g2_decap_8 FILLER_0_85_1171 ();
 sg13g2_decap_8 FILLER_0_85_1178 ();
 sg13g2_decap_8 FILLER_0_85_1185 ();
 sg13g2_decap_8 FILLER_0_85_1192 ();
 sg13g2_decap_8 FILLER_0_85_1199 ();
 sg13g2_decap_8 FILLER_0_85_1206 ();
 sg13g2_decap_8 FILLER_0_85_1213 ();
 sg13g2_decap_8 FILLER_0_85_1220 ();
 sg13g2_fill_1 FILLER_0_85_1227 ();
 sg13g2_decap_4 FILLER_0_86_0 ();
 sg13g2_decap_8 FILLER_0_86_40 ();
 sg13g2_decap_8 FILLER_0_86_47 ();
 sg13g2_fill_1 FILLER_0_86_54 ();
 sg13g2_decap_8 FILLER_0_86_63 ();
 sg13g2_decap_4 FILLER_0_86_88 ();
 sg13g2_decap_8 FILLER_0_86_152 ();
 sg13g2_decap_8 FILLER_0_86_159 ();
 sg13g2_fill_2 FILLER_0_86_166 ();
 sg13g2_fill_1 FILLER_0_86_168 ();
 sg13g2_fill_2 FILLER_0_86_174 ();
 sg13g2_fill_2 FILLER_0_86_186 ();
 sg13g2_fill_1 FILLER_0_86_188 ();
 sg13g2_decap_8 FILLER_0_86_228 ();
 sg13g2_fill_1 FILLER_0_86_239 ();
 sg13g2_fill_1 FILLER_0_86_286 ();
 sg13g2_decap_8 FILLER_0_86_301 ();
 sg13g2_decap_4 FILLER_0_86_308 ();
 sg13g2_fill_1 FILLER_0_86_316 ();
 sg13g2_fill_1 FILLER_0_86_321 ();
 sg13g2_fill_2 FILLER_0_86_327 ();
 sg13g2_fill_2 FILLER_0_86_339 ();
 sg13g2_fill_2 FILLER_0_86_367 ();
 sg13g2_fill_1 FILLER_0_86_369 ();
 sg13g2_decap_4 FILLER_0_86_396 ();
 sg13g2_fill_2 FILLER_0_86_400 ();
 sg13g2_decap_8 FILLER_0_86_407 ();
 sg13g2_decap_8 FILLER_0_86_414 ();
 sg13g2_decap_8 FILLER_0_86_421 ();
 sg13g2_decap_8 FILLER_0_86_428 ();
 sg13g2_decap_8 FILLER_0_86_435 ();
 sg13g2_decap_8 FILLER_0_86_442 ();
 sg13g2_decap_8 FILLER_0_86_449 ();
 sg13g2_decap_4 FILLER_0_86_456 ();
 sg13g2_fill_2 FILLER_0_86_465 ();
 sg13g2_fill_1 FILLER_0_86_467 ();
 sg13g2_fill_2 FILLER_0_86_525 ();
 sg13g2_decap_4 FILLER_0_86_553 ();
 sg13g2_fill_1 FILLER_0_86_557 ();
 sg13g2_decap_4 FILLER_0_86_563 ();
 sg13g2_fill_1 FILLER_0_86_571 ();
 sg13g2_fill_1 FILLER_0_86_582 ();
 sg13g2_fill_1 FILLER_0_86_609 ();
 sg13g2_fill_1 FILLER_0_86_641 ();
 sg13g2_fill_1 FILLER_0_86_646 ();
 sg13g2_decap_8 FILLER_0_86_681 ();
 sg13g2_decap_8 FILLER_0_86_688 ();
 sg13g2_decap_8 FILLER_0_86_695 ();
 sg13g2_decap_4 FILLER_0_86_702 ();
 sg13g2_fill_1 FILLER_0_86_706 ();
 sg13g2_decap_4 FILLER_0_86_711 ();
 sg13g2_fill_2 FILLER_0_86_715 ();
 sg13g2_decap_8 FILLER_0_86_722 ();
 sg13g2_decap_8 FILLER_0_86_729 ();
 sg13g2_decap_8 FILLER_0_86_736 ();
 sg13g2_fill_2 FILLER_0_86_743 ();
 sg13g2_fill_1 FILLER_0_86_745 ();
 sg13g2_fill_2 FILLER_0_86_750 ();
 sg13g2_fill_1 FILLER_0_86_752 ();
 sg13g2_fill_1 FILLER_0_86_801 ();
 sg13g2_fill_1 FILLER_0_86_812 ();
 sg13g2_fill_1 FILLER_0_86_817 ();
 sg13g2_fill_2 FILLER_0_86_828 ();
 sg13g2_fill_1 FILLER_0_86_860 ();
 sg13g2_decap_8 FILLER_0_86_897 ();
 sg13g2_decap_8 FILLER_0_86_904 ();
 sg13g2_decap_8 FILLER_0_86_911 ();
 sg13g2_decap_8 FILLER_0_86_918 ();
 sg13g2_decap_8 FILLER_0_86_925 ();
 sg13g2_decap_8 FILLER_0_86_932 ();
 sg13g2_decap_8 FILLER_0_86_939 ();
 sg13g2_decap_8 FILLER_0_86_946 ();
 sg13g2_decap_8 FILLER_0_86_953 ();
 sg13g2_decap_8 FILLER_0_86_960 ();
 sg13g2_decap_8 FILLER_0_86_967 ();
 sg13g2_decap_8 FILLER_0_86_974 ();
 sg13g2_decap_8 FILLER_0_86_981 ();
 sg13g2_decap_8 FILLER_0_86_988 ();
 sg13g2_decap_8 FILLER_0_86_995 ();
 sg13g2_decap_8 FILLER_0_86_1002 ();
 sg13g2_decap_8 FILLER_0_86_1009 ();
 sg13g2_decap_8 FILLER_0_86_1016 ();
 sg13g2_decap_8 FILLER_0_86_1023 ();
 sg13g2_decap_8 FILLER_0_86_1030 ();
 sg13g2_decap_8 FILLER_0_86_1037 ();
 sg13g2_decap_8 FILLER_0_86_1044 ();
 sg13g2_decap_8 FILLER_0_86_1051 ();
 sg13g2_decap_8 FILLER_0_86_1058 ();
 sg13g2_decap_8 FILLER_0_86_1065 ();
 sg13g2_decap_8 FILLER_0_86_1072 ();
 sg13g2_decap_8 FILLER_0_86_1079 ();
 sg13g2_decap_8 FILLER_0_86_1086 ();
 sg13g2_decap_8 FILLER_0_86_1093 ();
 sg13g2_decap_8 FILLER_0_86_1100 ();
 sg13g2_decap_8 FILLER_0_86_1107 ();
 sg13g2_decap_8 FILLER_0_86_1114 ();
 sg13g2_decap_8 FILLER_0_86_1121 ();
 sg13g2_decap_8 FILLER_0_86_1128 ();
 sg13g2_decap_8 FILLER_0_86_1135 ();
 sg13g2_decap_8 FILLER_0_86_1142 ();
 sg13g2_decap_8 FILLER_0_86_1149 ();
 sg13g2_decap_8 FILLER_0_86_1156 ();
 sg13g2_decap_8 FILLER_0_86_1163 ();
 sg13g2_decap_8 FILLER_0_86_1170 ();
 sg13g2_decap_8 FILLER_0_86_1177 ();
 sg13g2_decap_8 FILLER_0_86_1184 ();
 sg13g2_decap_8 FILLER_0_86_1191 ();
 sg13g2_decap_8 FILLER_0_86_1198 ();
 sg13g2_decap_8 FILLER_0_86_1205 ();
 sg13g2_decap_8 FILLER_0_86_1212 ();
 sg13g2_decap_8 FILLER_0_86_1219 ();
 sg13g2_fill_2 FILLER_0_86_1226 ();
 sg13g2_decap_8 FILLER_0_87_0 ();
 sg13g2_decap_4 FILLER_0_87_7 ();
 sg13g2_fill_2 FILLER_0_87_20 ();
 sg13g2_fill_1 FILLER_0_87_22 ();
 sg13g2_decap_8 FILLER_0_87_33 ();
 sg13g2_decap_8 FILLER_0_87_40 ();
 sg13g2_decap_8 FILLER_0_87_47 ();
 sg13g2_decap_8 FILLER_0_87_62 ();
 sg13g2_fill_1 FILLER_0_87_69 ();
 sg13g2_fill_1 FILLER_0_87_105 ();
 sg13g2_decap_4 FILLER_0_87_114 ();
 sg13g2_fill_1 FILLER_0_87_118 ();
 sg13g2_decap_8 FILLER_0_87_138 ();
 sg13g2_decap_4 FILLER_0_87_145 ();
 sg13g2_fill_1 FILLER_0_87_149 ();
 sg13g2_decap_4 FILLER_0_87_232 ();
 sg13g2_fill_2 FILLER_0_87_274 ();
 sg13g2_decap_8 FILLER_0_87_291 ();
 sg13g2_fill_2 FILLER_0_87_298 ();
 sg13g2_fill_1 FILLER_0_87_300 ();
 sg13g2_fill_1 FILLER_0_87_336 ();
 sg13g2_fill_1 FILLER_0_87_342 ();
 sg13g2_fill_2 FILLER_0_87_353 ();
 sg13g2_fill_2 FILLER_0_87_359 ();
 sg13g2_fill_1 FILLER_0_87_371 ();
 sg13g2_decap_8 FILLER_0_87_418 ();
 sg13g2_decap_8 FILLER_0_87_425 ();
 sg13g2_decap_8 FILLER_0_87_432 ();
 sg13g2_fill_1 FILLER_0_87_536 ();
 sg13g2_fill_1 FILLER_0_87_541 ();
 sg13g2_fill_2 FILLER_0_87_571 ();
 sg13g2_fill_2 FILLER_0_87_599 ();
 sg13g2_fill_1 FILLER_0_87_601 ();
 sg13g2_fill_2 FILLER_0_87_628 ();
 sg13g2_fill_1 FILLER_0_87_630 ();
 sg13g2_fill_1 FILLER_0_87_674 ();
 sg13g2_fill_1 FILLER_0_87_685 ();
 sg13g2_decap_4 FILLER_0_87_696 ();
 sg13g2_fill_2 FILLER_0_87_700 ();
 sg13g2_fill_1 FILLER_0_87_728 ();
 sg13g2_decap_8 FILLER_0_87_748 ();
 sg13g2_decap_8 FILLER_0_87_755 ();
 sg13g2_decap_8 FILLER_0_87_762 ();
 sg13g2_fill_1 FILLER_0_87_797 ();
 sg13g2_decap_8 FILLER_0_87_829 ();
 sg13g2_fill_2 FILLER_0_87_841 ();
 sg13g2_fill_2 FILLER_0_87_853 ();
 sg13g2_decap_8 FILLER_0_87_865 ();
 sg13g2_fill_2 FILLER_0_87_872 ();
 sg13g2_fill_1 FILLER_0_87_878 ();
 sg13g2_decap_8 FILLER_0_87_884 ();
 sg13g2_decap_8 FILLER_0_87_891 ();
 sg13g2_decap_8 FILLER_0_87_898 ();
 sg13g2_decap_8 FILLER_0_87_905 ();
 sg13g2_decap_8 FILLER_0_87_912 ();
 sg13g2_decap_8 FILLER_0_87_919 ();
 sg13g2_decap_8 FILLER_0_87_926 ();
 sg13g2_decap_8 FILLER_0_87_933 ();
 sg13g2_decap_8 FILLER_0_87_940 ();
 sg13g2_decap_8 FILLER_0_87_947 ();
 sg13g2_decap_8 FILLER_0_87_954 ();
 sg13g2_decap_8 FILLER_0_87_961 ();
 sg13g2_decap_8 FILLER_0_87_968 ();
 sg13g2_decap_8 FILLER_0_87_975 ();
 sg13g2_decap_8 FILLER_0_87_982 ();
 sg13g2_decap_8 FILLER_0_87_989 ();
 sg13g2_decap_8 FILLER_0_87_996 ();
 sg13g2_decap_8 FILLER_0_87_1003 ();
 sg13g2_decap_8 FILLER_0_87_1010 ();
 sg13g2_decap_8 FILLER_0_87_1017 ();
 sg13g2_decap_8 FILLER_0_87_1024 ();
 sg13g2_decap_8 FILLER_0_87_1031 ();
 sg13g2_decap_8 FILLER_0_87_1038 ();
 sg13g2_decap_8 FILLER_0_87_1045 ();
 sg13g2_decap_8 FILLER_0_87_1052 ();
 sg13g2_decap_8 FILLER_0_87_1059 ();
 sg13g2_decap_8 FILLER_0_87_1066 ();
 sg13g2_decap_8 FILLER_0_87_1073 ();
 sg13g2_decap_8 FILLER_0_87_1080 ();
 sg13g2_decap_8 FILLER_0_87_1087 ();
 sg13g2_decap_8 FILLER_0_87_1094 ();
 sg13g2_decap_8 FILLER_0_87_1101 ();
 sg13g2_decap_8 FILLER_0_87_1108 ();
 sg13g2_decap_8 FILLER_0_87_1115 ();
 sg13g2_decap_8 FILLER_0_87_1122 ();
 sg13g2_decap_8 FILLER_0_87_1129 ();
 sg13g2_decap_8 FILLER_0_87_1136 ();
 sg13g2_decap_8 FILLER_0_87_1143 ();
 sg13g2_decap_8 FILLER_0_87_1150 ();
 sg13g2_decap_8 FILLER_0_87_1157 ();
 sg13g2_decap_8 FILLER_0_87_1164 ();
 sg13g2_decap_8 FILLER_0_87_1171 ();
 sg13g2_decap_8 FILLER_0_87_1178 ();
 sg13g2_decap_8 FILLER_0_87_1185 ();
 sg13g2_decap_8 FILLER_0_87_1192 ();
 sg13g2_decap_8 FILLER_0_87_1199 ();
 sg13g2_decap_8 FILLER_0_87_1206 ();
 sg13g2_decap_8 FILLER_0_87_1213 ();
 sg13g2_decap_8 FILLER_0_87_1220 ();
 sg13g2_fill_1 FILLER_0_87_1227 ();
 sg13g2_decap_4 FILLER_0_88_0 ();
 sg13g2_fill_2 FILLER_0_88_4 ();
 sg13g2_fill_2 FILLER_0_88_37 ();
 sg13g2_fill_2 FILLER_0_88_65 ();
 sg13g2_decap_4 FILLER_0_88_74 ();
 sg13g2_fill_2 FILLER_0_88_78 ();
 sg13g2_fill_2 FILLER_0_88_103 ();
 sg13g2_fill_1 FILLER_0_88_105 ();
 sg13g2_decap_8 FILLER_0_88_147 ();
 sg13g2_decap_4 FILLER_0_88_154 ();
 sg13g2_fill_1 FILLER_0_88_158 ();
 sg13g2_fill_1 FILLER_0_88_217 ();
 sg13g2_decap_8 FILLER_0_88_222 ();
 sg13g2_decap_8 FILLER_0_88_229 ();
 sg13g2_decap_8 FILLER_0_88_236 ();
 sg13g2_decap_8 FILLER_0_88_243 ();
 sg13g2_decap_8 FILLER_0_88_254 ();
 sg13g2_decap_4 FILLER_0_88_261 ();
 sg13g2_fill_2 FILLER_0_88_304 ();
 sg13g2_fill_1 FILLER_0_88_311 ();
 sg13g2_fill_1 FILLER_0_88_317 ();
 sg13g2_fill_1 FILLER_0_88_323 ();
 sg13g2_fill_1 FILLER_0_88_339 ();
 sg13g2_decap_4 FILLER_0_88_355 ();
 sg13g2_fill_2 FILLER_0_88_359 ();
 sg13g2_fill_2 FILLER_0_88_378 ();
 sg13g2_fill_1 FILLER_0_88_380 ();
 sg13g2_fill_1 FILLER_0_88_386 ();
 sg13g2_fill_1 FILLER_0_88_397 ();
 sg13g2_fill_1 FILLER_0_88_403 ();
 sg13g2_fill_1 FILLER_0_88_435 ();
 sg13g2_fill_2 FILLER_0_88_495 ();
 sg13g2_fill_2 FILLER_0_88_507 ();
 sg13g2_fill_1 FILLER_0_88_509 ();
 sg13g2_decap_8 FILLER_0_88_524 ();
 sg13g2_decap_4 FILLER_0_88_531 ();
 sg13g2_fill_2 FILLER_0_88_535 ();
 sg13g2_fill_1 FILLER_0_88_586 ();
 sg13g2_fill_1 FILLER_0_88_591 ();
 sg13g2_fill_2 FILLER_0_88_637 ();
 sg13g2_fill_1 FILLER_0_88_674 ();
 sg13g2_decap_8 FILLER_0_88_680 ();
 sg13g2_decap_4 FILLER_0_88_687 ();
 sg13g2_decap_4 FILLER_0_88_762 ();
 sg13g2_fill_1 FILLER_0_88_766 ();
 sg13g2_fill_2 FILLER_0_88_793 ();
 sg13g2_fill_1 FILLER_0_88_795 ();
 sg13g2_decap_8 FILLER_0_88_804 ();
 sg13g2_fill_1 FILLER_0_88_815 ();
 sg13g2_fill_2 FILLER_0_88_829 ();
 sg13g2_fill_1 FILLER_0_88_831 ();
 sg13g2_decap_4 FILLER_0_88_875 ();
 sg13g2_decap_8 FILLER_0_88_883 ();
 sg13g2_decap_8 FILLER_0_88_890 ();
 sg13g2_decap_8 FILLER_0_88_897 ();
 sg13g2_decap_8 FILLER_0_88_904 ();
 sg13g2_decap_8 FILLER_0_88_911 ();
 sg13g2_fill_2 FILLER_0_88_918 ();
 sg13g2_fill_1 FILLER_0_88_920 ();
 sg13g2_fill_1 FILLER_0_88_925 ();
 sg13g2_fill_1 FILLER_0_88_931 ();
 sg13g2_fill_1 FILLER_0_88_942 ();
 sg13g2_fill_2 FILLER_0_88_947 ();
 sg13g2_decap_8 FILLER_0_88_954 ();
 sg13g2_decap_8 FILLER_0_88_961 ();
 sg13g2_decap_8 FILLER_0_88_968 ();
 sg13g2_decap_8 FILLER_0_88_975 ();
 sg13g2_decap_8 FILLER_0_88_982 ();
 sg13g2_decap_8 FILLER_0_88_989 ();
 sg13g2_decap_8 FILLER_0_88_996 ();
 sg13g2_decap_8 FILLER_0_88_1003 ();
 sg13g2_decap_8 FILLER_0_88_1010 ();
 sg13g2_decap_8 FILLER_0_88_1017 ();
 sg13g2_decap_8 FILLER_0_88_1024 ();
 sg13g2_decap_8 FILLER_0_88_1031 ();
 sg13g2_decap_8 FILLER_0_88_1038 ();
 sg13g2_decap_8 FILLER_0_88_1045 ();
 sg13g2_decap_8 FILLER_0_88_1052 ();
 sg13g2_decap_8 FILLER_0_88_1059 ();
 sg13g2_decap_8 FILLER_0_88_1066 ();
 sg13g2_decap_8 FILLER_0_88_1073 ();
 sg13g2_decap_8 FILLER_0_88_1080 ();
 sg13g2_decap_8 FILLER_0_88_1087 ();
 sg13g2_decap_8 FILLER_0_88_1094 ();
 sg13g2_decap_8 FILLER_0_88_1101 ();
 sg13g2_decap_8 FILLER_0_88_1108 ();
 sg13g2_decap_8 FILLER_0_88_1115 ();
 sg13g2_decap_8 FILLER_0_88_1122 ();
 sg13g2_decap_8 FILLER_0_88_1129 ();
 sg13g2_decap_8 FILLER_0_88_1136 ();
 sg13g2_decap_8 FILLER_0_88_1143 ();
 sg13g2_decap_8 FILLER_0_88_1150 ();
 sg13g2_decap_8 FILLER_0_88_1157 ();
 sg13g2_decap_8 FILLER_0_88_1164 ();
 sg13g2_decap_8 FILLER_0_88_1171 ();
 sg13g2_decap_8 FILLER_0_88_1178 ();
 sg13g2_decap_8 FILLER_0_88_1185 ();
 sg13g2_decap_8 FILLER_0_88_1192 ();
 sg13g2_decap_8 FILLER_0_88_1199 ();
 sg13g2_decap_8 FILLER_0_88_1206 ();
 sg13g2_decap_8 FILLER_0_88_1213 ();
 sg13g2_decap_8 FILLER_0_88_1220 ();
 sg13g2_fill_1 FILLER_0_88_1227 ();
 sg13g2_fill_1 FILLER_0_89_0 ();
 sg13g2_fill_1 FILLER_0_89_5 ();
 sg13g2_fill_1 FILLER_0_89_32 ();
 sg13g2_fill_1 FILLER_0_89_38 ();
 sg13g2_fill_1 FILLER_0_89_43 ();
 sg13g2_fill_2 FILLER_0_89_74 ();
 sg13g2_fill_2 FILLER_0_89_102 ();
 sg13g2_fill_1 FILLER_0_89_104 ();
 sg13g2_fill_2 FILLER_0_89_110 ();
 sg13g2_fill_1 FILLER_0_89_112 ();
 sg13g2_fill_2 FILLER_0_89_117 ();
 sg13g2_decap_4 FILLER_0_89_123 ();
 sg13g2_fill_2 FILLER_0_89_137 ();
 sg13g2_fill_1 FILLER_0_89_139 ();
 sg13g2_fill_2 FILLER_0_89_170 ();
 sg13g2_fill_2 FILLER_0_89_182 ();
 sg13g2_fill_1 FILLER_0_89_184 ();
 sg13g2_decap_4 FILLER_0_89_195 ();
 sg13g2_fill_1 FILLER_0_89_199 ();
 sg13g2_decap_8 FILLER_0_89_208 ();
 sg13g2_decap_4 FILLER_0_89_215 ();
 sg13g2_decap_8 FILLER_0_89_224 ();
 sg13g2_decap_8 FILLER_0_89_231 ();
 sg13g2_decap_4 FILLER_0_89_238 ();
 sg13g2_fill_1 FILLER_0_89_242 ();
 sg13g2_fill_1 FILLER_0_89_269 ();
 sg13g2_fill_1 FILLER_0_89_335 ();
 sg13g2_fill_2 FILLER_0_89_341 ();
 sg13g2_fill_2 FILLER_0_89_369 ();
 sg13g2_fill_1 FILLER_0_89_371 ();
 sg13g2_decap_4 FILLER_0_89_376 ();
 sg13g2_fill_2 FILLER_0_89_380 ();
 sg13g2_fill_2 FILLER_0_89_386 ();
 sg13g2_fill_1 FILLER_0_89_388 ();
 sg13g2_fill_2 FILLER_0_89_393 ();
 sg13g2_fill_1 FILLER_0_89_421 ();
 sg13g2_fill_1 FILLER_0_89_452 ();
 sg13g2_decap_4 FILLER_0_89_467 ();
 sg13g2_decap_8 FILLER_0_89_476 ();
 sg13g2_decap_8 FILLER_0_89_483 ();
 sg13g2_decap_4 FILLER_0_89_490 ();
 sg13g2_fill_1 FILLER_0_89_494 ();
 sg13g2_fill_1 FILLER_0_89_505 ();
 sg13g2_decap_8 FILLER_0_89_510 ();
 sg13g2_decap_4 FILLER_0_89_517 ();
 sg13g2_decap_4 FILLER_0_89_526 ();
 sg13g2_fill_2 FILLER_0_89_530 ();
 sg13g2_fill_1 FILLER_0_89_578 ();
 sg13g2_decap_8 FILLER_0_89_591 ();
 sg13g2_fill_2 FILLER_0_89_606 ();
 sg13g2_decap_4 FILLER_0_89_621 ();
 sg13g2_fill_2 FILLER_0_89_638 ();
 sg13g2_fill_1 FILLER_0_89_644 ();
 sg13g2_decap_8 FILLER_0_89_650 ();
 sg13g2_fill_1 FILLER_0_89_657 ();
 sg13g2_fill_1 FILLER_0_89_692 ();
 sg13g2_fill_2 FILLER_0_89_770 ();
 sg13g2_fill_1 FILLER_0_89_776 ();
 sg13g2_fill_2 FILLER_0_89_782 ();
 sg13g2_decap_4 FILLER_0_89_794 ();
 sg13g2_fill_2 FILLER_0_89_798 ();
 sg13g2_decap_8 FILLER_0_89_831 ();
 sg13g2_decap_8 FILLER_0_89_838 ();
 sg13g2_fill_1 FILLER_0_89_888 ();
 sg13g2_fill_1 FILLER_0_89_897 ();
 sg13g2_decap_8 FILLER_0_89_903 ();
 sg13g2_decap_4 FILLER_0_89_910 ();
 sg13g2_fill_1 FILLER_0_89_914 ();
 sg13g2_decap_8 FILLER_0_89_982 ();
 sg13g2_decap_8 FILLER_0_89_989 ();
 sg13g2_decap_8 FILLER_0_89_996 ();
 sg13g2_decap_8 FILLER_0_89_1003 ();
 sg13g2_decap_8 FILLER_0_89_1010 ();
 sg13g2_decap_8 FILLER_0_89_1017 ();
 sg13g2_decap_8 FILLER_0_89_1024 ();
 sg13g2_decap_8 FILLER_0_89_1031 ();
 sg13g2_decap_8 FILLER_0_89_1038 ();
 sg13g2_decap_8 FILLER_0_89_1045 ();
 sg13g2_decap_8 FILLER_0_89_1052 ();
 sg13g2_decap_8 FILLER_0_89_1059 ();
 sg13g2_decap_8 FILLER_0_89_1066 ();
 sg13g2_decap_8 FILLER_0_89_1073 ();
 sg13g2_decap_8 FILLER_0_89_1080 ();
 sg13g2_decap_8 FILLER_0_89_1087 ();
 sg13g2_decap_8 FILLER_0_89_1094 ();
 sg13g2_decap_8 FILLER_0_89_1101 ();
 sg13g2_decap_8 FILLER_0_89_1108 ();
 sg13g2_decap_8 FILLER_0_89_1115 ();
 sg13g2_decap_8 FILLER_0_89_1122 ();
 sg13g2_decap_8 FILLER_0_89_1129 ();
 sg13g2_decap_8 FILLER_0_89_1136 ();
 sg13g2_decap_8 FILLER_0_89_1143 ();
 sg13g2_decap_8 FILLER_0_89_1150 ();
 sg13g2_decap_8 FILLER_0_89_1157 ();
 sg13g2_decap_8 FILLER_0_89_1164 ();
 sg13g2_decap_8 FILLER_0_89_1171 ();
 sg13g2_decap_8 FILLER_0_89_1178 ();
 sg13g2_decap_8 FILLER_0_89_1185 ();
 sg13g2_decap_8 FILLER_0_89_1192 ();
 sg13g2_decap_8 FILLER_0_89_1199 ();
 sg13g2_decap_8 FILLER_0_89_1206 ();
 sg13g2_decap_8 FILLER_0_89_1213 ();
 sg13g2_decap_8 FILLER_0_89_1220 ();
 sg13g2_fill_1 FILLER_0_89_1227 ();
 sg13g2_fill_2 FILLER_0_90_0 ();
 sg13g2_fill_2 FILLER_0_90_6 ();
 sg13g2_fill_2 FILLER_0_90_13 ();
 sg13g2_fill_1 FILLER_0_90_15 ();
 sg13g2_fill_1 FILLER_0_90_26 ();
 sg13g2_fill_1 FILLER_0_90_47 ();
 sg13g2_fill_1 FILLER_0_90_52 ();
 sg13g2_fill_2 FILLER_0_90_65 ();
 sg13g2_fill_1 FILLER_0_90_86 ();
 sg13g2_fill_1 FILLER_0_90_97 ();
 sg13g2_fill_1 FILLER_0_90_106 ();
 sg13g2_decap_8 FILLER_0_90_143 ();
 sg13g2_fill_2 FILLER_0_90_150 ();
 sg13g2_decap_8 FILLER_0_90_156 ();
 sg13g2_decap_4 FILLER_0_90_163 ();
 sg13g2_fill_2 FILLER_0_90_193 ();
 sg13g2_fill_1 FILLER_0_90_195 ();
 sg13g2_fill_2 FILLER_0_90_201 ();
 sg13g2_decap_8 FILLER_0_90_207 ();
 sg13g2_decap_8 FILLER_0_90_214 ();
 sg13g2_decap_8 FILLER_0_90_221 ();
 sg13g2_fill_1 FILLER_0_90_299 ();
 sg13g2_fill_1 FILLER_0_90_326 ();
 sg13g2_fill_2 FILLER_0_90_337 ();
 sg13g2_fill_2 FILLER_0_90_343 ();
 sg13g2_decap_8 FILLER_0_90_354 ();
 sg13g2_decap_8 FILLER_0_90_371 ();
 sg13g2_decap_8 FILLER_0_90_378 ();
 sg13g2_decap_8 FILLER_0_90_385 ();
 sg13g2_decap_8 FILLER_0_90_392 ();
 sg13g2_decap_4 FILLER_0_90_399 ();
 sg13g2_fill_2 FILLER_0_90_436 ();
 sg13g2_fill_1 FILLER_0_90_438 ();
 sg13g2_fill_2 FILLER_0_90_443 ();
 sg13g2_fill_1 FILLER_0_90_445 ();
 sg13g2_decap_8 FILLER_0_90_454 ();
 sg13g2_decap_8 FILLER_0_90_461 ();
 sg13g2_decap_8 FILLER_0_90_468 ();
 sg13g2_decap_8 FILLER_0_90_475 ();
 sg13g2_fill_2 FILLER_0_90_482 ();
 sg13g2_fill_1 FILLER_0_90_510 ();
 sg13g2_fill_2 FILLER_0_90_537 ();
 sg13g2_fill_1 FILLER_0_90_544 ();
 sg13g2_fill_2 FILLER_0_90_555 ();
 sg13g2_fill_1 FILLER_0_90_561 ();
 sg13g2_decap_8 FILLER_0_90_573 ();
 sg13g2_decap_8 FILLER_0_90_580 ();
 sg13g2_decap_8 FILLER_0_90_587 ();
 sg13g2_decap_8 FILLER_0_90_594 ();
 sg13g2_decap_8 FILLER_0_90_601 ();
 sg13g2_decap_8 FILLER_0_90_608 ();
 sg13g2_decap_8 FILLER_0_90_615 ();
 sg13g2_fill_2 FILLER_0_90_634 ();
 sg13g2_decap_4 FILLER_0_90_667 ();
 sg13g2_decap_8 FILLER_0_90_675 ();
 sg13g2_decap_8 FILLER_0_90_682 ();
 sg13g2_decap_4 FILLER_0_90_694 ();
 sg13g2_fill_2 FILLER_0_90_698 ();
 sg13g2_decap_4 FILLER_0_90_709 ();
 sg13g2_fill_1 FILLER_0_90_713 ();
 sg13g2_fill_2 FILLER_0_90_718 ();
 sg13g2_decap_4 FILLER_0_90_742 ();
 sg13g2_fill_1 FILLER_0_90_750 ();
 sg13g2_decap_8 FILLER_0_90_790 ();
 sg13g2_fill_2 FILLER_0_90_797 ();
 sg13g2_fill_1 FILLER_0_90_811 ();
 sg13g2_fill_1 FILLER_0_90_817 ();
 sg13g2_fill_1 FILLER_0_90_828 ();
 sg13g2_fill_1 FILLER_0_90_834 ();
 sg13g2_fill_1 FILLER_0_90_845 ();
 sg13g2_fill_1 FILLER_0_90_856 ();
 sg13g2_fill_1 FILLER_0_90_892 ();
 sg13g2_fill_2 FILLER_0_90_943 ();
 sg13g2_decap_8 FILLER_0_90_955 ();
 sg13g2_decap_8 FILLER_0_90_966 ();
 sg13g2_decap_8 FILLER_0_90_973 ();
 sg13g2_decap_8 FILLER_0_90_980 ();
 sg13g2_decap_8 FILLER_0_90_987 ();
 sg13g2_decap_8 FILLER_0_90_994 ();
 sg13g2_decap_8 FILLER_0_90_1001 ();
 sg13g2_decap_8 FILLER_0_90_1008 ();
 sg13g2_decap_8 FILLER_0_90_1015 ();
 sg13g2_decap_8 FILLER_0_90_1022 ();
 sg13g2_decap_8 FILLER_0_90_1029 ();
 sg13g2_decap_8 FILLER_0_90_1036 ();
 sg13g2_decap_8 FILLER_0_90_1043 ();
 sg13g2_decap_8 FILLER_0_90_1050 ();
 sg13g2_decap_8 FILLER_0_90_1057 ();
 sg13g2_decap_8 FILLER_0_90_1064 ();
 sg13g2_decap_8 FILLER_0_90_1071 ();
 sg13g2_decap_8 FILLER_0_90_1078 ();
 sg13g2_decap_8 FILLER_0_90_1085 ();
 sg13g2_decap_8 FILLER_0_90_1092 ();
 sg13g2_decap_8 FILLER_0_90_1099 ();
 sg13g2_decap_8 FILLER_0_90_1106 ();
 sg13g2_decap_8 FILLER_0_90_1113 ();
 sg13g2_decap_8 FILLER_0_90_1120 ();
 sg13g2_decap_8 FILLER_0_90_1127 ();
 sg13g2_decap_8 FILLER_0_90_1134 ();
 sg13g2_decap_8 FILLER_0_90_1141 ();
 sg13g2_decap_8 FILLER_0_90_1148 ();
 sg13g2_decap_8 FILLER_0_90_1155 ();
 sg13g2_decap_8 FILLER_0_90_1162 ();
 sg13g2_decap_8 FILLER_0_90_1169 ();
 sg13g2_decap_8 FILLER_0_90_1176 ();
 sg13g2_decap_8 FILLER_0_90_1183 ();
 sg13g2_decap_8 FILLER_0_90_1190 ();
 sg13g2_decap_8 FILLER_0_90_1197 ();
 sg13g2_decap_8 FILLER_0_90_1204 ();
 sg13g2_decap_8 FILLER_0_90_1211 ();
 sg13g2_decap_8 FILLER_0_90_1218 ();
 sg13g2_fill_2 FILLER_0_90_1225 ();
 sg13g2_fill_1 FILLER_0_90_1227 ();
 sg13g2_decap_8 FILLER_0_91_0 ();
 sg13g2_decap_8 FILLER_0_91_7 ();
 sg13g2_decap_8 FILLER_0_91_14 ();
 sg13g2_fill_1 FILLER_0_91_25 ();
 sg13g2_fill_2 FILLER_0_91_49 ();
 sg13g2_fill_1 FILLER_0_91_55 ();
 sg13g2_fill_1 FILLER_0_91_66 ();
 sg13g2_fill_1 FILLER_0_91_71 ();
 sg13g2_fill_2 FILLER_0_91_107 ();
 sg13g2_fill_1 FILLER_0_91_109 ();
 sg13g2_fill_2 FILLER_0_91_136 ();
 sg13g2_fill_2 FILLER_0_91_143 ();
 sg13g2_fill_2 FILLER_0_91_171 ();
 sg13g2_fill_1 FILLER_0_91_173 ();
 sg13g2_decap_4 FILLER_0_91_178 ();
 sg13g2_fill_2 FILLER_0_91_182 ();
 sg13g2_fill_2 FILLER_0_91_210 ();
 sg13g2_fill_1 FILLER_0_91_212 ();
 sg13g2_decap_8 FILLER_0_91_227 ();
 sg13g2_decap_4 FILLER_0_91_234 ();
 sg13g2_fill_2 FILLER_0_91_242 ();
 sg13g2_fill_1 FILLER_0_91_249 ();
 sg13g2_fill_2 FILLER_0_91_260 ();
 sg13g2_fill_1 FILLER_0_91_272 ();
 sg13g2_fill_2 FILLER_0_91_278 ();
 sg13g2_fill_2 FILLER_0_91_284 ();
 sg13g2_decap_8 FILLER_0_91_290 ();
 sg13g2_fill_2 FILLER_0_91_297 ();
 sg13g2_fill_1 FILLER_0_91_299 ();
 sg13g2_decap_4 FILLER_0_91_309 ();
 sg13g2_fill_2 FILLER_0_91_313 ();
 sg13g2_fill_1 FILLER_0_91_338 ();
 sg13g2_decap_8 FILLER_0_91_369 ();
 sg13g2_fill_1 FILLER_0_91_376 ();
 sg13g2_decap_8 FILLER_0_91_385 ();
 sg13g2_decap_8 FILLER_0_91_392 ();
 sg13g2_decap_8 FILLER_0_91_399 ();
 sg13g2_decap_8 FILLER_0_91_406 ();
 sg13g2_decap_8 FILLER_0_91_413 ();
 sg13g2_decap_4 FILLER_0_91_420 ();
 sg13g2_fill_2 FILLER_0_91_424 ();
 sg13g2_decap_8 FILLER_0_91_431 ();
 sg13g2_decap_8 FILLER_0_91_438 ();
 sg13g2_decap_8 FILLER_0_91_445 ();
 sg13g2_decap_4 FILLER_0_91_452 ();
 sg13g2_decap_8 FILLER_0_91_461 ();
 sg13g2_fill_1 FILLER_0_91_468 ();
 sg13g2_fill_2 FILLER_0_91_473 ();
 sg13g2_fill_1 FILLER_0_91_475 ();
 sg13g2_fill_2 FILLER_0_91_483 ();
 sg13g2_decap_4 FILLER_0_91_495 ();
 sg13g2_fill_1 FILLER_0_91_499 ();
 sg13g2_fill_2 FILLER_0_91_513 ();
 sg13g2_fill_2 FILLER_0_91_525 ();
 sg13g2_decap_8 FILLER_0_91_553 ();
 sg13g2_fill_2 FILLER_0_91_560 ();
 sg13g2_fill_2 FILLER_0_91_565 ();
 sg13g2_fill_1 FILLER_0_91_567 ();
 sg13g2_decap_8 FILLER_0_91_599 ();
 sg13g2_decap_8 FILLER_0_91_606 ();
 sg13g2_fill_1 FILLER_0_91_613 ();
 sg13g2_fill_1 FILLER_0_91_622 ();
 sg13g2_fill_1 FILLER_0_91_649 ();
 sg13g2_fill_1 FILLER_0_91_676 ();
 sg13g2_fill_1 FILLER_0_91_695 ();
 sg13g2_fill_2 FILLER_0_91_706 ();
 sg13g2_decap_8 FILLER_0_91_712 ();
 sg13g2_fill_2 FILLER_0_91_719 ();
 sg13g2_decap_4 FILLER_0_91_755 ();
 sg13g2_fill_2 FILLER_0_91_759 ();
 sg13g2_decap_4 FILLER_0_91_766 ();
 sg13g2_fill_1 FILLER_0_91_770 ();
 sg13g2_fill_2 FILLER_0_91_900 ();
 sg13g2_fill_1 FILLER_0_91_938 ();
 sg13g2_decap_8 FILLER_0_91_975 ();
 sg13g2_decap_8 FILLER_0_91_982 ();
 sg13g2_decap_8 FILLER_0_91_989 ();
 sg13g2_decap_8 FILLER_0_91_996 ();
 sg13g2_decap_8 FILLER_0_91_1003 ();
 sg13g2_decap_8 FILLER_0_91_1010 ();
 sg13g2_decap_8 FILLER_0_91_1017 ();
 sg13g2_decap_8 FILLER_0_91_1024 ();
 sg13g2_decap_8 FILLER_0_91_1031 ();
 sg13g2_decap_8 FILLER_0_91_1038 ();
 sg13g2_decap_8 FILLER_0_91_1045 ();
 sg13g2_decap_8 FILLER_0_91_1052 ();
 sg13g2_decap_8 FILLER_0_91_1059 ();
 sg13g2_decap_8 FILLER_0_91_1066 ();
 sg13g2_decap_8 FILLER_0_91_1073 ();
 sg13g2_decap_8 FILLER_0_91_1080 ();
 sg13g2_decap_8 FILLER_0_91_1087 ();
 sg13g2_decap_8 FILLER_0_91_1094 ();
 sg13g2_decap_8 FILLER_0_91_1101 ();
 sg13g2_decap_8 FILLER_0_91_1108 ();
 sg13g2_decap_8 FILLER_0_91_1115 ();
 sg13g2_decap_8 FILLER_0_91_1122 ();
 sg13g2_decap_8 FILLER_0_91_1129 ();
 sg13g2_decap_8 FILLER_0_91_1136 ();
 sg13g2_decap_8 FILLER_0_91_1143 ();
 sg13g2_decap_8 FILLER_0_91_1150 ();
 sg13g2_decap_8 FILLER_0_91_1157 ();
 sg13g2_decap_8 FILLER_0_91_1164 ();
 sg13g2_decap_8 FILLER_0_91_1171 ();
 sg13g2_decap_8 FILLER_0_91_1178 ();
 sg13g2_decap_8 FILLER_0_91_1185 ();
 sg13g2_decap_8 FILLER_0_91_1192 ();
 sg13g2_decap_8 FILLER_0_91_1199 ();
 sg13g2_decap_8 FILLER_0_91_1206 ();
 sg13g2_decap_8 FILLER_0_91_1213 ();
 sg13g2_decap_8 FILLER_0_91_1220 ();
 sg13g2_fill_1 FILLER_0_91_1227 ();
 sg13g2_decap_4 FILLER_0_92_0 ();
 sg13g2_fill_2 FILLER_0_92_4 ();
 sg13g2_decap_4 FILLER_0_92_15 ();
 sg13g2_fill_1 FILLER_0_92_32 ();
 sg13g2_fill_1 FILLER_0_92_37 ();
 sg13g2_fill_2 FILLER_0_92_68 ();
 sg13g2_fill_2 FILLER_0_92_109 ();
 sg13g2_fill_1 FILLER_0_92_111 ();
 sg13g2_decap_4 FILLER_0_92_152 ();
 sg13g2_decap_4 FILLER_0_92_166 ();
 sg13g2_fill_2 FILLER_0_92_170 ();
 sg13g2_fill_2 FILLER_0_92_180 ();
 sg13g2_decap_4 FILLER_0_92_232 ();
 sg13g2_decap_8 FILLER_0_92_267 ();
 sg13g2_decap_8 FILLER_0_92_274 ();
 sg13g2_decap_8 FILLER_0_92_281 ();
 sg13g2_decap_8 FILLER_0_92_288 ();
 sg13g2_decap_4 FILLER_0_92_295 ();
 sg13g2_fill_2 FILLER_0_92_299 ();
 sg13g2_fill_1 FILLER_0_92_312 ();
 sg13g2_fill_2 FILLER_0_92_343 ();
 sg13g2_fill_1 FILLER_0_92_371 ();
 sg13g2_decap_4 FILLER_0_92_385 ();
 sg13g2_fill_2 FILLER_0_92_393 ();
 sg13g2_fill_1 FILLER_0_92_395 ();
 sg13g2_decap_8 FILLER_0_92_401 ();
 sg13g2_fill_1 FILLER_0_92_424 ();
 sg13g2_fill_1 FILLER_0_92_455 ();
 sg13g2_decap_4 FILLER_0_92_466 ();
 sg13g2_decap_8 FILLER_0_92_545 ();
 sg13g2_decap_8 FILLER_0_92_552 ();
 sg13g2_fill_2 FILLER_0_92_650 ();
 sg13g2_fill_1 FILLER_0_92_662 ();
 sg13g2_fill_1 FILLER_0_92_689 ();
 sg13g2_fill_2 FILLER_0_92_716 ();
 sg13g2_fill_2 FILLER_0_92_728 ();
 sg13g2_fill_1 FILLER_0_92_730 ();
 sg13g2_fill_2 FILLER_0_92_749 ();
 sg13g2_fill_2 FILLER_0_92_771 ();
 sg13g2_decap_4 FILLER_0_92_821 ();
 sg13g2_fill_1 FILLER_0_92_825 ();
 sg13g2_decap_4 FILLER_0_92_861 ();
 sg13g2_fill_2 FILLER_0_92_865 ();
 sg13g2_fill_1 FILLER_0_92_876 ();
 sg13g2_fill_1 FILLER_0_92_885 ();
 sg13g2_fill_1 FILLER_0_92_922 ();
 sg13g2_fill_2 FILLER_0_92_954 ();
 sg13g2_decap_8 FILLER_0_92_960 ();
 sg13g2_decap_8 FILLER_0_92_967 ();
 sg13g2_decap_8 FILLER_0_92_974 ();
 sg13g2_decap_8 FILLER_0_92_981 ();
 sg13g2_decap_8 FILLER_0_92_988 ();
 sg13g2_decap_8 FILLER_0_92_995 ();
 sg13g2_decap_8 FILLER_0_92_1002 ();
 sg13g2_decap_8 FILLER_0_92_1009 ();
 sg13g2_decap_8 FILLER_0_92_1016 ();
 sg13g2_decap_8 FILLER_0_92_1023 ();
 sg13g2_decap_8 FILLER_0_92_1030 ();
 sg13g2_decap_8 FILLER_0_92_1037 ();
 sg13g2_decap_8 FILLER_0_92_1044 ();
 sg13g2_decap_8 FILLER_0_92_1051 ();
 sg13g2_decap_8 FILLER_0_92_1058 ();
 sg13g2_decap_8 FILLER_0_92_1065 ();
 sg13g2_decap_8 FILLER_0_92_1072 ();
 sg13g2_decap_8 FILLER_0_92_1079 ();
 sg13g2_decap_8 FILLER_0_92_1086 ();
 sg13g2_decap_8 FILLER_0_92_1093 ();
 sg13g2_decap_8 FILLER_0_92_1100 ();
 sg13g2_decap_8 FILLER_0_92_1107 ();
 sg13g2_decap_8 FILLER_0_92_1114 ();
 sg13g2_decap_8 FILLER_0_92_1121 ();
 sg13g2_decap_8 FILLER_0_92_1128 ();
 sg13g2_decap_8 FILLER_0_92_1135 ();
 sg13g2_decap_8 FILLER_0_92_1142 ();
 sg13g2_decap_8 FILLER_0_92_1149 ();
 sg13g2_decap_8 FILLER_0_92_1156 ();
 sg13g2_decap_8 FILLER_0_92_1163 ();
 sg13g2_decap_8 FILLER_0_92_1170 ();
 sg13g2_decap_8 FILLER_0_92_1177 ();
 sg13g2_decap_8 FILLER_0_92_1184 ();
 sg13g2_decap_8 FILLER_0_92_1191 ();
 sg13g2_decap_8 FILLER_0_92_1198 ();
 sg13g2_decap_8 FILLER_0_92_1205 ();
 sg13g2_decap_8 FILLER_0_92_1212 ();
 sg13g2_decap_8 FILLER_0_92_1219 ();
 sg13g2_fill_2 FILLER_0_92_1226 ();
 sg13g2_decap_8 FILLER_0_93_0 ();
 sg13g2_fill_1 FILLER_0_93_7 ();
 sg13g2_fill_1 FILLER_0_93_42 ();
 sg13g2_decap_8 FILLER_0_93_53 ();
 sg13g2_decap_8 FILLER_0_93_60 ();
 sg13g2_fill_2 FILLER_0_93_67 ();
 sg13g2_decap_8 FILLER_0_93_99 ();
 sg13g2_decap_8 FILLER_0_93_106 ();
 sg13g2_decap_4 FILLER_0_93_113 ();
 sg13g2_decap_8 FILLER_0_93_121 ();
 sg13g2_decap_4 FILLER_0_93_128 ();
 sg13g2_fill_1 FILLER_0_93_132 ();
 sg13g2_fill_1 FILLER_0_93_142 ();
 sg13g2_fill_1 FILLER_0_93_148 ();
 sg13g2_fill_1 FILLER_0_93_154 ();
 sg13g2_fill_2 FILLER_0_93_186 ();
 sg13g2_decap_8 FILLER_0_93_272 ();
 sg13g2_decap_8 FILLER_0_93_279 ();
 sg13g2_decap_4 FILLER_0_93_286 ();
 sg13g2_fill_2 FILLER_0_93_290 ();
 sg13g2_fill_1 FILLER_0_93_297 ();
 sg13g2_fill_2 FILLER_0_93_308 ();
 sg13g2_decap_4 FILLER_0_93_340 ();
 sg13g2_fill_1 FILLER_0_93_344 ();
 sg13g2_decap_8 FILLER_0_93_380 ();
 sg13g2_decap_8 FILLER_0_93_387 ();
 sg13g2_decap_8 FILLER_0_93_394 ();
 sg13g2_fill_1 FILLER_0_93_401 ();
 sg13g2_decap_4 FILLER_0_93_496 ();
 sg13g2_fill_1 FILLER_0_93_500 ();
 sg13g2_fill_1 FILLER_0_93_520 ();
 sg13g2_decap_8 FILLER_0_93_525 ();
 sg13g2_decap_8 FILLER_0_93_532 ();
 sg13g2_fill_2 FILLER_0_93_539 ();
 sg13g2_fill_2 FILLER_0_93_572 ();
 sg13g2_fill_1 FILLER_0_93_574 ();
 sg13g2_fill_1 FILLER_0_93_579 ();
 sg13g2_fill_1 FILLER_0_93_590 ();
 sg13g2_fill_1 FILLER_0_93_601 ();
 sg13g2_fill_2 FILLER_0_93_645 ();
 sg13g2_fill_1 FILLER_0_93_651 ();
 sg13g2_fill_1 FILLER_0_93_657 ();
 sg13g2_fill_2 FILLER_0_93_662 ();
 sg13g2_fill_2 FILLER_0_93_674 ();
 sg13g2_fill_2 FILLER_0_93_680 ();
 sg13g2_fill_1 FILLER_0_93_682 ();
 sg13g2_decap_4 FILLER_0_93_688 ();
 sg13g2_fill_2 FILLER_0_93_692 ();
 sg13g2_fill_2 FILLER_0_93_698 ();
 sg13g2_fill_1 FILLER_0_93_700 ();
 sg13g2_fill_1 FILLER_0_93_727 ();
 sg13g2_fill_2 FILLER_0_93_773 ();
 sg13g2_fill_1 FILLER_0_93_775 ();
 sg13g2_decap_8 FILLER_0_93_815 ();
 sg13g2_decap_8 FILLER_0_93_822 ();
 sg13g2_decap_8 FILLER_0_93_829 ();
 sg13g2_decap_4 FILLER_0_93_836 ();
 sg13g2_decap_8 FILLER_0_93_848 ();
 sg13g2_decap_4 FILLER_0_93_855 ();
 sg13g2_fill_1 FILLER_0_93_859 ();
 sg13g2_fill_1 FILLER_0_93_878 ();
 sg13g2_decap_8 FILLER_0_93_884 ();
 sg13g2_decap_8 FILLER_0_93_891 ();
 sg13g2_decap_4 FILLER_0_93_898 ();
 sg13g2_decap_4 FILLER_0_93_906 ();
 sg13g2_fill_2 FILLER_0_93_910 ();
 sg13g2_fill_1 FILLER_0_93_921 ();
 sg13g2_decap_8 FILLER_0_93_926 ();
 sg13g2_fill_2 FILLER_0_93_933 ();
 sg13g2_decap_8 FILLER_0_93_976 ();
 sg13g2_decap_8 FILLER_0_93_983 ();
 sg13g2_decap_8 FILLER_0_93_990 ();
 sg13g2_decap_8 FILLER_0_93_997 ();
 sg13g2_decap_8 FILLER_0_93_1004 ();
 sg13g2_decap_8 FILLER_0_93_1011 ();
 sg13g2_decap_8 FILLER_0_93_1018 ();
 sg13g2_decap_8 FILLER_0_93_1025 ();
 sg13g2_decap_8 FILLER_0_93_1032 ();
 sg13g2_decap_8 FILLER_0_93_1039 ();
 sg13g2_decap_8 FILLER_0_93_1046 ();
 sg13g2_decap_8 FILLER_0_93_1053 ();
 sg13g2_decap_8 FILLER_0_93_1060 ();
 sg13g2_decap_8 FILLER_0_93_1067 ();
 sg13g2_decap_8 FILLER_0_93_1074 ();
 sg13g2_decap_8 FILLER_0_93_1081 ();
 sg13g2_decap_8 FILLER_0_93_1088 ();
 sg13g2_decap_8 FILLER_0_93_1095 ();
 sg13g2_decap_8 FILLER_0_93_1102 ();
 sg13g2_decap_8 FILLER_0_93_1109 ();
 sg13g2_decap_8 FILLER_0_93_1116 ();
 sg13g2_decap_8 FILLER_0_93_1123 ();
 sg13g2_decap_8 FILLER_0_93_1130 ();
 sg13g2_decap_8 FILLER_0_93_1137 ();
 sg13g2_decap_8 FILLER_0_93_1144 ();
 sg13g2_decap_8 FILLER_0_93_1151 ();
 sg13g2_decap_8 FILLER_0_93_1158 ();
 sg13g2_decap_8 FILLER_0_93_1165 ();
 sg13g2_decap_8 FILLER_0_93_1172 ();
 sg13g2_decap_8 FILLER_0_93_1179 ();
 sg13g2_decap_8 FILLER_0_93_1186 ();
 sg13g2_decap_8 FILLER_0_93_1193 ();
 sg13g2_decap_8 FILLER_0_93_1200 ();
 sg13g2_decap_8 FILLER_0_93_1207 ();
 sg13g2_decap_8 FILLER_0_93_1214 ();
 sg13g2_decap_8 FILLER_0_93_1221 ();
 sg13g2_decap_4 FILLER_0_94_0 ();
 sg13g2_fill_1 FILLER_0_94_4 ();
 sg13g2_decap_8 FILLER_0_94_45 ();
 sg13g2_decap_8 FILLER_0_94_52 ();
 sg13g2_decap_8 FILLER_0_94_59 ();
 sg13g2_fill_1 FILLER_0_94_66 ();
 sg13g2_decap_4 FILLER_0_94_72 ();
 sg13g2_fill_1 FILLER_0_94_76 ();
 sg13g2_decap_4 FILLER_0_94_117 ();
 sg13g2_fill_1 FILLER_0_94_121 ();
 sg13g2_fill_2 FILLER_0_94_163 ();
 sg13g2_fill_1 FILLER_0_94_165 ();
 sg13g2_fill_2 FILLER_0_94_170 ();
 sg13g2_fill_1 FILLER_0_94_172 ();
 sg13g2_decap_8 FILLER_0_94_177 ();
 sg13g2_fill_2 FILLER_0_94_184 ();
 sg13g2_decap_4 FILLER_0_94_190 ();
 sg13g2_fill_1 FILLER_0_94_194 ();
 sg13g2_fill_1 FILLER_0_94_200 ();
 sg13g2_decap_8 FILLER_0_94_209 ();
 sg13g2_fill_1 FILLER_0_94_225 ();
 sg13g2_fill_2 FILLER_0_94_236 ();
 sg13g2_fill_1 FILLER_0_94_242 ();
 sg13g2_fill_2 FILLER_0_94_269 ();
 sg13g2_decap_8 FILLER_0_94_276 ();
 sg13g2_fill_1 FILLER_0_94_283 ();
 sg13g2_fill_1 FILLER_0_94_310 ();
 sg13g2_decap_8 FILLER_0_94_326 ();
 sg13g2_decap_4 FILLER_0_94_333 ();
 sg13g2_fill_1 FILLER_0_94_347 ();
 sg13g2_decap_8 FILLER_0_94_383 ();
 sg13g2_decap_8 FILLER_0_94_390 ();
 sg13g2_fill_2 FILLER_0_94_397 ();
 sg13g2_fill_1 FILLER_0_94_399 ();
 sg13g2_fill_1 FILLER_0_94_420 ();
 sg13g2_decap_8 FILLER_0_94_471 ();
 sg13g2_fill_1 FILLER_0_94_478 ();
 sg13g2_decap_8 FILLER_0_94_494 ();
 sg13g2_decap_8 FILLER_0_94_501 ();
 sg13g2_decap_8 FILLER_0_94_508 ();
 sg13g2_decap_8 FILLER_0_94_515 ();
 sg13g2_decap_8 FILLER_0_94_522 ();
 sg13g2_decap_8 FILLER_0_94_529 ();
 sg13g2_decap_4 FILLER_0_94_536 ();
 sg13g2_fill_1 FILLER_0_94_540 ();
 sg13g2_decap_4 FILLER_0_94_550 ();
 sg13g2_fill_1 FILLER_0_94_558 ();
 sg13g2_fill_2 FILLER_0_94_569 ();
 sg13g2_fill_1 FILLER_0_94_571 ();
 sg13g2_decap_8 FILLER_0_94_580 ();
 sg13g2_fill_2 FILLER_0_94_587 ();
 sg13g2_fill_1 FILLER_0_94_601 ();
 sg13g2_fill_2 FILLER_0_94_617 ();
 sg13g2_fill_2 FILLER_0_94_645 ();
 sg13g2_fill_2 FILLER_0_94_655 ();
 sg13g2_fill_1 FILLER_0_94_657 ();
 sg13g2_decap_8 FILLER_0_94_662 ();
 sg13g2_decap_8 FILLER_0_94_669 ();
 sg13g2_decap_8 FILLER_0_94_676 ();
 sg13g2_decap_8 FILLER_0_94_683 ();
 sg13g2_decap_8 FILLER_0_94_690 ();
 sg13g2_decap_8 FILLER_0_94_697 ();
 sg13g2_decap_4 FILLER_0_94_713 ();
 sg13g2_fill_2 FILLER_0_94_717 ();
 sg13g2_decap_4 FILLER_0_94_729 ();
 sg13g2_fill_1 FILLER_0_94_733 ();
 sg13g2_decap_8 FILLER_0_94_769 ();
 sg13g2_decap_8 FILLER_0_94_776 ();
 sg13g2_decap_8 FILLER_0_94_783 ();
 sg13g2_decap_4 FILLER_0_94_790 ();
 sg13g2_decap_8 FILLER_0_94_824 ();
 sg13g2_decap_4 FILLER_0_94_831 ();
 sg13g2_fill_2 FILLER_0_94_835 ();
 sg13g2_fill_2 FILLER_0_94_868 ();
 sg13g2_fill_1 FILLER_0_94_870 ();
 sg13g2_decap_8 FILLER_0_94_897 ();
 sg13g2_fill_1 FILLER_0_94_904 ();
 sg13g2_decap_8 FILLER_0_94_936 ();
 sg13g2_decap_4 FILLER_0_94_948 ();
 sg13g2_fill_1 FILLER_0_94_952 ();
 sg13g2_decap_8 FILLER_0_94_957 ();
 sg13g2_fill_1 FILLER_0_94_964 ();
 sg13g2_decap_8 FILLER_0_94_973 ();
 sg13g2_decap_8 FILLER_0_94_980 ();
 sg13g2_decap_8 FILLER_0_94_987 ();
 sg13g2_decap_8 FILLER_0_94_994 ();
 sg13g2_decap_8 FILLER_0_94_1001 ();
 sg13g2_decap_8 FILLER_0_94_1008 ();
 sg13g2_decap_8 FILLER_0_94_1015 ();
 sg13g2_decap_8 FILLER_0_94_1022 ();
 sg13g2_decap_8 FILLER_0_94_1029 ();
 sg13g2_decap_8 FILLER_0_94_1036 ();
 sg13g2_decap_8 FILLER_0_94_1043 ();
 sg13g2_decap_8 FILLER_0_94_1050 ();
 sg13g2_decap_8 FILLER_0_94_1057 ();
 sg13g2_decap_8 FILLER_0_94_1064 ();
 sg13g2_decap_8 FILLER_0_94_1071 ();
 sg13g2_decap_8 FILLER_0_94_1078 ();
 sg13g2_decap_8 FILLER_0_94_1085 ();
 sg13g2_decap_8 FILLER_0_94_1092 ();
 sg13g2_decap_8 FILLER_0_94_1099 ();
 sg13g2_decap_8 FILLER_0_94_1106 ();
 sg13g2_decap_8 FILLER_0_94_1113 ();
 sg13g2_decap_8 FILLER_0_94_1120 ();
 sg13g2_decap_8 FILLER_0_94_1127 ();
 sg13g2_decap_8 FILLER_0_94_1134 ();
 sg13g2_decap_8 FILLER_0_94_1141 ();
 sg13g2_decap_8 FILLER_0_94_1148 ();
 sg13g2_decap_8 FILLER_0_94_1155 ();
 sg13g2_decap_8 FILLER_0_94_1162 ();
 sg13g2_decap_8 FILLER_0_94_1169 ();
 sg13g2_decap_8 FILLER_0_94_1176 ();
 sg13g2_decap_8 FILLER_0_94_1183 ();
 sg13g2_decap_8 FILLER_0_94_1190 ();
 sg13g2_decap_8 FILLER_0_94_1197 ();
 sg13g2_decap_8 FILLER_0_94_1204 ();
 sg13g2_decap_8 FILLER_0_94_1211 ();
 sg13g2_decap_8 FILLER_0_94_1218 ();
 sg13g2_fill_2 FILLER_0_94_1225 ();
 sg13g2_fill_1 FILLER_0_94_1227 ();
 sg13g2_fill_1 FILLER_0_95_0 ();
 sg13g2_decap_8 FILLER_0_95_42 ();
 sg13g2_decap_8 FILLER_0_95_49 ();
 sg13g2_decap_8 FILLER_0_95_56 ();
 sg13g2_decap_8 FILLER_0_95_63 ();
 sg13g2_fill_2 FILLER_0_95_70 ();
 sg13g2_fill_2 FILLER_0_95_77 ();
 sg13g2_fill_1 FILLER_0_95_79 ();
 sg13g2_fill_2 FILLER_0_95_94 ();
 sg13g2_fill_1 FILLER_0_95_96 ();
 sg13g2_decap_8 FILLER_0_95_112 ();
 sg13g2_decap_8 FILLER_0_95_129 ();
 sg13g2_fill_2 FILLER_0_95_136 ();
 sg13g2_fill_2 FILLER_0_95_169 ();
 sg13g2_fill_1 FILLER_0_95_179 ();
 sg13g2_fill_2 FILLER_0_95_185 ();
 sg13g2_decap_8 FILLER_0_95_202 ();
 sg13g2_decap_4 FILLER_0_95_209 ();
 sg13g2_fill_1 FILLER_0_95_213 ();
 sg13g2_decap_8 FILLER_0_95_240 ();
 sg13g2_fill_2 FILLER_0_95_277 ();
 sg13g2_decap_8 FILLER_0_95_314 ();
 sg13g2_decap_4 FILLER_0_95_321 ();
 sg13g2_fill_2 FILLER_0_95_325 ();
 sg13g2_decap_8 FILLER_0_95_373 ();
 sg13g2_decap_8 FILLER_0_95_380 ();
 sg13g2_fill_2 FILLER_0_95_387 ();
 sg13g2_fill_1 FILLER_0_95_389 ();
 sg13g2_decap_4 FILLER_0_95_431 ();
 sg13g2_fill_2 FILLER_0_95_435 ();
 sg13g2_decap_8 FILLER_0_95_472 ();
 sg13g2_fill_2 FILLER_0_95_479 ();
 sg13g2_decap_8 FILLER_0_95_507 ();
 sg13g2_decap_8 FILLER_0_95_514 ();
 sg13g2_decap_8 FILLER_0_95_521 ();
 sg13g2_decap_8 FILLER_0_95_528 ();
 sg13g2_decap_4 FILLER_0_95_535 ();
 sg13g2_decap_4 FILLER_0_95_565 ();
 sg13g2_fill_1 FILLER_0_95_569 ();
 sg13g2_fill_2 FILLER_0_95_580 ();
 sg13g2_decap_4 FILLER_0_95_625 ();
 sg13g2_fill_1 FILLER_0_95_629 ();
 sg13g2_decap_4 FILLER_0_95_640 ();
 sg13g2_fill_2 FILLER_0_95_644 ();
 sg13g2_decap_8 FILLER_0_95_677 ();
 sg13g2_decap_8 FILLER_0_95_684 ();
 sg13g2_decap_8 FILLER_0_95_691 ();
 sg13g2_fill_2 FILLER_0_95_698 ();
 sg13g2_fill_1 FILLER_0_95_700 ();
 sg13g2_decap_8 FILLER_0_95_732 ();
 sg13g2_decap_8 FILLER_0_95_739 ();
 sg13g2_fill_2 FILLER_0_95_746 ();
 sg13g2_decap_4 FILLER_0_95_788 ();
 sg13g2_decap_8 FILLER_0_95_821 ();
 sg13g2_decap_8 FILLER_0_95_828 ();
 sg13g2_decap_8 FILLER_0_95_835 ();
 sg13g2_decap_8 FILLER_0_95_842 ();
 sg13g2_fill_2 FILLER_0_95_849 ();
 sg13g2_fill_1 FILLER_0_95_851 ();
 sg13g2_fill_2 FILLER_0_95_867 ();
 sg13g2_fill_1 FILLER_0_95_869 ();
 sg13g2_fill_1 FILLER_0_95_875 ();
 sg13g2_decap_8 FILLER_0_95_886 ();
 sg13g2_decap_8 FILLER_0_95_980 ();
 sg13g2_fill_2 FILLER_0_95_987 ();
 sg13g2_decap_8 FILLER_0_95_993 ();
 sg13g2_decap_8 FILLER_0_95_1000 ();
 sg13g2_decap_8 FILLER_0_95_1015 ();
 sg13g2_decap_8 FILLER_0_95_1022 ();
 sg13g2_decap_8 FILLER_0_95_1029 ();
 sg13g2_decap_8 FILLER_0_95_1036 ();
 sg13g2_decap_8 FILLER_0_95_1043 ();
 sg13g2_decap_8 FILLER_0_95_1050 ();
 sg13g2_decap_8 FILLER_0_95_1057 ();
 sg13g2_decap_8 FILLER_0_95_1064 ();
 sg13g2_decap_8 FILLER_0_95_1071 ();
 sg13g2_decap_8 FILLER_0_95_1078 ();
 sg13g2_decap_8 FILLER_0_95_1085 ();
 sg13g2_decap_8 FILLER_0_95_1092 ();
 sg13g2_decap_8 FILLER_0_95_1099 ();
 sg13g2_decap_8 FILLER_0_95_1106 ();
 sg13g2_decap_8 FILLER_0_95_1113 ();
 sg13g2_decap_8 FILLER_0_95_1120 ();
 sg13g2_decap_8 FILLER_0_95_1127 ();
 sg13g2_decap_8 FILLER_0_95_1134 ();
 sg13g2_decap_8 FILLER_0_95_1141 ();
 sg13g2_decap_8 FILLER_0_95_1148 ();
 sg13g2_decap_8 FILLER_0_95_1155 ();
 sg13g2_decap_8 FILLER_0_95_1162 ();
 sg13g2_decap_8 FILLER_0_95_1169 ();
 sg13g2_decap_8 FILLER_0_95_1176 ();
 sg13g2_decap_8 FILLER_0_95_1183 ();
 sg13g2_decap_8 FILLER_0_95_1190 ();
 sg13g2_decap_8 FILLER_0_95_1197 ();
 sg13g2_decap_8 FILLER_0_95_1204 ();
 sg13g2_decap_8 FILLER_0_95_1211 ();
 sg13g2_decap_8 FILLER_0_95_1218 ();
 sg13g2_fill_2 FILLER_0_95_1225 ();
 sg13g2_fill_1 FILLER_0_95_1227 ();
 sg13g2_decap_8 FILLER_0_96_0 ();
 sg13g2_decap_4 FILLER_0_96_7 ();
 sg13g2_decap_8 FILLER_0_96_15 ();
 sg13g2_decap_4 FILLER_0_96_22 ();
 sg13g2_decap_8 FILLER_0_96_41 ();
 sg13g2_decap_4 FILLER_0_96_61 ();
 sg13g2_decap_8 FILLER_0_96_70 ();
 sg13g2_decap_8 FILLER_0_96_77 ();
 sg13g2_decap_8 FILLER_0_96_84 ();
 sg13g2_decap_4 FILLER_0_96_91 ();
 sg13g2_fill_2 FILLER_0_96_95 ();
 sg13g2_decap_8 FILLER_0_96_136 ();
 sg13g2_decap_8 FILLER_0_96_143 ();
 sg13g2_fill_2 FILLER_0_96_150 ();
 sg13g2_fill_1 FILLER_0_96_178 ();
 sg13g2_decap_8 FILLER_0_96_236 ();
 sg13g2_decap_8 FILLER_0_96_243 ();
 sg13g2_fill_2 FILLER_0_96_250 ();
 sg13g2_fill_1 FILLER_0_96_252 ();
 sg13g2_decap_8 FILLER_0_96_272 ();
 sg13g2_decap_8 FILLER_0_96_279 ();
 sg13g2_decap_4 FILLER_0_96_286 ();
 sg13g2_decap_4 FILLER_0_96_294 ();
 sg13g2_fill_1 FILLER_0_96_298 ();
 sg13g2_decap_4 FILLER_0_96_309 ();
 sg13g2_fill_2 FILLER_0_96_317 ();
 sg13g2_fill_1 FILLER_0_96_319 ();
 sg13g2_decap_4 FILLER_0_96_351 ();
 sg13g2_fill_1 FILLER_0_96_355 ();
 sg13g2_decap_8 FILLER_0_96_360 ();
 sg13g2_decap_8 FILLER_0_96_367 ();
 sg13g2_decap_8 FILLER_0_96_374 ();
 sg13g2_decap_4 FILLER_0_96_381 ();
 sg13g2_fill_2 FILLER_0_96_389 ();
 sg13g2_decap_8 FILLER_0_96_421 ();
 sg13g2_decap_8 FILLER_0_96_428 ();
 sg13g2_decap_8 FILLER_0_96_435 ();
 sg13g2_decap_8 FILLER_0_96_442 ();
 sg13g2_fill_1 FILLER_0_96_449 ();
 sg13g2_decap_4 FILLER_0_96_454 ();
 sg13g2_decap_8 FILLER_0_96_463 ();
 sg13g2_decap_8 FILLER_0_96_470 ();
 sg13g2_decap_8 FILLER_0_96_477 ();
 sg13g2_fill_2 FILLER_0_96_484 ();
 sg13g2_decap_8 FILLER_0_96_526 ();
 sg13g2_decap_4 FILLER_0_96_533 ();
 sg13g2_fill_2 FILLER_0_96_537 ();
 sg13g2_decap_8 FILLER_0_96_570 ();
 sg13g2_decap_8 FILLER_0_96_577 ();
 sg13g2_fill_2 FILLER_0_96_584 ();
 sg13g2_fill_1 FILLER_0_96_586 ();
 sg13g2_fill_1 FILLER_0_96_651 ();
 sg13g2_decap_8 FILLER_0_96_693 ();
 sg13g2_fill_2 FILLER_0_96_700 ();
 sg13g2_fill_1 FILLER_0_96_702 ();
 sg13g2_decap_8 FILLER_0_96_722 ();
 sg13g2_decap_8 FILLER_0_96_729 ();
 sg13g2_decap_8 FILLER_0_96_741 ();
 sg13g2_fill_2 FILLER_0_96_748 ();
 sg13g2_fill_1 FILLER_0_96_750 ();
 sg13g2_fill_2 FILLER_0_96_766 ();
 sg13g2_fill_2 FILLER_0_96_794 ();
 sg13g2_fill_1 FILLER_0_96_835 ();
 sg13g2_decap_8 FILLER_0_96_903 ();
 sg13g2_fill_2 FILLER_0_96_910 ();
 sg13g2_fill_1 FILLER_0_96_912 ();
 sg13g2_decap_8 FILLER_0_96_937 ();
 sg13g2_fill_2 FILLER_0_96_948 ();
 sg13g2_fill_1 FILLER_0_96_950 ();
 sg13g2_decap_8 FILLER_0_96_1025 ();
 sg13g2_decap_8 FILLER_0_96_1032 ();
 sg13g2_decap_8 FILLER_0_96_1039 ();
 sg13g2_decap_8 FILLER_0_96_1046 ();
 sg13g2_decap_8 FILLER_0_96_1053 ();
 sg13g2_decap_8 FILLER_0_96_1060 ();
 sg13g2_decap_8 FILLER_0_96_1067 ();
 sg13g2_decap_8 FILLER_0_96_1074 ();
 sg13g2_decap_8 FILLER_0_96_1081 ();
 sg13g2_decap_8 FILLER_0_96_1088 ();
 sg13g2_decap_8 FILLER_0_96_1095 ();
 sg13g2_decap_8 FILLER_0_96_1102 ();
 sg13g2_decap_8 FILLER_0_96_1109 ();
 sg13g2_decap_8 FILLER_0_96_1116 ();
 sg13g2_decap_8 FILLER_0_96_1123 ();
 sg13g2_decap_8 FILLER_0_96_1130 ();
 sg13g2_decap_8 FILLER_0_96_1137 ();
 sg13g2_decap_8 FILLER_0_96_1144 ();
 sg13g2_decap_8 FILLER_0_96_1151 ();
 sg13g2_decap_8 FILLER_0_96_1158 ();
 sg13g2_decap_8 FILLER_0_96_1165 ();
 sg13g2_decap_8 FILLER_0_96_1172 ();
 sg13g2_decap_8 FILLER_0_96_1179 ();
 sg13g2_decap_8 FILLER_0_96_1186 ();
 sg13g2_decap_8 FILLER_0_96_1193 ();
 sg13g2_decap_8 FILLER_0_96_1200 ();
 sg13g2_decap_8 FILLER_0_96_1207 ();
 sg13g2_decap_8 FILLER_0_96_1214 ();
 sg13g2_decap_8 FILLER_0_96_1221 ();
 sg13g2_decap_8 FILLER_0_97_0 ();
 sg13g2_decap_8 FILLER_0_97_7 ();
 sg13g2_fill_2 FILLER_0_97_14 ();
 sg13g2_fill_2 FILLER_0_97_42 ();
 sg13g2_fill_1 FILLER_0_97_44 ();
 sg13g2_decap_8 FILLER_0_97_81 ();
 sg13g2_decap_8 FILLER_0_97_88 ();
 sg13g2_decap_8 FILLER_0_97_95 ();
 sg13g2_decap_8 FILLER_0_97_102 ();
 sg13g2_fill_1 FILLER_0_97_119 ();
 sg13g2_fill_1 FILLER_0_97_124 ();
 sg13g2_decap_4 FILLER_0_97_135 ();
 sg13g2_fill_1 FILLER_0_97_139 ();
 sg13g2_fill_1 FILLER_0_97_145 ();
 sg13g2_fill_2 FILLER_0_97_172 ();
 sg13g2_fill_1 FILLER_0_97_225 ();
 sg13g2_fill_2 FILLER_0_97_230 ();
 sg13g2_decap_8 FILLER_0_97_242 ();
 sg13g2_decap_8 FILLER_0_97_249 ();
 sg13g2_decap_4 FILLER_0_97_256 ();
 sg13g2_fill_2 FILLER_0_97_260 ();
 sg13g2_decap_8 FILLER_0_97_267 ();
 sg13g2_decap_8 FILLER_0_97_274 ();
 sg13g2_decap_8 FILLER_0_97_281 ();
 sg13g2_fill_2 FILLER_0_97_288 ();
 sg13g2_fill_1 FILLER_0_97_290 ();
 sg13g2_decap_4 FILLER_0_97_296 ();
 sg13g2_fill_2 FILLER_0_97_300 ();
 sg13g2_fill_1 FILLER_0_97_312 ();
 sg13g2_decap_8 FILLER_0_97_347 ();
 sg13g2_decap_8 FILLER_0_97_358 ();
 sg13g2_fill_2 FILLER_0_97_365 ();
 sg13g2_decap_8 FILLER_0_97_417 ();
 sg13g2_decap_8 FILLER_0_97_424 ();
 sg13g2_decap_8 FILLER_0_97_431 ();
 sg13g2_fill_2 FILLER_0_97_438 ();
 sg13g2_fill_1 FILLER_0_97_440 ();
 sg13g2_decap_4 FILLER_0_97_493 ();
 sg13g2_fill_2 FILLER_0_97_502 ();
 sg13g2_fill_1 FILLER_0_97_504 ();
 sg13g2_fill_2 FILLER_0_97_531 ();
 sg13g2_fill_2 FILLER_0_97_538 ();
 sg13g2_fill_1 FILLER_0_97_540 ();
 sg13g2_fill_1 FILLER_0_97_549 ();
 sg13g2_decap_4 FILLER_0_97_585 ();
 sg13g2_fill_2 FILLER_0_97_597 ();
 sg13g2_decap_8 FILLER_0_97_613 ();
 sg13g2_decap_4 FILLER_0_97_620 ();
 sg13g2_fill_2 FILLER_0_97_624 ();
 sg13g2_fill_2 FILLER_0_97_650 ();
 sg13g2_fill_1 FILLER_0_97_652 ();
 sg13g2_fill_2 FILLER_0_97_658 ();
 sg13g2_fill_1 FILLER_0_97_660 ();
 sg13g2_fill_2 FILLER_0_97_665 ();
 sg13g2_fill_1 FILLER_0_97_667 ();
 sg13g2_decap_4 FILLER_0_97_694 ();
 sg13g2_fill_2 FILLER_0_97_724 ();
 sg13g2_fill_2 FILLER_0_97_770 ();
 sg13g2_fill_1 FILLER_0_97_772 ();
 sg13g2_fill_2 FILLER_0_97_782 ();
 sg13g2_decap_4 FILLER_0_97_794 ();
 sg13g2_decap_4 FILLER_0_97_803 ();
 sg13g2_fill_2 FILLER_0_97_811 ();
 sg13g2_fill_1 FILLER_0_97_813 ();
 sg13g2_decap_8 FILLER_0_97_824 ();
 sg13g2_decap_8 FILLER_0_97_831 ();
 sg13g2_decap_4 FILLER_0_97_838 ();
 sg13g2_decap_8 FILLER_0_97_850 ();
 sg13g2_fill_2 FILLER_0_97_857 ();
 sg13g2_fill_1 FILLER_0_97_904 ();
 sg13g2_decap_8 FILLER_0_97_936 ();
 sg13g2_decap_8 FILLER_0_97_943 ();
 sg13g2_fill_1 FILLER_0_97_950 ();
 sg13g2_decap_8 FILLER_0_97_1044 ();
 sg13g2_decap_8 FILLER_0_97_1051 ();
 sg13g2_decap_8 FILLER_0_97_1058 ();
 sg13g2_decap_8 FILLER_0_97_1065 ();
 sg13g2_decap_8 FILLER_0_97_1072 ();
 sg13g2_decap_8 FILLER_0_97_1079 ();
 sg13g2_decap_8 FILLER_0_97_1086 ();
 sg13g2_decap_8 FILLER_0_97_1093 ();
 sg13g2_decap_8 FILLER_0_97_1100 ();
 sg13g2_decap_8 FILLER_0_97_1107 ();
 sg13g2_decap_8 FILLER_0_97_1114 ();
 sg13g2_decap_8 FILLER_0_97_1121 ();
 sg13g2_decap_8 FILLER_0_97_1128 ();
 sg13g2_decap_8 FILLER_0_97_1135 ();
 sg13g2_decap_8 FILLER_0_97_1142 ();
 sg13g2_decap_8 FILLER_0_97_1149 ();
 sg13g2_decap_8 FILLER_0_97_1156 ();
 sg13g2_decap_8 FILLER_0_97_1163 ();
 sg13g2_decap_8 FILLER_0_97_1170 ();
 sg13g2_decap_8 FILLER_0_97_1177 ();
 sg13g2_decap_8 FILLER_0_97_1184 ();
 sg13g2_decap_8 FILLER_0_97_1191 ();
 sg13g2_decap_8 FILLER_0_97_1198 ();
 sg13g2_decap_8 FILLER_0_97_1205 ();
 sg13g2_decap_8 FILLER_0_97_1212 ();
 sg13g2_decap_8 FILLER_0_97_1219 ();
 sg13g2_fill_2 FILLER_0_97_1226 ();
 sg13g2_decap_8 FILLER_0_98_0 ();
 sg13g2_decap_8 FILLER_0_98_7 ();
 sg13g2_decap_8 FILLER_0_98_14 ();
 sg13g2_fill_2 FILLER_0_98_21 ();
 sg13g2_fill_1 FILLER_0_98_23 ();
 sg13g2_decap_8 FILLER_0_98_85 ();
 sg13g2_decap_4 FILLER_0_98_92 ();
 sg13g2_fill_1 FILLER_0_98_96 ();
 sg13g2_fill_1 FILLER_0_98_137 ();
 sg13g2_fill_2 FILLER_0_98_168 ();
 sg13g2_fill_1 FILLER_0_98_170 ();
 sg13g2_fill_1 FILLER_0_98_184 ();
 sg13g2_decap_8 FILLER_0_98_208 ();
 sg13g2_fill_2 FILLER_0_98_215 ();
 sg13g2_fill_1 FILLER_0_98_217 ();
 sg13g2_fill_2 FILLER_0_98_244 ();
 sg13g2_fill_1 FILLER_0_98_246 ();
 sg13g2_fill_1 FILLER_0_98_256 ();
 sg13g2_fill_1 FILLER_0_98_283 ();
 sg13g2_fill_1 FILLER_0_98_310 ();
 sg13g2_fill_1 FILLER_0_98_323 ();
 sg13g2_fill_2 FILLER_0_98_344 ();
 sg13g2_fill_1 FILLER_0_98_346 ();
 sg13g2_decap_8 FILLER_0_98_409 ();
 sg13g2_decap_4 FILLER_0_98_416 ();
 sg13g2_fill_2 FILLER_0_98_424 ();
 sg13g2_fill_1 FILLER_0_98_426 ();
 sg13g2_decap_8 FILLER_0_98_436 ();
 sg13g2_decap_8 FILLER_0_98_443 ();
 sg13g2_fill_2 FILLER_0_98_450 ();
 sg13g2_fill_2 FILLER_0_98_462 ();
 sg13g2_decap_4 FILLER_0_98_485 ();
 sg13g2_fill_2 FILLER_0_98_493 ();
 sg13g2_fill_2 FILLER_0_98_513 ();
 sg13g2_fill_1 FILLER_0_98_515 ();
 sg13g2_fill_1 FILLER_0_98_526 ();
 sg13g2_fill_1 FILLER_0_98_553 ();
 sg13g2_fill_1 FILLER_0_98_564 ();
 sg13g2_fill_1 FILLER_0_98_569 ();
 sg13g2_fill_1 FILLER_0_98_596 ();
 sg13g2_decap_8 FILLER_0_98_601 ();
 sg13g2_decap_4 FILLER_0_98_608 ();
 sg13g2_fill_2 FILLER_0_98_612 ();
 sg13g2_fill_2 FILLER_0_98_619 ();
 sg13g2_decap_8 FILLER_0_98_647 ();
 sg13g2_decap_8 FILLER_0_98_654 ();
 sg13g2_decap_8 FILLER_0_98_661 ();
 sg13g2_fill_2 FILLER_0_98_673 ();
 sg13g2_fill_2 FILLER_0_98_679 ();
 sg13g2_decap_4 FILLER_0_98_691 ();
 sg13g2_decap_4 FILLER_0_98_721 ();
 sg13g2_decap_8 FILLER_0_98_760 ();
 sg13g2_decap_4 FILLER_0_98_767 ();
 sg13g2_fill_1 FILLER_0_98_797 ();
 sg13g2_decap_8 FILLER_0_98_824 ();
 sg13g2_decap_4 FILLER_0_98_831 ();
 sg13g2_decap_8 FILLER_0_98_866 ();
 sg13g2_fill_1 FILLER_0_98_873 ();
 sg13g2_decap_8 FILLER_0_98_882 ();
 sg13g2_decap_4 FILLER_0_98_910 ();
 sg13g2_decap_8 FILLER_0_98_918 ();
 sg13g2_decap_8 FILLER_0_98_925 ();
 sg13g2_decap_4 FILLER_0_98_932 ();
 sg13g2_fill_2 FILLER_0_98_936 ();
 sg13g2_decap_8 FILLER_0_98_943 ();
 sg13g2_decap_8 FILLER_0_98_950 ();
 sg13g2_fill_1 FILLER_0_98_957 ();
 sg13g2_decap_8 FILLER_0_98_971 ();
 sg13g2_decap_4 FILLER_0_98_978 ();
 sg13g2_decap_8 FILLER_0_98_1012 ();
 sg13g2_fill_1 FILLER_0_98_1024 ();
 sg13g2_fill_1 FILLER_0_98_1029 ();
 sg13g2_fill_2 FILLER_0_98_1040 ();
 sg13g2_decap_8 FILLER_0_98_1046 ();
 sg13g2_decap_8 FILLER_0_98_1053 ();
 sg13g2_decap_8 FILLER_0_98_1060 ();
 sg13g2_decap_8 FILLER_0_98_1067 ();
 sg13g2_decap_8 FILLER_0_98_1074 ();
 sg13g2_decap_8 FILLER_0_98_1081 ();
 sg13g2_decap_8 FILLER_0_98_1088 ();
 sg13g2_decap_8 FILLER_0_98_1095 ();
 sg13g2_decap_8 FILLER_0_98_1102 ();
 sg13g2_decap_8 FILLER_0_98_1109 ();
 sg13g2_decap_8 FILLER_0_98_1116 ();
 sg13g2_decap_8 FILLER_0_98_1123 ();
 sg13g2_decap_8 FILLER_0_98_1130 ();
 sg13g2_decap_8 FILLER_0_98_1137 ();
 sg13g2_decap_8 FILLER_0_98_1144 ();
 sg13g2_decap_8 FILLER_0_98_1151 ();
 sg13g2_decap_8 FILLER_0_98_1158 ();
 sg13g2_decap_8 FILLER_0_98_1165 ();
 sg13g2_decap_8 FILLER_0_98_1172 ();
 sg13g2_decap_8 FILLER_0_98_1179 ();
 sg13g2_decap_8 FILLER_0_98_1186 ();
 sg13g2_decap_8 FILLER_0_98_1193 ();
 sg13g2_decap_8 FILLER_0_98_1200 ();
 sg13g2_decap_8 FILLER_0_98_1207 ();
 sg13g2_decap_8 FILLER_0_98_1214 ();
 sg13g2_decap_8 FILLER_0_98_1221 ();
 sg13g2_decap_8 FILLER_0_99_0 ();
 sg13g2_decap_8 FILLER_0_99_7 ();
 sg13g2_decap_8 FILLER_0_99_14 ();
 sg13g2_decap_8 FILLER_0_99_21 ();
 sg13g2_fill_1 FILLER_0_99_33 ();
 sg13g2_fill_1 FILLER_0_99_38 ();
 sg13g2_fill_1 FILLER_0_99_49 ();
 sg13g2_fill_2 FILLER_0_99_60 ();
 sg13g2_decap_8 FILLER_0_99_96 ();
 sg13g2_decap_4 FILLER_0_99_103 ();
 sg13g2_fill_1 FILLER_0_99_107 ();
 sg13g2_decap_4 FILLER_0_99_134 ();
 sg13g2_decap_4 FILLER_0_99_143 ();
 sg13g2_fill_1 FILLER_0_99_147 ();
 sg13g2_fill_1 FILLER_0_99_152 ();
 sg13g2_fill_2 FILLER_0_99_173 ();
 sg13g2_decap_8 FILLER_0_99_206 ();
 sg13g2_fill_1 FILLER_0_99_213 ();
 sg13g2_fill_2 FILLER_0_99_250 ();
 sg13g2_fill_1 FILLER_0_99_282 ();
 sg13g2_decap_8 FILLER_0_99_301 ();
 sg13g2_decap_4 FILLER_0_99_308 ();
 sg13g2_fill_2 FILLER_0_99_312 ();
 sg13g2_fill_1 FILLER_0_99_340 ();
 sg13g2_fill_2 FILLER_0_99_346 ();
 sg13g2_fill_1 FILLER_0_99_353 ();
 sg13g2_fill_2 FILLER_0_99_359 ();
 sg13g2_fill_2 FILLER_0_99_394 ();
 sg13g2_decap_4 FILLER_0_99_404 ();
 sg13g2_fill_2 FILLER_0_99_455 ();
 sg13g2_decap_8 FILLER_0_99_501 ();
 sg13g2_fill_2 FILLER_0_99_508 ();
 sg13g2_fill_1 FILLER_0_99_543 ();
 sg13g2_decap_8 FILLER_0_99_552 ();
 sg13g2_decap_8 FILLER_0_99_559 ();
 sg13g2_fill_2 FILLER_0_99_566 ();
 sg13g2_fill_1 FILLER_0_99_568 ();
 sg13g2_fill_2 FILLER_0_99_584 ();
 sg13g2_fill_1 FILLER_0_99_586 ();
 sg13g2_decap_8 FILLER_0_99_597 ();
 sg13g2_decap_8 FILLER_0_99_604 ();
 sg13g2_decap_8 FILLER_0_99_611 ();
 sg13g2_decap_8 FILLER_0_99_618 ();
 sg13g2_fill_2 FILLER_0_99_625 ();
 sg13g2_decap_8 FILLER_0_99_631 ();
 sg13g2_decap_4 FILLER_0_99_638 ();
 sg13g2_fill_1 FILLER_0_99_642 ();
 sg13g2_decap_8 FILLER_0_99_658 ();
 sg13g2_decap_8 FILLER_0_99_665 ();
 sg13g2_fill_1 FILLER_0_99_686 ();
 sg13g2_decap_8 FILLER_0_99_695 ();
 sg13g2_fill_1 FILLER_0_99_711 ();
 sg13g2_fill_1 FILLER_0_99_722 ();
 sg13g2_fill_1 FILLER_0_99_733 ();
 sg13g2_fill_1 FILLER_0_99_738 ();
 sg13g2_fill_1 FILLER_0_99_765 ();
 sg13g2_decap_8 FILLER_0_99_800 ();
 sg13g2_fill_2 FILLER_0_99_807 ();
 sg13g2_decap_8 FILLER_0_99_828 ();
 sg13g2_decap_8 FILLER_0_99_835 ();
 sg13g2_decap_8 FILLER_0_99_842 ();
 sg13g2_decap_8 FILLER_0_99_849 ();
 sg13g2_decap_8 FILLER_0_99_856 ();
 sg13g2_decap_8 FILLER_0_99_863 ();
 sg13g2_decap_8 FILLER_0_99_870 ();
 sg13g2_decap_8 FILLER_0_99_877 ();
 sg13g2_fill_1 FILLER_0_99_884 ();
 sg13g2_fill_1 FILLER_0_99_890 ();
 sg13g2_decap_8 FILLER_0_99_971 ();
 sg13g2_decap_8 FILLER_0_99_978 ();
 sg13g2_decap_4 FILLER_0_99_985 ();
 sg13g2_fill_1 FILLER_0_99_989 ();
 sg13g2_fill_2 FILLER_0_99_1001 ();
 sg13g2_decap_8 FILLER_0_99_1007 ();
 sg13g2_fill_2 FILLER_0_99_1014 ();
 sg13g2_decap_4 FILLER_0_99_1021 ();
 sg13g2_fill_1 FILLER_0_99_1025 ();
 sg13g2_decap_8 FILLER_0_99_1057 ();
 sg13g2_decap_8 FILLER_0_99_1064 ();
 sg13g2_decap_8 FILLER_0_99_1071 ();
 sg13g2_decap_8 FILLER_0_99_1078 ();
 sg13g2_decap_8 FILLER_0_99_1085 ();
 sg13g2_decap_8 FILLER_0_99_1092 ();
 sg13g2_decap_8 FILLER_0_99_1099 ();
 sg13g2_decap_8 FILLER_0_99_1106 ();
 sg13g2_decap_8 FILLER_0_99_1113 ();
 sg13g2_decap_8 FILLER_0_99_1120 ();
 sg13g2_decap_8 FILLER_0_99_1127 ();
 sg13g2_decap_8 FILLER_0_99_1134 ();
 sg13g2_decap_8 FILLER_0_99_1141 ();
 sg13g2_decap_8 FILLER_0_99_1148 ();
 sg13g2_decap_8 FILLER_0_99_1155 ();
 sg13g2_decap_8 FILLER_0_99_1162 ();
 sg13g2_decap_8 FILLER_0_99_1169 ();
 sg13g2_decap_8 FILLER_0_99_1176 ();
 sg13g2_decap_8 FILLER_0_99_1183 ();
 sg13g2_decap_8 FILLER_0_99_1190 ();
 sg13g2_decap_8 FILLER_0_99_1197 ();
 sg13g2_decap_8 FILLER_0_99_1204 ();
 sg13g2_decap_8 FILLER_0_99_1211 ();
 sg13g2_decap_8 FILLER_0_99_1218 ();
 sg13g2_fill_2 FILLER_0_99_1225 ();
 sg13g2_fill_1 FILLER_0_99_1227 ();
 sg13g2_decap_8 FILLER_0_100_0 ();
 sg13g2_decap_8 FILLER_0_100_7 ();
 sg13g2_decap_8 FILLER_0_100_14 ();
 sg13g2_decap_8 FILLER_0_100_21 ();
 sg13g2_decap_8 FILLER_0_100_28 ();
 sg13g2_decap_8 FILLER_0_100_35 ();
 sg13g2_decap_8 FILLER_0_100_42 ();
 sg13g2_decap_8 FILLER_0_100_86 ();
 sg13g2_decap_8 FILLER_0_100_93 ();
 sg13g2_decap_8 FILLER_0_100_100 ();
 sg13g2_fill_1 FILLER_0_100_107 ();
 sg13g2_decap_4 FILLER_0_100_113 ();
 sg13g2_fill_1 FILLER_0_100_121 ();
 sg13g2_fill_2 FILLER_0_100_132 ();
 sg13g2_fill_1 FILLER_0_100_134 ();
 sg13g2_decap_8 FILLER_0_100_174 ();
 sg13g2_fill_2 FILLER_0_100_181 ();
 sg13g2_decap_8 FILLER_0_100_202 ();
 sg13g2_decap_4 FILLER_0_100_209 ();
 sg13g2_fill_1 FILLER_0_100_216 ();
 sg13g2_decap_8 FILLER_0_100_221 ();
 sg13g2_decap_4 FILLER_0_100_242 ();
 sg13g2_fill_1 FILLER_0_100_266 ();
 sg13g2_fill_2 FILLER_0_100_272 ();
 sg13g2_decap_8 FILLER_0_100_300 ();
 sg13g2_decap_8 FILLER_0_100_307 ();
 sg13g2_decap_4 FILLER_0_100_314 ();
 sg13g2_fill_1 FILLER_0_100_318 ();
 sg13g2_fill_2 FILLER_0_100_331 ();
 sg13g2_fill_1 FILLER_0_100_333 ();
 sg13g2_fill_2 FILLER_0_100_344 ();
 sg13g2_fill_1 FILLER_0_100_350 ();
 sg13g2_decap_8 FILLER_0_100_377 ();
 sg13g2_fill_1 FILLER_0_100_409 ();
 sg13g2_fill_2 FILLER_0_100_420 ();
 sg13g2_decap_8 FILLER_0_100_493 ();
 sg13g2_fill_2 FILLER_0_100_500 ();
 sg13g2_decap_8 FILLER_0_100_512 ();
 sg13g2_fill_2 FILLER_0_100_519 ();
 sg13g2_fill_1 FILLER_0_100_521 ();
 sg13g2_decap_4 FILLER_0_100_548 ();
 sg13g2_decap_8 FILLER_0_100_556 ();
 sg13g2_decap_8 FILLER_0_100_563 ();
 sg13g2_decap_4 FILLER_0_100_570 ();
 sg13g2_fill_1 FILLER_0_100_574 ();
 sg13g2_decap_8 FILLER_0_100_611 ();
 sg13g2_fill_2 FILLER_0_100_618 ();
 sg13g2_decap_4 FILLER_0_100_651 ();
 sg13g2_fill_2 FILLER_0_100_655 ();
 sg13g2_decap_8 FILLER_0_100_697 ();
 sg13g2_decap_8 FILLER_0_100_704 ();
 sg13g2_decap_4 FILLER_0_100_711 ();
 sg13g2_fill_2 FILLER_0_100_715 ();
 sg13g2_decap_8 FILLER_0_100_722 ();
 sg13g2_fill_2 FILLER_0_100_729 ();
 sg13g2_fill_1 FILLER_0_100_731 ();
 sg13g2_fill_2 FILLER_0_100_755 ();
 sg13g2_fill_2 FILLER_0_100_767 ();
 sg13g2_fill_1 FILLER_0_100_769 ();
 sg13g2_decap_8 FILLER_0_100_785 ();
 sg13g2_decap_8 FILLER_0_100_792 ();
 sg13g2_decap_8 FILLER_0_100_799 ();
 sg13g2_fill_2 FILLER_0_100_806 ();
 sg13g2_decap_8 FILLER_0_100_834 ();
 sg13g2_decap_8 FILLER_0_100_841 ();
 sg13g2_fill_2 FILLER_0_100_853 ();
 sg13g2_fill_1 FILLER_0_100_855 ();
 sg13g2_decap_8 FILLER_0_100_860 ();
 sg13g2_decap_8 FILLER_0_100_867 ();
 sg13g2_fill_2 FILLER_0_100_874 ();
 sg13g2_fill_1 FILLER_0_100_876 ();
 sg13g2_decap_4 FILLER_0_100_917 ();
 sg13g2_fill_1 FILLER_0_100_921 ();
 sg13g2_fill_1 FILLER_0_100_953 ();
 sg13g2_fill_1 FILLER_0_100_980 ();
 sg13g2_fill_1 FILLER_0_100_1007 ();
 sg13g2_fill_2 FILLER_0_100_1028 ();
 sg13g2_fill_1 FILLER_0_100_1040 ();
 sg13g2_decap_8 FILLER_0_100_1045 ();
 sg13g2_decap_8 FILLER_0_100_1052 ();
 sg13g2_decap_8 FILLER_0_100_1059 ();
 sg13g2_decap_8 FILLER_0_100_1066 ();
 sg13g2_decap_8 FILLER_0_100_1073 ();
 sg13g2_decap_8 FILLER_0_100_1080 ();
 sg13g2_decap_8 FILLER_0_100_1087 ();
 sg13g2_decap_8 FILLER_0_100_1094 ();
 sg13g2_decap_8 FILLER_0_100_1101 ();
 sg13g2_decap_8 FILLER_0_100_1108 ();
 sg13g2_decap_8 FILLER_0_100_1115 ();
 sg13g2_decap_8 FILLER_0_100_1122 ();
 sg13g2_decap_8 FILLER_0_100_1129 ();
 sg13g2_decap_8 FILLER_0_100_1136 ();
 sg13g2_decap_8 FILLER_0_100_1143 ();
 sg13g2_decap_8 FILLER_0_100_1150 ();
 sg13g2_decap_8 FILLER_0_100_1157 ();
 sg13g2_decap_8 FILLER_0_100_1164 ();
 sg13g2_decap_8 FILLER_0_100_1171 ();
 sg13g2_decap_8 FILLER_0_100_1178 ();
 sg13g2_decap_8 FILLER_0_100_1185 ();
 sg13g2_decap_8 FILLER_0_100_1192 ();
 sg13g2_decap_8 FILLER_0_100_1199 ();
 sg13g2_decap_8 FILLER_0_100_1206 ();
 sg13g2_decap_8 FILLER_0_100_1213 ();
 sg13g2_decap_8 FILLER_0_100_1220 ();
 sg13g2_fill_1 FILLER_0_100_1227 ();
 sg13g2_decap_8 FILLER_0_101_0 ();
 sg13g2_decap_8 FILLER_0_101_7 ();
 sg13g2_decap_8 FILLER_0_101_14 ();
 sg13g2_decap_8 FILLER_0_101_21 ();
 sg13g2_decap_8 FILLER_0_101_28 ();
 sg13g2_decap_8 FILLER_0_101_35 ();
 sg13g2_decap_8 FILLER_0_101_42 ();
 sg13g2_decap_8 FILLER_0_101_49 ();
 sg13g2_fill_1 FILLER_0_101_56 ();
 sg13g2_decap_8 FILLER_0_101_88 ();
 sg13g2_decap_8 FILLER_0_101_95 ();
 sg13g2_decap_4 FILLER_0_101_102 ();
 sg13g2_decap_8 FILLER_0_101_137 ();
 sg13g2_decap_4 FILLER_0_101_144 ();
 sg13g2_fill_1 FILLER_0_101_148 ();
 sg13g2_decap_8 FILLER_0_101_164 ();
 sg13g2_decap_8 FILLER_0_101_171 ();
 sg13g2_decap_8 FILLER_0_101_178 ();
 sg13g2_fill_1 FILLER_0_101_185 ();
 sg13g2_fill_1 FILLER_0_101_212 ();
 sg13g2_fill_2 FILLER_0_101_225 ();
 sg13g2_fill_1 FILLER_0_101_227 ();
 sg13g2_decap_4 FILLER_0_101_242 ();
 sg13g2_fill_1 FILLER_0_101_246 ();
 sg13g2_fill_2 FILLER_0_101_255 ();
 sg13g2_fill_1 FILLER_0_101_257 ();
 sg13g2_decap_8 FILLER_0_101_262 ();
 sg13g2_decap_4 FILLER_0_101_269 ();
 sg13g2_fill_2 FILLER_0_101_273 ();
 sg13g2_decap_4 FILLER_0_101_280 ();
 sg13g2_fill_2 FILLER_0_101_284 ();
 sg13g2_decap_8 FILLER_0_101_300 ();
 sg13g2_decap_8 FILLER_0_101_307 ();
 sg13g2_decap_8 FILLER_0_101_345 ();
 sg13g2_decap_8 FILLER_0_101_352 ();
 sg13g2_fill_2 FILLER_0_101_359 ();
 sg13g2_fill_1 FILLER_0_101_370 ();
 sg13g2_fill_1 FILLER_0_101_437 ();
 sg13g2_fill_2 FILLER_0_101_442 ();
 sg13g2_fill_2 FILLER_0_101_454 ();
 sg13g2_fill_1 FILLER_0_101_456 ();
 sg13g2_decap_4 FILLER_0_101_467 ();
 sg13g2_decap_8 FILLER_0_101_475 ();
 sg13g2_decap_8 FILLER_0_101_482 ();
 sg13g2_decap_4 FILLER_0_101_489 ();
 sg13g2_fill_1 FILLER_0_101_493 ();
 sg13g2_decap_4 FILLER_0_101_504 ();
 sg13g2_fill_1 FILLER_0_101_508 ();
 sg13g2_decap_4 FILLER_0_101_571 ();
 sg13g2_decap_4 FILLER_0_101_652 ();
 sg13g2_decap_8 FILLER_0_101_692 ();
 sg13g2_decap_8 FILLER_0_101_699 ();
 sg13g2_decap_8 FILLER_0_101_706 ();
 sg13g2_decap_8 FILLER_0_101_713 ();
 sg13g2_decap_8 FILLER_0_101_720 ();
 sg13g2_decap_4 FILLER_0_101_727 ();
 sg13g2_fill_1 FILLER_0_101_731 ();
 sg13g2_decap_8 FILLER_0_101_752 ();
 sg13g2_fill_1 FILLER_0_101_759 ();
 sg13g2_decap_8 FILLER_0_101_771 ();
 sg13g2_decap_8 FILLER_0_101_778 ();
 sg13g2_decap_8 FILLER_0_101_785 ();
 sg13g2_decap_8 FILLER_0_101_792 ();
 sg13g2_decap_8 FILLER_0_101_799 ();
 sg13g2_decap_8 FILLER_0_101_806 ();
 sg13g2_fill_1 FILLER_0_101_844 ();
 sg13g2_decap_8 FILLER_0_101_871 ();
 sg13g2_decap_8 FILLER_0_101_878 ();
 sg13g2_fill_1 FILLER_0_101_885 ();
 sg13g2_fill_1 FILLER_0_101_890 ();
 sg13g2_fill_1 FILLER_0_101_917 ();
 sg13g2_fill_1 FILLER_0_101_944 ();
 sg13g2_fill_2 FILLER_0_101_955 ();
 sg13g2_fill_1 FILLER_0_101_983 ();
 sg13g2_fill_2 FILLER_0_101_1020 ();
 sg13g2_decap_8 FILLER_0_101_1053 ();
 sg13g2_decap_8 FILLER_0_101_1060 ();
 sg13g2_decap_8 FILLER_0_101_1067 ();
 sg13g2_decap_8 FILLER_0_101_1074 ();
 sg13g2_decap_8 FILLER_0_101_1081 ();
 sg13g2_decap_8 FILLER_0_101_1088 ();
 sg13g2_decap_8 FILLER_0_101_1095 ();
 sg13g2_decap_8 FILLER_0_101_1102 ();
 sg13g2_decap_8 FILLER_0_101_1109 ();
 sg13g2_decap_8 FILLER_0_101_1116 ();
 sg13g2_decap_8 FILLER_0_101_1123 ();
 sg13g2_decap_8 FILLER_0_101_1130 ();
 sg13g2_decap_8 FILLER_0_101_1137 ();
 sg13g2_decap_8 FILLER_0_101_1144 ();
 sg13g2_decap_8 FILLER_0_101_1151 ();
 sg13g2_decap_8 FILLER_0_101_1158 ();
 sg13g2_decap_8 FILLER_0_101_1165 ();
 sg13g2_decap_8 FILLER_0_101_1172 ();
 sg13g2_decap_8 FILLER_0_101_1179 ();
 sg13g2_decap_8 FILLER_0_101_1186 ();
 sg13g2_decap_8 FILLER_0_101_1193 ();
 sg13g2_decap_8 FILLER_0_101_1200 ();
 sg13g2_decap_8 FILLER_0_101_1207 ();
 sg13g2_decap_8 FILLER_0_101_1214 ();
 sg13g2_decap_8 FILLER_0_101_1221 ();
 sg13g2_decap_8 FILLER_0_102_0 ();
 sg13g2_decap_8 FILLER_0_102_7 ();
 sg13g2_decap_8 FILLER_0_102_14 ();
 sg13g2_decap_8 FILLER_0_102_21 ();
 sg13g2_decap_8 FILLER_0_102_28 ();
 sg13g2_decap_8 FILLER_0_102_35 ();
 sg13g2_decap_8 FILLER_0_102_42 ();
 sg13g2_fill_2 FILLER_0_102_49 ();
 sg13g2_fill_1 FILLER_0_102_51 ();
 sg13g2_decap_8 FILLER_0_102_62 ();
 sg13g2_fill_1 FILLER_0_102_69 ();
 sg13g2_decap_8 FILLER_0_102_74 ();
 sg13g2_decap_8 FILLER_0_102_81 ();
 sg13g2_decap_8 FILLER_0_102_88 ();
 sg13g2_fill_1 FILLER_0_102_112 ();
 sg13g2_fill_1 FILLER_0_102_117 ();
 sg13g2_fill_1 FILLER_0_102_128 ();
 sg13g2_fill_2 FILLER_0_102_139 ();
 sg13g2_decap_8 FILLER_0_102_171 ();
 sg13g2_fill_2 FILLER_0_102_178 ();
 sg13g2_fill_1 FILLER_0_102_211 ();
 sg13g2_decap_8 FILLER_0_102_243 ();
 sg13g2_decap_4 FILLER_0_102_250 ();
 sg13g2_fill_1 FILLER_0_102_259 ();
 sg13g2_fill_2 FILLER_0_102_277 ();
 sg13g2_fill_1 FILLER_0_102_279 ();
 sg13g2_decap_8 FILLER_0_102_306 ();
 sg13g2_fill_2 FILLER_0_102_313 ();
 sg13g2_decap_4 FILLER_0_102_346 ();
 sg13g2_fill_2 FILLER_0_102_350 ();
 sg13g2_decap_4 FILLER_0_102_378 ();
 sg13g2_fill_2 FILLER_0_102_423 ();
 sg13g2_decap_8 FILLER_0_102_438 ();
 sg13g2_decap_8 FILLER_0_102_445 ();
 sg13g2_decap_4 FILLER_0_102_452 ();
 sg13g2_fill_1 FILLER_0_102_456 ();
 sg13g2_decap_8 FILLER_0_102_462 ();
 sg13g2_decap_8 FILLER_0_102_469 ();
 sg13g2_fill_1 FILLER_0_102_476 ();
 sg13g2_decap_8 FILLER_0_102_482 ();
 sg13g2_fill_2 FILLER_0_102_489 ();
 sg13g2_fill_1 FILLER_0_102_491 ();
 sg13g2_fill_1 FILLER_0_102_496 ();
 sg13g2_fill_1 FILLER_0_102_502 ();
 sg13g2_fill_2 FILLER_0_102_529 ();
 sg13g2_fill_1 FILLER_0_102_545 ();
 sg13g2_fill_1 FILLER_0_102_551 ();
 sg13g2_fill_1 FILLER_0_102_562 ();
 sg13g2_fill_1 FILLER_0_102_567 ();
 sg13g2_fill_1 FILLER_0_102_617 ();
 sg13g2_decap_4 FILLER_0_102_622 ();
 sg13g2_fill_1 FILLER_0_102_626 ();
 sg13g2_fill_1 FILLER_0_102_636 ();
 sg13g2_fill_2 FILLER_0_102_647 ();
 sg13g2_fill_1 FILLER_0_102_649 ();
 sg13g2_decap_4 FILLER_0_102_680 ();
 sg13g2_fill_1 FILLER_0_102_684 ();
 sg13g2_decap_4 FILLER_0_102_720 ();
 sg13g2_fill_1 FILLER_0_102_724 ();
 sg13g2_fill_2 FILLER_0_102_756 ();
 sg13g2_fill_1 FILLER_0_102_758 ();
 sg13g2_decap_8 FILLER_0_102_785 ();
 sg13g2_decap_8 FILLER_0_102_792 ();
 sg13g2_decap_8 FILLER_0_102_799 ();
 sg13g2_decap_4 FILLER_0_102_806 ();
 sg13g2_fill_2 FILLER_0_102_815 ();
 sg13g2_fill_1 FILLER_0_102_817 ();
 sg13g2_fill_2 FILLER_0_102_828 ();
 sg13g2_fill_1 FILLER_0_102_830 ();
 sg13g2_fill_2 FILLER_0_102_857 ();
 sg13g2_fill_1 FILLER_0_102_859 ();
 sg13g2_fill_1 FILLER_0_102_886 ();
 sg13g2_decap_4 FILLER_0_102_910 ();
 sg13g2_fill_2 FILLER_0_102_914 ();
 sg13g2_decap_4 FILLER_0_102_921 ();
 sg13g2_fill_2 FILLER_0_102_929 ();
 sg13g2_fill_1 FILLER_0_102_931 ();
 sg13g2_decap_8 FILLER_0_102_936 ();
 sg13g2_decap_4 FILLER_0_102_943 ();
 sg13g2_decap_4 FILLER_0_102_951 ();
 sg13g2_decap_8 FILLER_0_102_1050 ();
 sg13g2_decap_8 FILLER_0_102_1057 ();
 sg13g2_decap_8 FILLER_0_102_1064 ();
 sg13g2_decap_8 FILLER_0_102_1071 ();
 sg13g2_decap_8 FILLER_0_102_1078 ();
 sg13g2_decap_8 FILLER_0_102_1085 ();
 sg13g2_decap_8 FILLER_0_102_1092 ();
 sg13g2_decap_8 FILLER_0_102_1099 ();
 sg13g2_decap_8 FILLER_0_102_1106 ();
 sg13g2_decap_8 FILLER_0_102_1113 ();
 sg13g2_decap_8 FILLER_0_102_1120 ();
 sg13g2_decap_8 FILLER_0_102_1127 ();
 sg13g2_decap_8 FILLER_0_102_1134 ();
 sg13g2_decap_8 FILLER_0_102_1141 ();
 sg13g2_decap_8 FILLER_0_102_1148 ();
 sg13g2_decap_8 FILLER_0_102_1155 ();
 sg13g2_decap_8 FILLER_0_102_1162 ();
 sg13g2_decap_8 FILLER_0_102_1169 ();
 sg13g2_decap_8 FILLER_0_102_1176 ();
 sg13g2_decap_8 FILLER_0_102_1183 ();
 sg13g2_decap_8 FILLER_0_102_1190 ();
 sg13g2_decap_8 FILLER_0_102_1197 ();
 sg13g2_decap_8 FILLER_0_102_1204 ();
 sg13g2_decap_8 FILLER_0_102_1211 ();
 sg13g2_decap_8 FILLER_0_102_1218 ();
 sg13g2_fill_2 FILLER_0_102_1225 ();
 sg13g2_fill_1 FILLER_0_102_1227 ();
 sg13g2_decap_8 FILLER_0_103_0 ();
 sg13g2_decap_8 FILLER_0_103_7 ();
 sg13g2_decap_8 FILLER_0_103_14 ();
 sg13g2_decap_8 FILLER_0_103_21 ();
 sg13g2_decap_8 FILLER_0_103_28 ();
 sg13g2_decap_8 FILLER_0_103_35 ();
 sg13g2_decap_8 FILLER_0_103_42 ();
 sg13g2_decap_8 FILLER_0_103_49 ();
 sg13g2_fill_1 FILLER_0_103_56 ();
 sg13g2_decap_8 FILLER_0_103_88 ();
 sg13g2_decap_8 FILLER_0_103_95 ();
 sg13g2_fill_1 FILLER_0_103_102 ();
 sg13g2_decap_8 FILLER_0_103_134 ();
 sg13g2_fill_2 FILLER_0_103_172 ();
 sg13g2_fill_2 FILLER_0_103_183 ();
 sg13g2_fill_1 FILLER_0_103_185 ();
 sg13g2_fill_2 FILLER_0_103_210 ();
 sg13g2_fill_1 FILLER_0_103_212 ();
 sg13g2_decap_4 FILLER_0_103_249 ();
 sg13g2_decap_8 FILLER_0_103_279 ();
 sg13g2_fill_2 FILLER_0_103_286 ();
 sg13g2_decap_8 FILLER_0_103_307 ();
 sg13g2_decap_8 FILLER_0_103_314 ();
 sg13g2_fill_2 FILLER_0_103_325 ();
 sg13g2_fill_1 FILLER_0_103_348 ();
 sg13g2_fill_1 FILLER_0_103_379 ();
 sg13g2_fill_1 FILLER_0_103_388 ();
 sg13g2_decap_4 FILLER_0_103_408 ();
 sg13g2_fill_2 FILLER_0_103_412 ();
 sg13g2_decap_8 FILLER_0_103_449 ();
 sg13g2_decap_8 FILLER_0_103_456 ();
 sg13g2_decap_8 FILLER_0_103_463 ();
 sg13g2_fill_1 FILLER_0_103_470 ();
 sg13g2_decap_8 FILLER_0_103_515 ();
 sg13g2_decap_8 FILLER_0_103_522 ();
 sg13g2_fill_1 FILLER_0_103_529 ();
 sg13g2_fill_1 FILLER_0_103_542 ();
 sg13g2_decap_8 FILLER_0_103_569 ();
 sg13g2_decap_8 FILLER_0_103_576 ();
 sg13g2_decap_8 FILLER_0_103_583 ();
 sg13g2_fill_1 FILLER_0_103_594 ();
 sg13g2_decap_8 FILLER_0_103_599 ();
 sg13g2_decap_8 FILLER_0_103_606 ();
 sg13g2_decap_8 FILLER_0_103_613 ();
 sg13g2_decap_4 FILLER_0_103_620 ();
 sg13g2_fill_2 FILLER_0_103_624 ();
 sg13g2_fill_2 FILLER_0_103_652 ();
 sg13g2_decap_8 FILLER_0_103_682 ();
 sg13g2_fill_2 FILLER_0_103_689 ();
 sg13g2_fill_1 FILLER_0_103_691 ();
 sg13g2_fill_1 FILLER_0_103_733 ();
 sg13g2_decap_4 FILLER_0_103_760 ();
 sg13g2_fill_2 FILLER_0_103_814 ();
 sg13g2_fill_2 FILLER_0_103_838 ();
 sg13g2_fill_1 FILLER_0_103_840 ();
 sg13g2_fill_2 FILLER_0_103_866 ();
 sg13g2_decap_8 FILLER_0_103_872 ();
 sg13g2_decap_8 FILLER_0_103_883 ();
 sg13g2_fill_2 FILLER_0_103_890 ();
 sg13g2_fill_2 FILLER_0_103_897 ();
 sg13g2_fill_1 FILLER_0_103_899 ();
 sg13g2_decap_8 FILLER_0_103_926 ();
 sg13g2_decap_8 FILLER_0_103_933 ();
 sg13g2_decap_8 FILLER_0_103_940 ();
 sg13g2_decap_8 FILLER_0_103_947 ();
 sg13g2_fill_2 FILLER_0_103_954 ();
 sg13g2_decap_8 FILLER_0_103_973 ();
 sg13g2_decap_8 FILLER_0_103_980 ();
 sg13g2_decap_8 FILLER_0_103_987 ();
 sg13g2_decap_4 FILLER_0_103_994 ();
 sg13g2_fill_2 FILLER_0_103_1002 ();
 sg13g2_decap_4 FILLER_0_103_1009 ();
 sg13g2_fill_2 FILLER_0_103_1023 ();
 sg13g2_decap_8 FILLER_0_103_1045 ();
 sg13g2_decap_8 FILLER_0_103_1052 ();
 sg13g2_decap_8 FILLER_0_103_1059 ();
 sg13g2_decap_8 FILLER_0_103_1066 ();
 sg13g2_decap_8 FILLER_0_103_1073 ();
 sg13g2_decap_8 FILLER_0_103_1080 ();
 sg13g2_decap_8 FILLER_0_103_1087 ();
 sg13g2_decap_8 FILLER_0_103_1094 ();
 sg13g2_decap_8 FILLER_0_103_1101 ();
 sg13g2_decap_8 FILLER_0_103_1108 ();
 sg13g2_decap_8 FILLER_0_103_1115 ();
 sg13g2_decap_8 FILLER_0_103_1122 ();
 sg13g2_decap_8 FILLER_0_103_1129 ();
 sg13g2_decap_8 FILLER_0_103_1136 ();
 sg13g2_decap_8 FILLER_0_103_1143 ();
 sg13g2_decap_8 FILLER_0_103_1150 ();
 sg13g2_decap_8 FILLER_0_103_1157 ();
 sg13g2_decap_8 FILLER_0_103_1164 ();
 sg13g2_decap_8 FILLER_0_103_1171 ();
 sg13g2_decap_8 FILLER_0_103_1178 ();
 sg13g2_decap_8 FILLER_0_103_1185 ();
 sg13g2_decap_8 FILLER_0_103_1192 ();
 sg13g2_decap_8 FILLER_0_103_1199 ();
 sg13g2_decap_8 FILLER_0_103_1206 ();
 sg13g2_decap_8 FILLER_0_103_1213 ();
 sg13g2_decap_8 FILLER_0_103_1220 ();
 sg13g2_fill_1 FILLER_0_103_1227 ();
 sg13g2_decap_8 FILLER_0_104_0 ();
 sg13g2_decap_8 FILLER_0_104_7 ();
 sg13g2_decap_8 FILLER_0_104_14 ();
 sg13g2_decap_8 FILLER_0_104_21 ();
 sg13g2_decap_8 FILLER_0_104_28 ();
 sg13g2_decap_8 FILLER_0_104_35 ();
 sg13g2_decap_8 FILLER_0_104_42 ();
 sg13g2_decap_8 FILLER_0_104_49 ();
 sg13g2_fill_1 FILLER_0_104_56 ();
 sg13g2_fill_2 FILLER_0_104_98 ();
 sg13g2_fill_1 FILLER_0_104_100 ();
 sg13g2_decap_8 FILLER_0_104_127 ();
 sg13g2_decap_8 FILLER_0_104_134 ();
 sg13g2_decap_8 FILLER_0_104_141 ();
 sg13g2_decap_8 FILLER_0_104_148 ();
 sg13g2_fill_2 FILLER_0_104_155 ();
 sg13g2_decap_8 FILLER_0_104_167 ();
 sg13g2_fill_2 FILLER_0_104_174 ();
 sg13g2_decap_8 FILLER_0_104_202 ();
 sg13g2_decap_8 FILLER_0_104_209 ();
 sg13g2_fill_2 FILLER_0_104_216 ();
 sg13g2_fill_1 FILLER_0_104_218 ();
 sg13g2_fill_1 FILLER_0_104_223 ();
 sg13g2_fill_2 FILLER_0_104_228 ();
 sg13g2_fill_1 FILLER_0_104_256 ();
 sg13g2_fill_2 FILLER_0_104_283 ();
 sg13g2_fill_1 FILLER_0_104_311 ();
 sg13g2_decap_8 FILLER_0_104_342 ();
 sg13g2_decap_8 FILLER_0_104_349 ();
 sg13g2_fill_1 FILLER_0_104_356 ();
 sg13g2_decap_8 FILLER_0_104_372 ();
 sg13g2_fill_1 FILLER_0_104_379 ();
 sg13g2_fill_2 FILLER_0_104_384 ();
 sg13g2_decap_4 FILLER_0_104_412 ();
 sg13g2_fill_1 FILLER_0_104_416 ();
 sg13g2_fill_1 FILLER_0_104_457 ();
 sg13g2_decap_8 FILLER_0_104_492 ();
 sg13g2_decap_8 FILLER_0_104_499 ();
 sg13g2_decap_8 FILLER_0_104_506 ();
 sg13g2_decap_8 FILLER_0_104_513 ();
 sg13g2_decap_8 FILLER_0_104_520 ();
 sg13g2_decap_8 FILLER_0_104_527 ();
 sg13g2_decap_4 FILLER_0_104_534 ();
 sg13g2_fill_1 FILLER_0_104_538 ();
 sg13g2_decap_8 FILLER_0_104_543 ();
 sg13g2_decap_8 FILLER_0_104_550 ();
 sg13g2_decap_8 FILLER_0_104_557 ();
 sg13g2_decap_8 FILLER_0_104_564 ();
 sg13g2_decap_8 FILLER_0_104_571 ();
 sg13g2_decap_8 FILLER_0_104_578 ();
 sg13g2_decap_8 FILLER_0_104_585 ();
 sg13g2_decap_4 FILLER_0_104_592 ();
 sg13g2_fill_1 FILLER_0_104_596 ();
 sg13g2_decap_8 FILLER_0_104_602 ();
 sg13g2_fill_1 FILLER_0_104_609 ();
 sg13g2_decap_8 FILLER_0_104_620 ();
 sg13g2_decap_4 FILLER_0_104_627 ();
 sg13g2_fill_2 FILLER_0_104_631 ();
 sg13g2_decap_4 FILLER_0_104_643 ();
 sg13g2_fill_2 FILLER_0_104_647 ();
 sg13g2_fill_2 FILLER_0_104_690 ();
 sg13g2_fill_1 FILLER_0_104_692 ();
 sg13g2_fill_2 FILLER_0_104_697 ();
 sg13g2_fill_1 FILLER_0_104_699 ();
 sg13g2_fill_2 FILLER_0_104_710 ();
 sg13g2_fill_1 FILLER_0_104_712 ();
 sg13g2_fill_1 FILLER_0_104_717 ();
 sg13g2_fill_2 FILLER_0_104_728 ();
 sg13g2_fill_1 FILLER_0_104_730 ();
 sg13g2_fill_1 FILLER_0_104_746 ();
 sg13g2_decap_8 FILLER_0_104_762 ();
 sg13g2_decap_4 FILLER_0_104_783 ();
 sg13g2_decap_8 FILLER_0_104_797 ();
 sg13g2_decap_8 FILLER_0_104_830 ();
 sg13g2_fill_1 FILLER_0_104_837 ();
 sg13g2_fill_1 FILLER_0_104_842 ();
 sg13g2_decap_8 FILLER_0_104_853 ();
 sg13g2_fill_1 FILLER_0_104_860 ();
 sg13g2_fill_2 FILLER_0_104_897 ();
 sg13g2_fill_1 FILLER_0_104_899 ();
 sg13g2_fill_2 FILLER_0_104_913 ();
 sg13g2_fill_1 FILLER_0_104_915 ();
 sg13g2_decap_4 FILLER_0_104_942 ();
 sg13g2_decap_8 FILLER_0_104_980 ();
 sg13g2_decap_4 FILLER_0_104_987 ();
 sg13g2_fill_1 FILLER_0_104_991 ();
 sg13g2_decap_8 FILLER_0_104_996 ();
 sg13g2_decap_8 FILLER_0_104_1003 ();
 sg13g2_decap_8 FILLER_0_104_1010 ();
 sg13g2_decap_8 FILLER_0_104_1017 ();
 sg13g2_decap_8 FILLER_0_104_1024 ();
 sg13g2_decap_8 FILLER_0_104_1031 ();
 sg13g2_decap_8 FILLER_0_104_1038 ();
 sg13g2_decap_8 FILLER_0_104_1045 ();
 sg13g2_decap_8 FILLER_0_104_1052 ();
 sg13g2_decap_8 FILLER_0_104_1059 ();
 sg13g2_decap_8 FILLER_0_104_1066 ();
 sg13g2_decap_8 FILLER_0_104_1073 ();
 sg13g2_decap_8 FILLER_0_104_1080 ();
 sg13g2_decap_8 FILLER_0_104_1087 ();
 sg13g2_decap_8 FILLER_0_104_1094 ();
 sg13g2_decap_8 FILLER_0_104_1101 ();
 sg13g2_decap_8 FILLER_0_104_1108 ();
 sg13g2_decap_8 FILLER_0_104_1115 ();
 sg13g2_decap_8 FILLER_0_104_1122 ();
 sg13g2_decap_8 FILLER_0_104_1129 ();
 sg13g2_decap_8 FILLER_0_104_1136 ();
 sg13g2_decap_8 FILLER_0_104_1143 ();
 sg13g2_decap_8 FILLER_0_104_1150 ();
 sg13g2_decap_8 FILLER_0_104_1157 ();
 sg13g2_decap_8 FILLER_0_104_1164 ();
 sg13g2_decap_8 FILLER_0_104_1171 ();
 sg13g2_decap_8 FILLER_0_104_1178 ();
 sg13g2_decap_8 FILLER_0_104_1185 ();
 sg13g2_decap_8 FILLER_0_104_1192 ();
 sg13g2_decap_8 FILLER_0_104_1199 ();
 sg13g2_decap_8 FILLER_0_104_1206 ();
 sg13g2_decap_8 FILLER_0_104_1213 ();
 sg13g2_decap_8 FILLER_0_104_1220 ();
 sg13g2_fill_1 FILLER_0_104_1227 ();
 sg13g2_decap_8 FILLER_0_105_0 ();
 sg13g2_decap_8 FILLER_0_105_7 ();
 sg13g2_decap_8 FILLER_0_105_14 ();
 sg13g2_decap_8 FILLER_0_105_21 ();
 sg13g2_decap_8 FILLER_0_105_28 ();
 sg13g2_decap_8 FILLER_0_105_35 ();
 sg13g2_decap_4 FILLER_0_105_42 ();
 sg13g2_decap_8 FILLER_0_105_91 ();
 sg13g2_fill_1 FILLER_0_105_117 ();
 sg13g2_fill_1 FILLER_0_105_128 ();
 sg13g2_fill_1 FILLER_0_105_147 ();
 sg13g2_fill_2 FILLER_0_105_153 ();
 sg13g2_fill_1 FILLER_0_105_190 ();
 sg13g2_decap_4 FILLER_0_105_195 ();
 sg13g2_decap_8 FILLER_0_105_209 ();
 sg13g2_decap_8 FILLER_0_105_216 ();
 sg13g2_decap_4 FILLER_0_105_223 ();
 sg13g2_fill_1 FILLER_0_105_227 ();
 sg13g2_fill_1 FILLER_0_105_238 ();
 sg13g2_fill_2 FILLER_0_105_249 ();
 sg13g2_fill_2 FILLER_0_105_261 ();
 sg13g2_fill_2 FILLER_0_105_273 ();
 sg13g2_decap_8 FILLER_0_105_279 ();
 sg13g2_decap_8 FILLER_0_105_286 ();
 sg13g2_decap_8 FILLER_0_105_293 ();
 sg13g2_decap_8 FILLER_0_105_300 ();
 sg13g2_fill_2 FILLER_0_105_307 ();
 sg13g2_decap_4 FILLER_0_105_317 ();
 sg13g2_fill_1 FILLER_0_105_321 ();
 sg13g2_decap_8 FILLER_0_105_337 ();
 sg13g2_decap_8 FILLER_0_105_378 ();
 sg13g2_decap_8 FILLER_0_105_385 ();
 sg13g2_fill_2 FILLER_0_105_392 ();
 sg13g2_decap_8 FILLER_0_105_398 ();
 sg13g2_decap_8 FILLER_0_105_405 ();
 sg13g2_decap_8 FILLER_0_105_412 ();
 sg13g2_fill_2 FILLER_0_105_419 ();
 sg13g2_decap_8 FILLER_0_105_452 ();
 sg13g2_fill_1 FILLER_0_105_459 ();
 sg13g2_decap_4 FILLER_0_105_464 ();
 sg13g2_fill_2 FILLER_0_105_473 ();
 sg13g2_fill_2 FILLER_0_105_485 ();
 sg13g2_decap_4 FILLER_0_105_513 ();
 sg13g2_decap_4 FILLER_0_105_522 ();
 sg13g2_decap_4 FILLER_0_105_536 ();
 sg13g2_fill_1 FILLER_0_105_647 ();
 sg13g2_fill_2 FILLER_0_105_666 ();
 sg13g2_fill_1 FILLER_0_105_668 ();
 sg13g2_decap_4 FILLER_0_105_677 ();
 sg13g2_fill_1 FILLER_0_105_681 ();
 sg13g2_decap_8 FILLER_0_105_713 ();
 sg13g2_decap_8 FILLER_0_105_720 ();
 sg13g2_decap_8 FILLER_0_105_727 ();
 sg13g2_decap_8 FILLER_0_105_734 ();
 sg13g2_decap_8 FILLER_0_105_741 ();
 sg13g2_decap_8 FILLER_0_105_748 ();
 sg13g2_decap_4 FILLER_0_105_755 ();
 sg13g2_fill_2 FILLER_0_105_759 ();
 sg13g2_decap_8 FILLER_0_105_771 ();
 sg13g2_decap_8 FILLER_0_105_778 ();
 sg13g2_fill_1 FILLER_0_105_785 ();
 sg13g2_fill_1 FILLER_0_105_796 ();
 sg13g2_fill_2 FILLER_0_105_802 ();
 sg13g2_fill_2 FILLER_0_105_830 ();
 sg13g2_decap_4 FILLER_0_105_873 ();
 sg13g2_fill_2 FILLER_0_105_877 ();
 sg13g2_fill_2 FILLER_0_105_915 ();
 sg13g2_fill_1 FILLER_0_105_927 ();
 sg13g2_fill_1 FILLER_0_105_954 ();
 sg13g2_fill_1 FILLER_0_105_986 ();
 sg13g2_decap_8 FILLER_0_105_1027 ();
 sg13g2_decap_8 FILLER_0_105_1034 ();
 sg13g2_decap_8 FILLER_0_105_1041 ();
 sg13g2_decap_8 FILLER_0_105_1048 ();
 sg13g2_decap_8 FILLER_0_105_1055 ();
 sg13g2_decap_8 FILLER_0_105_1062 ();
 sg13g2_decap_8 FILLER_0_105_1069 ();
 sg13g2_decap_8 FILLER_0_105_1076 ();
 sg13g2_decap_8 FILLER_0_105_1083 ();
 sg13g2_decap_8 FILLER_0_105_1090 ();
 sg13g2_decap_8 FILLER_0_105_1097 ();
 sg13g2_decap_8 FILLER_0_105_1104 ();
 sg13g2_decap_8 FILLER_0_105_1111 ();
 sg13g2_decap_8 FILLER_0_105_1118 ();
 sg13g2_decap_8 FILLER_0_105_1125 ();
 sg13g2_decap_8 FILLER_0_105_1132 ();
 sg13g2_decap_8 FILLER_0_105_1139 ();
 sg13g2_decap_8 FILLER_0_105_1146 ();
 sg13g2_decap_8 FILLER_0_105_1153 ();
 sg13g2_decap_8 FILLER_0_105_1160 ();
 sg13g2_decap_8 FILLER_0_105_1167 ();
 sg13g2_decap_8 FILLER_0_105_1174 ();
 sg13g2_decap_8 FILLER_0_105_1181 ();
 sg13g2_decap_8 FILLER_0_105_1188 ();
 sg13g2_decap_8 FILLER_0_105_1195 ();
 sg13g2_decap_8 FILLER_0_105_1202 ();
 sg13g2_decap_8 FILLER_0_105_1209 ();
 sg13g2_decap_8 FILLER_0_105_1216 ();
 sg13g2_decap_4 FILLER_0_105_1223 ();
 sg13g2_fill_1 FILLER_0_105_1227 ();
 sg13g2_decap_8 FILLER_0_106_0 ();
 sg13g2_decap_8 FILLER_0_106_7 ();
 sg13g2_decap_8 FILLER_0_106_14 ();
 sg13g2_decap_8 FILLER_0_106_21 ();
 sg13g2_decap_8 FILLER_0_106_28 ();
 sg13g2_fill_2 FILLER_0_106_35 ();
 sg13g2_fill_1 FILLER_0_106_37 ();
 sg13g2_decap_4 FILLER_0_106_68 ();
 sg13g2_decap_8 FILLER_0_106_82 ();
 sg13g2_fill_2 FILLER_0_106_89 ();
 sg13g2_fill_1 FILLER_0_106_91 ();
 sg13g2_fill_2 FILLER_0_106_106 ();
 sg13g2_decap_4 FILLER_0_106_156 ();
 sg13g2_decap_8 FILLER_0_106_164 ();
 sg13g2_decap_4 FILLER_0_106_171 ();
 sg13g2_fill_1 FILLER_0_106_175 ();
 sg13g2_fill_1 FILLER_0_106_184 ();
 sg13g2_decap_8 FILLER_0_106_211 ();
 sg13g2_decap_8 FILLER_0_106_218 ();
 sg13g2_decap_8 FILLER_0_106_225 ();
 sg13g2_decap_8 FILLER_0_106_232 ();
 sg13g2_decap_8 FILLER_0_106_243 ();
 sg13g2_decap_8 FILLER_0_106_250 ();
 sg13g2_decap_4 FILLER_0_106_257 ();
 sg13g2_fill_1 FILLER_0_106_261 ();
 sg13g2_decap_8 FILLER_0_106_266 ();
 sg13g2_decap_8 FILLER_0_106_273 ();
 sg13g2_fill_2 FILLER_0_106_280 ();
 sg13g2_fill_1 FILLER_0_106_282 ();
 sg13g2_fill_2 FILLER_0_106_292 ();
 sg13g2_fill_1 FILLER_0_106_294 ();
 sg13g2_fill_2 FILLER_0_106_348 ();
 sg13g2_fill_1 FILLER_0_106_350 ();
 sg13g2_decap_8 FILLER_0_106_388 ();
 sg13g2_decap_8 FILLER_0_106_395 ();
 sg13g2_decap_8 FILLER_0_106_402 ();
 sg13g2_decap_8 FILLER_0_106_409 ();
 sg13g2_decap_8 FILLER_0_106_416 ();
 sg13g2_fill_2 FILLER_0_106_423 ();
 sg13g2_fill_1 FILLER_0_106_425 ();
 sg13g2_fill_1 FILLER_0_106_453 ();
 sg13g2_fill_1 FILLER_0_106_480 ();
 sg13g2_fill_1 FILLER_0_106_491 ();
 sg13g2_fill_1 FILLER_0_106_497 ();
 sg13g2_fill_1 FILLER_0_106_503 ();
 sg13g2_fill_1 FILLER_0_106_530 ();
 sg13g2_fill_1 FILLER_0_106_597 ();
 sg13g2_fill_1 FILLER_0_106_628 ();
 sg13g2_fill_1 FILLER_0_106_634 ();
 sg13g2_fill_2 FILLER_0_106_639 ();
 sg13g2_fill_1 FILLER_0_106_641 ();
 sg13g2_decap_4 FILLER_0_106_668 ();
 sg13g2_fill_1 FILLER_0_106_676 ();
 sg13g2_fill_2 FILLER_0_106_703 ();
 sg13g2_fill_1 FILLER_0_106_705 ();
 sg13g2_decap_4 FILLER_0_106_711 ();
 sg13g2_decap_4 FILLER_0_106_745 ();
 sg13g2_fill_1 FILLER_0_106_749 ();
 sg13g2_fill_2 FILLER_0_106_760 ();
 sg13g2_fill_2 FILLER_0_106_828 ();
 sg13g2_fill_1 FILLER_0_106_830 ();
 sg13g2_fill_2 FILLER_0_106_836 ();
 sg13g2_fill_1 FILLER_0_106_838 ();
 sg13g2_fill_2 FILLER_0_106_843 ();
 sg13g2_fill_1 FILLER_0_106_845 ();
 sg13g2_fill_2 FILLER_0_106_885 ();
 sg13g2_decap_4 FILLER_0_106_891 ();
 sg13g2_fill_2 FILLER_0_106_905 ();
 sg13g2_fill_1 FILLER_0_106_907 ();
 sg13g2_fill_2 FILLER_0_106_912 ();
 sg13g2_fill_1 FILLER_0_106_919 ();
 sg13g2_fill_1 FILLER_0_106_930 ();
 sg13g2_fill_1 FILLER_0_106_936 ();
 sg13g2_fill_2 FILLER_0_106_941 ();
 sg13g2_fill_2 FILLER_0_106_948 ();
 sg13g2_fill_2 FILLER_0_106_974 ();
 sg13g2_decap_4 FILLER_0_106_1002 ();
 sg13g2_decap_8 FILLER_0_106_1032 ();
 sg13g2_decap_8 FILLER_0_106_1039 ();
 sg13g2_decap_8 FILLER_0_106_1046 ();
 sg13g2_decap_8 FILLER_0_106_1053 ();
 sg13g2_decap_8 FILLER_0_106_1060 ();
 sg13g2_decap_8 FILLER_0_106_1067 ();
 sg13g2_decap_8 FILLER_0_106_1074 ();
 sg13g2_decap_8 FILLER_0_106_1081 ();
 sg13g2_decap_8 FILLER_0_106_1088 ();
 sg13g2_decap_8 FILLER_0_106_1095 ();
 sg13g2_decap_8 FILLER_0_106_1102 ();
 sg13g2_decap_8 FILLER_0_106_1109 ();
 sg13g2_decap_8 FILLER_0_106_1116 ();
 sg13g2_decap_8 FILLER_0_106_1123 ();
 sg13g2_decap_8 FILLER_0_106_1130 ();
 sg13g2_decap_8 FILLER_0_106_1137 ();
 sg13g2_decap_8 FILLER_0_106_1144 ();
 sg13g2_decap_8 FILLER_0_106_1151 ();
 sg13g2_decap_8 FILLER_0_106_1158 ();
 sg13g2_decap_8 FILLER_0_106_1165 ();
 sg13g2_decap_8 FILLER_0_106_1172 ();
 sg13g2_decap_8 FILLER_0_106_1179 ();
 sg13g2_decap_8 FILLER_0_106_1186 ();
 sg13g2_decap_8 FILLER_0_106_1193 ();
 sg13g2_decap_8 FILLER_0_106_1200 ();
 sg13g2_decap_8 FILLER_0_106_1207 ();
 sg13g2_decap_8 FILLER_0_106_1214 ();
 sg13g2_decap_8 FILLER_0_106_1221 ();
 sg13g2_decap_8 FILLER_0_107_0 ();
 sg13g2_decap_8 FILLER_0_107_7 ();
 sg13g2_decap_8 FILLER_0_107_14 ();
 sg13g2_decap_8 FILLER_0_107_21 ();
 sg13g2_decap_8 FILLER_0_107_28 ();
 sg13g2_decap_4 FILLER_0_107_35 ();
 sg13g2_fill_1 FILLER_0_107_39 ();
 sg13g2_fill_2 FILLER_0_107_45 ();
 sg13g2_fill_1 FILLER_0_107_47 ();
 sg13g2_fill_1 FILLER_0_107_57 ();
 sg13g2_decap_4 FILLER_0_107_72 ();
 sg13g2_fill_1 FILLER_0_107_76 ();
 sg13g2_fill_2 FILLER_0_107_85 ();
 sg13g2_fill_1 FILLER_0_107_87 ();
 sg13g2_decap_4 FILLER_0_107_122 ();
 sg13g2_fill_1 FILLER_0_107_126 ();
 sg13g2_decap_4 FILLER_0_107_158 ();
 sg13g2_fill_2 FILLER_0_107_171 ();
 sg13g2_decap_8 FILLER_0_107_217 ();
 sg13g2_decap_8 FILLER_0_107_224 ();
 sg13g2_decap_8 FILLER_0_107_231 ();
 sg13g2_decap_8 FILLER_0_107_238 ();
 sg13g2_decap_4 FILLER_0_107_245 ();
 sg13g2_decap_4 FILLER_0_107_280 ();
 sg13g2_fill_1 FILLER_0_107_284 ();
 sg13g2_fill_2 FILLER_0_107_311 ();
 sg13g2_fill_2 FILLER_0_107_318 ();
 sg13g2_fill_2 FILLER_0_107_324 ();
 sg13g2_fill_1 FILLER_0_107_326 ();
 sg13g2_fill_1 FILLER_0_107_337 ();
 sg13g2_fill_2 FILLER_0_107_348 ();
 sg13g2_fill_1 FILLER_0_107_350 ();
 sg13g2_decap_8 FILLER_0_107_386 ();
 sg13g2_decap_8 FILLER_0_107_393 ();
 sg13g2_decap_8 FILLER_0_107_400 ();
 sg13g2_decap_8 FILLER_0_107_407 ();
 sg13g2_decap_8 FILLER_0_107_414 ();
 sg13g2_decap_8 FILLER_0_107_421 ();
 sg13g2_fill_1 FILLER_0_107_428 ();
 sg13g2_fill_2 FILLER_0_107_455 ();
 sg13g2_fill_2 FILLER_0_107_490 ();
 sg13g2_fill_1 FILLER_0_107_492 ();
 sg13g2_fill_2 FILLER_0_107_497 ();
 sg13g2_fill_2 FILLER_0_107_537 ();
 sg13g2_decap_4 FILLER_0_107_553 ();
 sg13g2_fill_2 FILLER_0_107_583 ();
 sg13g2_fill_1 FILLER_0_107_585 ();
 sg13g2_fill_2 FILLER_0_107_596 ();
 sg13g2_decap_4 FILLER_0_107_608 ();
 sg13g2_fill_1 FILLER_0_107_612 ();
 sg13g2_decap_8 FILLER_0_107_618 ();
 sg13g2_decap_4 FILLER_0_107_625 ();
 sg13g2_fill_1 FILLER_0_107_629 ();
 sg13g2_decap_8 FILLER_0_107_661 ();
 sg13g2_decap_4 FILLER_0_107_668 ();
 sg13g2_decap_4 FILLER_0_107_677 ();
 sg13g2_decap_8 FILLER_0_107_699 ();
 sg13g2_fill_1 FILLER_0_107_706 ();
 sg13g2_decap_4 FILLER_0_107_711 ();
 sg13g2_fill_1 FILLER_0_107_715 ();
 sg13g2_decap_8 FILLER_0_107_782 ();
 sg13g2_decap_4 FILLER_0_107_799 ();
 sg13g2_fill_1 FILLER_0_107_803 ();
 sg13g2_decap_4 FILLER_0_107_808 ();
 sg13g2_fill_1 FILLER_0_107_812 ();
 sg13g2_decap_8 FILLER_0_107_817 ();
 sg13g2_decap_8 FILLER_0_107_824 ();
 sg13g2_fill_2 FILLER_0_107_831 ();
 sg13g2_fill_1 FILLER_0_107_833 ();
 sg13g2_decap_8 FILLER_0_107_842 ();
 sg13g2_fill_2 FILLER_0_107_849 ();
 sg13g2_fill_1 FILLER_0_107_851 ();
 sg13g2_decap_4 FILLER_0_107_856 ();
 sg13g2_fill_1 FILLER_0_107_860 ();
 sg13g2_decap_8 FILLER_0_107_866 ();
 sg13g2_decap_4 FILLER_0_107_873 ();
 sg13g2_fill_1 FILLER_0_107_877 ();
 sg13g2_fill_1 FILLER_0_107_881 ();
 sg13g2_decap_8 FILLER_0_107_890 ();
 sg13g2_fill_2 FILLER_0_107_897 ();
 sg13g2_fill_1 FILLER_0_107_899 ();
 sg13g2_decap_4 FILLER_0_107_905 ();
 sg13g2_fill_1 FILLER_0_107_909 ();
 sg13g2_decap_4 FILLER_0_107_914 ();
 sg13g2_fill_2 FILLER_0_107_922 ();
 sg13g2_fill_2 FILLER_0_107_928 ();
 sg13g2_fill_1 FILLER_0_107_930 ();
 sg13g2_decap_8 FILLER_0_107_935 ();
 sg13g2_decap_8 FILLER_0_107_942 ();
 sg13g2_fill_2 FILLER_0_107_949 ();
 sg13g2_decap_8 FILLER_0_107_955 ();
 sg13g2_decap_8 FILLER_0_107_962 ();
 sg13g2_decap_4 FILLER_0_107_969 ();
 sg13g2_fill_1 FILLER_0_107_973 ();
 sg13g2_fill_1 FILLER_0_107_979 ();
 sg13g2_fill_1 FILLER_0_107_990 ();
 sg13g2_fill_1 FILLER_0_107_996 ();
 sg13g2_fill_1 FILLER_0_107_1007 ();
 sg13g2_decap_8 FILLER_0_107_1051 ();
 sg13g2_decap_8 FILLER_0_107_1058 ();
 sg13g2_decap_8 FILLER_0_107_1065 ();
 sg13g2_decap_8 FILLER_0_107_1072 ();
 sg13g2_decap_8 FILLER_0_107_1079 ();
 sg13g2_decap_8 FILLER_0_107_1086 ();
 sg13g2_decap_8 FILLER_0_107_1093 ();
 sg13g2_decap_8 FILLER_0_107_1100 ();
 sg13g2_decap_8 FILLER_0_107_1107 ();
 sg13g2_decap_8 FILLER_0_107_1114 ();
 sg13g2_decap_8 FILLER_0_107_1121 ();
 sg13g2_decap_8 FILLER_0_107_1128 ();
 sg13g2_decap_8 FILLER_0_107_1135 ();
 sg13g2_decap_8 FILLER_0_107_1142 ();
 sg13g2_decap_8 FILLER_0_107_1149 ();
 sg13g2_decap_8 FILLER_0_107_1156 ();
 sg13g2_decap_8 FILLER_0_107_1163 ();
 sg13g2_decap_8 FILLER_0_107_1170 ();
 sg13g2_decap_8 FILLER_0_107_1177 ();
 sg13g2_decap_8 FILLER_0_107_1184 ();
 sg13g2_decap_8 FILLER_0_107_1191 ();
 sg13g2_decap_8 FILLER_0_107_1198 ();
 sg13g2_decap_8 FILLER_0_107_1205 ();
 sg13g2_decap_8 FILLER_0_107_1212 ();
 sg13g2_decap_8 FILLER_0_107_1219 ();
 sg13g2_fill_2 FILLER_0_107_1226 ();
 sg13g2_decap_8 FILLER_0_108_0 ();
 sg13g2_decap_8 FILLER_0_108_7 ();
 sg13g2_decap_8 FILLER_0_108_14 ();
 sg13g2_decap_8 FILLER_0_108_21 ();
 sg13g2_decap_8 FILLER_0_108_28 ();
 sg13g2_decap_8 FILLER_0_108_35 ();
 sg13g2_decap_8 FILLER_0_108_42 ();
 sg13g2_fill_1 FILLER_0_108_106 ();
 sg13g2_fill_1 FILLER_0_108_117 ();
 sg13g2_fill_2 FILLER_0_108_123 ();
 sg13g2_fill_2 FILLER_0_108_151 ();
 sg13g2_decap_8 FILLER_0_108_192 ();
 sg13g2_decap_8 FILLER_0_108_199 ();
 sg13g2_decap_8 FILLER_0_108_206 ();
 sg13g2_decap_4 FILLER_0_108_213 ();
 sg13g2_decap_8 FILLER_0_108_222 ();
 sg13g2_decap_8 FILLER_0_108_229 ();
 sg13g2_fill_2 FILLER_0_108_236 ();
 sg13g2_fill_1 FILLER_0_108_238 ();
 sg13g2_decap_8 FILLER_0_108_244 ();
 sg13g2_decap_4 FILLER_0_108_251 ();
 sg13g2_fill_1 FILLER_0_108_255 ();
 sg13g2_decap_4 FILLER_0_108_276 ();
 sg13g2_fill_1 FILLER_0_108_280 ();
 sg13g2_fill_2 FILLER_0_108_296 ();
 sg13g2_decap_4 FILLER_0_108_324 ();
 sg13g2_fill_2 FILLER_0_108_333 ();
 sg13g2_fill_2 FILLER_0_108_365 ();
 sg13g2_fill_1 FILLER_0_108_367 ();
 sg13g2_decap_4 FILLER_0_108_372 ();
 sg13g2_fill_2 FILLER_0_108_390 ();
 sg13g2_decap_8 FILLER_0_108_397 ();
 sg13g2_decap_8 FILLER_0_108_404 ();
 sg13g2_fill_1 FILLER_0_108_411 ();
 sg13g2_fill_1 FILLER_0_108_422 ();
 sg13g2_fill_1 FILLER_0_108_449 ();
 sg13g2_fill_1 FILLER_0_108_455 ();
 sg13g2_fill_1 FILLER_0_108_460 ();
 sg13g2_decap_8 FILLER_0_108_487 ();
 sg13g2_fill_2 FILLER_0_108_494 ();
 sg13g2_fill_1 FILLER_0_108_496 ();
 sg13g2_decap_8 FILLER_0_108_539 ();
 sg13g2_decap_8 FILLER_0_108_546 ();
 sg13g2_decap_8 FILLER_0_108_553 ();
 sg13g2_fill_2 FILLER_0_108_560 ();
 sg13g2_fill_1 FILLER_0_108_575 ();
 sg13g2_decap_4 FILLER_0_108_586 ();
 sg13g2_fill_2 FILLER_0_108_590 ();
 sg13g2_decap_4 FILLER_0_108_609 ();
 sg13g2_decap_4 FILLER_0_108_654 ();
 sg13g2_fill_1 FILLER_0_108_658 ();
 sg13g2_fill_2 FILLER_0_108_689 ();
 sg13g2_fill_1 FILLER_0_108_731 ();
 sg13g2_decap_8 FILLER_0_108_742 ();
 sg13g2_fill_1 FILLER_0_108_758 ();
 sg13g2_fill_2 FILLER_0_108_763 ();
 sg13g2_decap_8 FILLER_0_108_769 ();
 sg13g2_fill_1 FILLER_0_108_776 ();
 sg13g2_fill_2 FILLER_0_108_784 ();
 sg13g2_fill_1 FILLER_0_108_789 ();
 sg13g2_decap_8 FILLER_0_108_794 ();
 sg13g2_fill_2 FILLER_0_108_801 ();
 sg13g2_fill_2 FILLER_0_108_811 ();
 sg13g2_fill_2 FILLER_0_108_817 ();
 sg13g2_fill_1 FILLER_0_108_819 ();
 sg13g2_fill_1 FILLER_0_108_824 ();
 sg13g2_decap_8 FILLER_0_108_830 ();
 sg13g2_fill_2 FILLER_0_108_841 ();
 sg13g2_decap_4 FILLER_0_108_869 ();
 sg13g2_fill_1 FILLER_0_108_881 ();
 sg13g2_fill_1 FILLER_0_108_891 ();
 sg13g2_fill_2 FILLER_0_108_901 ();
 sg13g2_fill_1 FILLER_0_108_929 ();
 sg13g2_decap_8 FILLER_0_108_964 ();
 sg13g2_decap_8 FILLER_0_108_971 ();
 sg13g2_decap_8 FILLER_0_108_978 ();
 sg13g2_decap_8 FILLER_0_108_985 ();
 sg13g2_fill_2 FILLER_0_108_992 ();
 sg13g2_fill_1 FILLER_0_108_994 ();
 sg13g2_decap_8 FILLER_0_108_999 ();
 sg13g2_decap_8 FILLER_0_108_1006 ();
 sg13g2_fill_1 FILLER_0_108_1013 ();
 sg13g2_decap_8 FILLER_0_108_1059 ();
 sg13g2_decap_8 FILLER_0_108_1066 ();
 sg13g2_decap_8 FILLER_0_108_1073 ();
 sg13g2_decap_8 FILLER_0_108_1080 ();
 sg13g2_decap_8 FILLER_0_108_1087 ();
 sg13g2_decap_8 FILLER_0_108_1094 ();
 sg13g2_decap_8 FILLER_0_108_1101 ();
 sg13g2_decap_8 FILLER_0_108_1108 ();
 sg13g2_decap_8 FILLER_0_108_1115 ();
 sg13g2_decap_8 FILLER_0_108_1122 ();
 sg13g2_decap_8 FILLER_0_108_1129 ();
 sg13g2_decap_8 FILLER_0_108_1136 ();
 sg13g2_decap_8 FILLER_0_108_1143 ();
 sg13g2_decap_8 FILLER_0_108_1150 ();
 sg13g2_decap_8 FILLER_0_108_1157 ();
 sg13g2_decap_8 FILLER_0_108_1164 ();
 sg13g2_decap_8 FILLER_0_108_1171 ();
 sg13g2_decap_8 FILLER_0_108_1178 ();
 sg13g2_decap_8 FILLER_0_108_1185 ();
 sg13g2_decap_8 FILLER_0_108_1192 ();
 sg13g2_decap_8 FILLER_0_108_1199 ();
 sg13g2_decap_8 FILLER_0_108_1206 ();
 sg13g2_decap_8 FILLER_0_108_1213 ();
 sg13g2_decap_8 FILLER_0_108_1220 ();
 sg13g2_fill_1 FILLER_0_108_1227 ();
 sg13g2_decap_8 FILLER_0_109_0 ();
 sg13g2_decap_8 FILLER_0_109_7 ();
 sg13g2_decap_8 FILLER_0_109_14 ();
 sg13g2_decap_8 FILLER_0_109_21 ();
 sg13g2_decap_8 FILLER_0_109_28 ();
 sg13g2_decap_4 FILLER_0_109_35 ();
 sg13g2_fill_2 FILLER_0_109_80 ();
 sg13g2_fill_1 FILLER_0_109_82 ();
 sg13g2_decap_8 FILLER_0_109_109 ();
 sg13g2_decap_4 FILLER_0_109_116 ();
 sg13g2_decap_4 FILLER_0_109_125 ();
 sg13g2_fill_1 FILLER_0_109_129 ();
 sg13g2_fill_1 FILLER_0_109_142 ();
 sg13g2_decap_4 FILLER_0_109_153 ();
 sg13g2_fill_1 FILLER_0_109_161 ();
 sg13g2_decap_4 FILLER_0_109_172 ();
 sg13g2_fill_1 FILLER_0_109_201 ();
 sg13g2_decap_8 FILLER_0_109_210 ();
 sg13g2_decap_8 FILLER_0_109_217 ();
 sg13g2_decap_8 FILLER_0_109_224 ();
 sg13g2_decap_8 FILLER_0_109_231 ();
 sg13g2_decap_4 FILLER_0_109_238 ();
 sg13g2_decap_4 FILLER_0_109_268 ();
 sg13g2_fill_2 FILLER_0_109_276 ();
 sg13g2_decap_8 FILLER_0_109_308 ();
 sg13g2_decap_4 FILLER_0_109_315 ();
 sg13g2_fill_1 FILLER_0_109_319 ();
 sg13g2_fill_2 FILLER_0_109_346 ();
 sg13g2_decap_4 FILLER_0_109_359 ();
 sg13g2_fill_1 FILLER_0_109_363 ();
 sg13g2_fill_2 FILLER_0_109_421 ();
 sg13g2_decap_8 FILLER_0_109_449 ();
 sg13g2_decap_4 FILLER_0_109_456 ();
 sg13g2_fill_2 FILLER_0_109_460 ();
 sg13g2_fill_1 FILLER_0_109_466 ();
 sg13g2_decap_4 FILLER_0_109_492 ();
 sg13g2_fill_2 FILLER_0_109_496 ();
 sg13g2_decap_8 FILLER_0_109_531 ();
 sg13g2_decap_8 FILLER_0_109_538 ();
 sg13g2_decap_8 FILLER_0_109_545 ();
 sg13g2_decap_8 FILLER_0_109_578 ();
 sg13g2_decap_8 FILLER_0_109_585 ();
 sg13g2_fill_1 FILLER_0_109_600 ();
 sg13g2_decap_4 FILLER_0_109_632 ();
 sg13g2_fill_1 FILLER_0_109_636 ();
 sg13g2_fill_2 FILLER_0_109_641 ();
 sg13g2_fill_2 FILLER_0_109_654 ();
 sg13g2_fill_2 FILLER_0_109_669 ();
 sg13g2_fill_1 FILLER_0_109_671 ();
 sg13g2_decap_8 FILLER_0_109_698 ();
 sg13g2_fill_2 FILLER_0_109_731 ();
 sg13g2_decap_8 FILLER_0_109_746 ();
 sg13g2_decap_4 FILLER_0_109_753 ();
 sg13g2_fill_2 FILLER_0_109_757 ();
 sg13g2_fill_2 FILLER_0_109_768 ();
 sg13g2_fill_1 FILLER_0_109_776 ();
 sg13g2_fill_1 FILLER_0_109_861 ();
 sg13g2_fill_2 FILLER_0_109_887 ();
 sg13g2_fill_1 FILLER_0_109_889 ();
 sg13g2_fill_1 FILLER_0_109_931 ();
 sg13g2_fill_1 FILLER_0_109_936 ();
 sg13g2_fill_2 FILLER_0_109_976 ();
 sg13g2_fill_1 FILLER_0_109_978 ();
 sg13g2_fill_1 FILLER_0_109_985 ();
 sg13g2_fill_1 FILLER_0_109_998 ();
 sg13g2_decap_8 FILLER_0_109_1012 ();
 sg13g2_decap_4 FILLER_0_109_1019 ();
 sg13g2_decap_8 FILLER_0_109_1052 ();
 sg13g2_decap_8 FILLER_0_109_1059 ();
 sg13g2_decap_8 FILLER_0_109_1066 ();
 sg13g2_decap_8 FILLER_0_109_1073 ();
 sg13g2_decap_8 FILLER_0_109_1080 ();
 sg13g2_decap_8 FILLER_0_109_1087 ();
 sg13g2_decap_8 FILLER_0_109_1094 ();
 sg13g2_decap_8 FILLER_0_109_1101 ();
 sg13g2_decap_8 FILLER_0_109_1108 ();
 sg13g2_decap_8 FILLER_0_109_1115 ();
 sg13g2_decap_8 FILLER_0_109_1122 ();
 sg13g2_decap_8 FILLER_0_109_1129 ();
 sg13g2_decap_8 FILLER_0_109_1136 ();
 sg13g2_decap_8 FILLER_0_109_1143 ();
 sg13g2_decap_8 FILLER_0_109_1150 ();
 sg13g2_decap_8 FILLER_0_109_1157 ();
 sg13g2_decap_8 FILLER_0_109_1164 ();
 sg13g2_decap_8 FILLER_0_109_1171 ();
 sg13g2_decap_8 FILLER_0_109_1178 ();
 sg13g2_decap_8 FILLER_0_109_1185 ();
 sg13g2_decap_8 FILLER_0_109_1192 ();
 sg13g2_decap_8 FILLER_0_109_1199 ();
 sg13g2_decap_8 FILLER_0_109_1206 ();
 sg13g2_decap_8 FILLER_0_109_1213 ();
 sg13g2_decap_8 FILLER_0_109_1220 ();
 sg13g2_fill_1 FILLER_0_109_1227 ();
 sg13g2_decap_8 FILLER_0_110_0 ();
 sg13g2_decap_8 FILLER_0_110_7 ();
 sg13g2_decap_8 FILLER_0_110_14 ();
 sg13g2_decap_8 FILLER_0_110_21 ();
 sg13g2_decap_8 FILLER_0_110_28 ();
 sg13g2_decap_8 FILLER_0_110_35 ();
 sg13g2_decap_4 FILLER_0_110_42 ();
 sg13g2_fill_1 FILLER_0_110_46 ();
 sg13g2_decap_8 FILLER_0_110_56 ();
 sg13g2_decap_4 FILLER_0_110_63 ();
 sg13g2_decap_8 FILLER_0_110_108 ();
 sg13g2_decap_8 FILLER_0_110_141 ();
 sg13g2_decap_4 FILLER_0_110_148 ();
 sg13g2_decap_4 FILLER_0_110_178 ();
 sg13g2_fill_1 FILLER_0_110_182 ();
 sg13g2_decap_8 FILLER_0_110_213 ();
 sg13g2_decap_8 FILLER_0_110_220 ();
 sg13g2_decap_8 FILLER_0_110_227 ();
 sg13g2_decap_8 FILLER_0_110_234 ();
 sg13g2_decap_8 FILLER_0_110_241 ();
 sg13g2_fill_1 FILLER_0_110_252 ();
 sg13g2_decap_8 FILLER_0_110_264 ();
 sg13g2_decap_8 FILLER_0_110_271 ();
 sg13g2_decap_8 FILLER_0_110_278 ();
 sg13g2_fill_2 FILLER_0_110_285 ();
 sg13g2_fill_1 FILLER_0_110_287 ();
 sg13g2_decap_8 FILLER_0_110_303 ();
 sg13g2_fill_2 FILLER_0_110_310 ();
 sg13g2_fill_1 FILLER_0_110_312 ();
 sg13g2_fill_2 FILLER_0_110_330 ();
 sg13g2_fill_1 FILLER_0_110_332 ();
 sg13g2_decap_8 FILLER_0_110_353 ();
 sg13g2_decap_4 FILLER_0_110_360 ();
 sg13g2_fill_2 FILLER_0_110_364 ();
 sg13g2_decap_8 FILLER_0_110_392 ();
 sg13g2_fill_2 FILLER_0_110_399 ();
 sg13g2_fill_1 FILLER_0_110_401 ();
 sg13g2_fill_1 FILLER_0_110_406 ();
 sg13g2_fill_1 FILLER_0_110_411 ();
 sg13g2_decap_4 FILLER_0_110_422 ();
 sg13g2_decap_8 FILLER_0_110_451 ();
 sg13g2_fill_2 FILLER_0_110_458 ();
 sg13g2_decap_4 FILLER_0_110_496 ();
 sg13g2_fill_2 FILLER_0_110_500 ();
 sg13g2_decap_8 FILLER_0_110_532 ();
 sg13g2_decap_8 FILLER_0_110_539 ();
 sg13g2_decap_4 FILLER_0_110_546 ();
 sg13g2_fill_1 FILLER_0_110_550 ();
 sg13g2_decap_8 FILLER_0_110_581 ();
 sg13g2_decap_4 FILLER_0_110_588 ();
 sg13g2_fill_1 FILLER_0_110_618 ();
 sg13g2_fill_1 FILLER_0_110_671 ();
 sg13g2_fill_2 FILLER_0_110_682 ();
 sg13g2_decap_8 FILLER_0_110_688 ();
 sg13g2_decap_8 FILLER_0_110_695 ();
 sg13g2_decap_8 FILLER_0_110_702 ();
 sg13g2_decap_4 FILLER_0_110_709 ();
 sg13g2_fill_2 FILLER_0_110_713 ();
 sg13g2_decap_4 FILLER_0_110_719 ();
 sg13g2_fill_2 FILLER_0_110_745 ();
 sg13g2_fill_2 FILLER_0_110_782 ();
 sg13g2_fill_1 FILLER_0_110_789 ();
 sg13g2_fill_1 FILLER_0_110_795 ();
 sg13g2_fill_2 FILLER_0_110_832 ();
 sg13g2_decap_8 FILLER_0_110_916 ();
 sg13g2_decap_4 FILLER_0_110_923 ();
 sg13g2_fill_2 FILLER_0_110_940 ();
 sg13g2_fill_1 FILLER_0_110_942 ();
 sg13g2_decap_8 FILLER_0_110_1015 ();
 sg13g2_decap_8 FILLER_0_110_1022 ();
 sg13g2_fill_2 FILLER_0_110_1029 ();
 sg13g2_decap_8 FILLER_0_110_1062 ();
 sg13g2_decap_8 FILLER_0_110_1069 ();
 sg13g2_decap_8 FILLER_0_110_1076 ();
 sg13g2_decap_8 FILLER_0_110_1083 ();
 sg13g2_decap_8 FILLER_0_110_1090 ();
 sg13g2_decap_8 FILLER_0_110_1097 ();
 sg13g2_decap_8 FILLER_0_110_1104 ();
 sg13g2_decap_8 FILLER_0_110_1111 ();
 sg13g2_decap_8 FILLER_0_110_1118 ();
 sg13g2_decap_8 FILLER_0_110_1125 ();
 sg13g2_decap_8 FILLER_0_110_1132 ();
 sg13g2_decap_8 FILLER_0_110_1139 ();
 sg13g2_decap_8 FILLER_0_110_1146 ();
 sg13g2_decap_8 FILLER_0_110_1153 ();
 sg13g2_decap_8 FILLER_0_110_1160 ();
 sg13g2_decap_8 FILLER_0_110_1167 ();
 sg13g2_decap_8 FILLER_0_110_1174 ();
 sg13g2_decap_8 FILLER_0_110_1181 ();
 sg13g2_decap_8 FILLER_0_110_1188 ();
 sg13g2_decap_8 FILLER_0_110_1195 ();
 sg13g2_decap_8 FILLER_0_110_1202 ();
 sg13g2_decap_8 FILLER_0_110_1209 ();
 sg13g2_decap_8 FILLER_0_110_1216 ();
 sg13g2_decap_4 FILLER_0_110_1223 ();
 sg13g2_fill_1 FILLER_0_110_1227 ();
 sg13g2_decap_8 FILLER_0_111_0 ();
 sg13g2_decap_8 FILLER_0_111_7 ();
 sg13g2_decap_8 FILLER_0_111_14 ();
 sg13g2_decap_8 FILLER_0_111_21 ();
 sg13g2_decap_8 FILLER_0_111_28 ();
 sg13g2_decap_8 FILLER_0_111_35 ();
 sg13g2_decap_4 FILLER_0_111_42 ();
 sg13g2_decap_8 FILLER_0_111_72 ();
 sg13g2_fill_2 FILLER_0_111_79 ();
 sg13g2_fill_1 FILLER_0_111_85 ();
 sg13g2_fill_1 FILLER_0_111_91 ();
 sg13g2_decap_8 FILLER_0_111_118 ();
 sg13g2_fill_2 FILLER_0_111_125 ();
 sg13g2_fill_2 FILLER_0_111_132 ();
 sg13g2_decap_4 FILLER_0_111_175 ();
 sg13g2_fill_1 FILLER_0_111_179 ();
 sg13g2_fill_2 FILLER_0_111_237 ();
 sg13g2_decap_8 FILLER_0_111_270 ();
 sg13g2_decap_8 FILLER_0_111_277 ();
 sg13g2_decap_4 FILLER_0_111_284 ();
 sg13g2_fill_1 FILLER_0_111_288 ();
 sg13g2_decap_8 FILLER_0_111_293 ();
 sg13g2_decap_8 FILLER_0_111_300 ();
 sg13g2_decap_8 FILLER_0_111_307 ();
 sg13g2_decap_8 FILLER_0_111_314 ();
 sg13g2_fill_2 FILLER_0_111_321 ();
 sg13g2_fill_2 FILLER_0_111_367 ();
 sg13g2_fill_2 FILLER_0_111_378 ();
 sg13g2_fill_2 FILLER_0_111_390 ();
 sg13g2_fill_1 FILLER_0_111_392 ();
 sg13g2_decap_8 FILLER_0_111_424 ();
 sg13g2_decap_4 FILLER_0_111_431 ();
 sg13g2_fill_1 FILLER_0_111_435 ();
 sg13g2_decap_8 FILLER_0_111_441 ();
 sg13g2_decap_8 FILLER_0_111_448 ();
 sg13g2_decap_4 FILLER_0_111_455 ();
 sg13g2_fill_2 FILLER_0_111_459 ();
 sg13g2_fill_2 FILLER_0_111_491 ();
 sg13g2_fill_1 FILLER_0_111_493 ();
 sg13g2_fill_2 FILLER_0_111_499 ();
 sg13g2_decap_4 FILLER_0_111_552 ();
 sg13g2_fill_1 FILLER_0_111_556 ();
 sg13g2_fill_1 FILLER_0_111_561 ();
 sg13g2_fill_2 FILLER_0_111_618 ();
 sg13g2_fill_1 FILLER_0_111_620 ();
 sg13g2_decap_8 FILLER_0_111_635 ();
 sg13g2_fill_1 FILLER_0_111_642 ();
 sg13g2_fill_2 FILLER_0_111_662 ();
 sg13g2_decap_4 FILLER_0_111_725 ();
 sg13g2_fill_1 FILLER_0_111_780 ();
 sg13g2_fill_1 FILLER_0_111_849 ();
 sg13g2_decap_8 FILLER_0_111_855 ();
 sg13g2_decap_8 FILLER_0_111_907 ();
 sg13g2_fill_1 FILLER_0_111_914 ();
 sg13g2_fill_2 FILLER_0_111_951 ();
 sg13g2_fill_2 FILLER_0_111_957 ();
 sg13g2_fill_1 FILLER_0_111_985 ();
 sg13g2_fill_1 FILLER_0_111_994 ();
 sg13g2_fill_1 FILLER_0_111_999 ();
 sg13g2_fill_1 FILLER_0_111_1009 ();
 sg13g2_decap_4 FILLER_0_111_1035 ();
 sg13g2_fill_1 FILLER_0_111_1039 ();
 sg13g2_decap_8 FILLER_0_111_1049 ();
 sg13g2_decap_8 FILLER_0_111_1056 ();
 sg13g2_decap_8 FILLER_0_111_1063 ();
 sg13g2_decap_8 FILLER_0_111_1070 ();
 sg13g2_decap_8 FILLER_0_111_1077 ();
 sg13g2_decap_8 FILLER_0_111_1084 ();
 sg13g2_decap_8 FILLER_0_111_1091 ();
 sg13g2_decap_8 FILLER_0_111_1098 ();
 sg13g2_decap_8 FILLER_0_111_1105 ();
 sg13g2_decap_8 FILLER_0_111_1112 ();
 sg13g2_decap_8 FILLER_0_111_1119 ();
 sg13g2_decap_8 FILLER_0_111_1126 ();
 sg13g2_decap_8 FILLER_0_111_1133 ();
 sg13g2_decap_8 FILLER_0_111_1140 ();
 sg13g2_decap_8 FILLER_0_111_1147 ();
 sg13g2_decap_8 FILLER_0_111_1154 ();
 sg13g2_decap_8 FILLER_0_111_1161 ();
 sg13g2_decap_8 FILLER_0_111_1168 ();
 sg13g2_decap_8 FILLER_0_111_1175 ();
 sg13g2_decap_8 FILLER_0_111_1182 ();
 sg13g2_decap_8 FILLER_0_111_1189 ();
 sg13g2_decap_8 FILLER_0_111_1196 ();
 sg13g2_decap_8 FILLER_0_111_1203 ();
 sg13g2_decap_8 FILLER_0_111_1210 ();
 sg13g2_decap_8 FILLER_0_111_1217 ();
 sg13g2_decap_4 FILLER_0_111_1224 ();
 sg13g2_decap_8 FILLER_0_112_0 ();
 sg13g2_decap_8 FILLER_0_112_7 ();
 sg13g2_decap_8 FILLER_0_112_14 ();
 sg13g2_decap_8 FILLER_0_112_21 ();
 sg13g2_decap_8 FILLER_0_112_28 ();
 sg13g2_decap_8 FILLER_0_112_35 ();
 sg13g2_decap_8 FILLER_0_112_42 ();
 sg13g2_fill_2 FILLER_0_112_49 ();
 sg13g2_decap_4 FILLER_0_112_64 ();
 sg13g2_fill_2 FILLER_0_112_68 ();
 sg13g2_decap_8 FILLER_0_112_80 ();
 sg13g2_decap_4 FILLER_0_112_87 ();
 sg13g2_fill_1 FILLER_0_112_91 ();
 sg13g2_fill_1 FILLER_0_112_116 ();
 sg13g2_fill_2 FILLER_0_112_150 ();
 sg13g2_decap_8 FILLER_0_112_182 ();
 sg13g2_decap_4 FILLER_0_112_189 ();
 sg13g2_decap_8 FILLER_0_112_197 ();
 sg13g2_decap_8 FILLER_0_112_204 ();
 sg13g2_decap_4 FILLER_0_112_211 ();
 sg13g2_fill_2 FILLER_0_112_215 ();
 sg13g2_decap_4 FILLER_0_112_248 ();
 sg13g2_decap_8 FILLER_0_112_313 ();
 sg13g2_decap_4 FILLER_0_112_320 ();
 sg13g2_fill_2 FILLER_0_112_324 ();
 sg13g2_decap_8 FILLER_0_112_356 ();
 sg13g2_fill_2 FILLER_0_112_363 ();
 sg13g2_fill_2 FILLER_0_112_401 ();
 sg13g2_fill_1 FILLER_0_112_403 ();
 sg13g2_decap_4 FILLER_0_112_409 ();
 sg13g2_fill_1 FILLER_0_112_413 ();
 sg13g2_fill_2 FILLER_0_112_424 ();
 sg13g2_fill_1 FILLER_0_112_426 ();
 sg13g2_decap_8 FILLER_0_112_432 ();
 sg13g2_decap_8 FILLER_0_112_439 ();
 sg13g2_decap_8 FILLER_0_112_446 ();
 sg13g2_decap_8 FILLER_0_112_453 ();
 sg13g2_decap_8 FILLER_0_112_460 ();
 sg13g2_fill_2 FILLER_0_112_467 ();
 sg13g2_fill_1 FILLER_0_112_469 ();
 sg13g2_decap_8 FILLER_0_112_501 ();
 sg13g2_decap_8 FILLER_0_112_508 ();
 sg13g2_fill_2 FILLER_0_112_515 ();
 sg13g2_fill_1 FILLER_0_112_517 ();
 sg13g2_fill_1 FILLER_0_112_533 ();
 sg13g2_fill_2 FILLER_0_112_565 ();
 sg13g2_fill_2 FILLER_0_112_577 ();
 sg13g2_fill_2 FILLER_0_112_589 ();
 sg13g2_fill_1 FILLER_0_112_591 ();
 sg13g2_fill_1 FILLER_0_112_596 ();
 sg13g2_fill_2 FILLER_0_112_605 ();
 sg13g2_fill_1 FILLER_0_112_607 ();
 sg13g2_decap_8 FILLER_0_112_623 ();
 sg13g2_decap_8 FILLER_0_112_630 ();
 sg13g2_decap_8 FILLER_0_112_637 ();
 sg13g2_decap_8 FILLER_0_112_644 ();
 sg13g2_decap_4 FILLER_0_112_666 ();
 sg13g2_fill_2 FILLER_0_112_674 ();
 sg13g2_fill_1 FILLER_0_112_676 ();
 sg13g2_fill_2 FILLER_0_112_726 ();
 sg13g2_fill_1 FILLER_0_112_728 ();
 sg13g2_fill_2 FILLER_0_112_747 ();
 sg13g2_fill_1 FILLER_0_112_771 ();
 sg13g2_fill_1 FILLER_0_112_775 ();
 sg13g2_fill_2 FILLER_0_112_798 ();
 sg13g2_decap_8 FILLER_0_112_804 ();
 sg13g2_decap_8 FILLER_0_112_815 ();
 sg13g2_decap_8 FILLER_0_112_822 ();
 sg13g2_fill_2 FILLER_0_112_864 ();
 sg13g2_decap_4 FILLER_0_112_896 ();
 sg13g2_fill_1 FILLER_0_112_900 ();
 sg13g2_decap_8 FILLER_0_112_911 ();
 sg13g2_decap_4 FILLER_0_112_918 ();
 sg13g2_decap_4 FILLER_0_112_926 ();
 sg13g2_fill_1 FILLER_0_112_930 ();
 sg13g2_fill_1 FILLER_0_112_939 ();
 sg13g2_fill_2 FILLER_0_112_945 ();
 sg13g2_decap_8 FILLER_0_112_956 ();
 sg13g2_fill_2 FILLER_0_112_963 ();
 sg13g2_fill_1 FILLER_0_112_965 ();
 sg13g2_fill_1 FILLER_0_112_1011 ();
 sg13g2_fill_2 FILLER_0_112_1044 ();
 sg13g2_decap_8 FILLER_0_112_1056 ();
 sg13g2_decap_8 FILLER_0_112_1063 ();
 sg13g2_decap_8 FILLER_0_112_1070 ();
 sg13g2_decap_8 FILLER_0_112_1077 ();
 sg13g2_decap_8 FILLER_0_112_1084 ();
 sg13g2_decap_8 FILLER_0_112_1091 ();
 sg13g2_decap_8 FILLER_0_112_1098 ();
 sg13g2_decap_8 FILLER_0_112_1105 ();
 sg13g2_decap_8 FILLER_0_112_1112 ();
 sg13g2_decap_8 FILLER_0_112_1119 ();
 sg13g2_decap_8 FILLER_0_112_1126 ();
 sg13g2_decap_8 FILLER_0_112_1133 ();
 sg13g2_decap_8 FILLER_0_112_1140 ();
 sg13g2_decap_8 FILLER_0_112_1147 ();
 sg13g2_decap_8 FILLER_0_112_1154 ();
 sg13g2_decap_8 FILLER_0_112_1161 ();
 sg13g2_decap_8 FILLER_0_112_1168 ();
 sg13g2_decap_8 FILLER_0_112_1175 ();
 sg13g2_decap_8 FILLER_0_112_1182 ();
 sg13g2_decap_8 FILLER_0_112_1189 ();
 sg13g2_decap_8 FILLER_0_112_1196 ();
 sg13g2_decap_8 FILLER_0_112_1203 ();
 sg13g2_decap_8 FILLER_0_112_1210 ();
 sg13g2_decap_8 FILLER_0_112_1217 ();
 sg13g2_decap_4 FILLER_0_112_1224 ();
 sg13g2_decap_8 FILLER_0_113_0 ();
 sg13g2_decap_8 FILLER_0_113_7 ();
 sg13g2_decap_8 FILLER_0_113_14 ();
 sg13g2_decap_8 FILLER_0_113_21 ();
 sg13g2_decap_8 FILLER_0_113_28 ();
 sg13g2_decap_8 FILLER_0_113_35 ();
 sg13g2_decap_8 FILLER_0_113_42 ();
 sg13g2_fill_1 FILLER_0_113_49 ();
 sg13g2_decap_8 FILLER_0_113_80 ();
 sg13g2_decap_8 FILLER_0_113_87 ();
 sg13g2_decap_8 FILLER_0_113_94 ();
 sg13g2_decap_8 FILLER_0_113_101 ();
 sg13g2_decap_8 FILLER_0_113_108 ();
 sg13g2_decap_8 FILLER_0_113_115 ();
 sg13g2_decap_8 FILLER_0_113_122 ();
 sg13g2_decap_8 FILLER_0_113_129 ();
 sg13g2_decap_8 FILLER_0_113_136 ();
 sg13g2_decap_8 FILLER_0_113_143 ();
 sg13g2_decap_4 FILLER_0_113_150 ();
 sg13g2_decap_8 FILLER_0_113_179 ();
 sg13g2_decap_8 FILLER_0_113_186 ();
 sg13g2_decap_8 FILLER_0_113_193 ();
 sg13g2_decap_8 FILLER_0_113_200 ();
 sg13g2_decap_4 FILLER_0_113_212 ();
 sg13g2_fill_2 FILLER_0_113_216 ();
 sg13g2_fill_1 FILLER_0_113_222 ();
 sg13g2_fill_1 FILLER_0_113_233 ();
 sg13g2_fill_1 FILLER_0_113_238 ();
 sg13g2_fill_1 FILLER_0_113_244 ();
 sg13g2_fill_1 FILLER_0_113_255 ();
 sg13g2_decap_4 FILLER_0_113_327 ();
 sg13g2_fill_1 FILLER_0_113_331 ();
 sg13g2_decap_8 FILLER_0_113_342 ();
 sg13g2_decap_8 FILLER_0_113_349 ();
 sg13g2_decap_8 FILLER_0_113_360 ();
 sg13g2_fill_2 FILLER_0_113_367 ();
 sg13g2_fill_1 FILLER_0_113_369 ();
 sg13g2_decap_8 FILLER_0_113_374 ();
 sg13g2_decap_4 FILLER_0_113_381 ();
 sg13g2_decap_8 FILLER_0_113_390 ();
 sg13g2_decap_8 FILLER_0_113_397 ();
 sg13g2_fill_1 FILLER_0_113_404 ();
 sg13g2_decap_4 FILLER_0_113_457 ();
 sg13g2_fill_1 FILLER_0_113_461 ();
 sg13g2_fill_1 FILLER_0_113_491 ();
 sg13g2_decap_8 FILLER_0_113_496 ();
 sg13g2_decap_8 FILLER_0_113_503 ();
 sg13g2_decap_8 FILLER_0_113_510 ();
 sg13g2_decap_4 FILLER_0_113_517 ();
 sg13g2_fill_1 FILLER_0_113_521 ();
 sg13g2_fill_2 FILLER_0_113_548 ();
 sg13g2_decap_4 FILLER_0_113_560 ();
 sg13g2_fill_2 FILLER_0_113_564 ();
 sg13g2_decap_8 FILLER_0_113_622 ();
 sg13g2_decap_8 FILLER_0_113_629 ();
 sg13g2_decap_8 FILLER_0_113_666 ();
 sg13g2_decap_8 FILLER_0_113_673 ();
 sg13g2_decap_8 FILLER_0_113_680 ();
 sg13g2_fill_2 FILLER_0_113_687 ();
 sg13g2_decap_8 FILLER_0_113_708 ();
 sg13g2_fill_2 FILLER_0_113_756 ();
 sg13g2_fill_2 FILLER_0_113_773 ();
 sg13g2_decap_8 FILLER_0_113_806 ();
 sg13g2_decap_8 FILLER_0_113_813 ();
 sg13g2_decap_8 FILLER_0_113_820 ();
 sg13g2_decap_8 FILLER_0_113_827 ();
 sg13g2_fill_1 FILLER_0_113_839 ();
 sg13g2_fill_2 FILLER_0_113_871 ();
 sg13g2_fill_1 FILLER_0_113_882 ();
 sg13g2_fill_1 FILLER_0_113_886 ();
 sg13g2_fill_1 FILLER_0_113_945 ();
 sg13g2_fill_2 FILLER_0_113_950 ();
 sg13g2_decap_4 FILLER_0_113_956 ();
 sg13g2_decap_8 FILLER_0_113_970 ();
 sg13g2_fill_2 FILLER_0_113_977 ();
 sg13g2_fill_1 FILLER_0_113_986 ();
 sg13g2_fill_1 FILLER_0_113_997 ();
 sg13g2_fill_2 FILLER_0_113_1003 ();
 sg13g2_fill_2 FILLER_0_113_1035 ();
 sg13g2_decap_8 FILLER_0_113_1063 ();
 sg13g2_decap_8 FILLER_0_113_1070 ();
 sg13g2_decap_8 FILLER_0_113_1077 ();
 sg13g2_decap_8 FILLER_0_113_1084 ();
 sg13g2_decap_8 FILLER_0_113_1091 ();
 sg13g2_decap_8 FILLER_0_113_1098 ();
 sg13g2_decap_8 FILLER_0_113_1105 ();
 sg13g2_decap_8 FILLER_0_113_1112 ();
 sg13g2_decap_8 FILLER_0_113_1119 ();
 sg13g2_decap_8 FILLER_0_113_1126 ();
 sg13g2_decap_8 FILLER_0_113_1133 ();
 sg13g2_decap_8 FILLER_0_113_1140 ();
 sg13g2_decap_8 FILLER_0_113_1147 ();
 sg13g2_decap_8 FILLER_0_113_1154 ();
 sg13g2_decap_8 FILLER_0_113_1161 ();
 sg13g2_decap_8 FILLER_0_113_1168 ();
 sg13g2_decap_8 FILLER_0_113_1175 ();
 sg13g2_decap_8 FILLER_0_113_1182 ();
 sg13g2_decap_8 FILLER_0_113_1189 ();
 sg13g2_decap_8 FILLER_0_113_1196 ();
 sg13g2_decap_8 FILLER_0_113_1203 ();
 sg13g2_decap_8 FILLER_0_113_1210 ();
 sg13g2_decap_8 FILLER_0_113_1217 ();
 sg13g2_decap_4 FILLER_0_113_1224 ();
 sg13g2_decap_8 FILLER_0_114_0 ();
 sg13g2_decap_8 FILLER_0_114_7 ();
 sg13g2_decap_8 FILLER_0_114_14 ();
 sg13g2_decap_8 FILLER_0_114_21 ();
 sg13g2_decap_8 FILLER_0_114_28 ();
 sg13g2_decap_8 FILLER_0_114_35 ();
 sg13g2_decap_4 FILLER_0_114_42 ();
 sg13g2_decap_8 FILLER_0_114_87 ();
 sg13g2_decap_8 FILLER_0_114_94 ();
 sg13g2_decap_8 FILLER_0_114_101 ();
 sg13g2_decap_8 FILLER_0_114_108 ();
 sg13g2_decap_8 FILLER_0_114_115 ();
 sg13g2_decap_8 FILLER_0_114_122 ();
 sg13g2_decap_8 FILLER_0_114_129 ();
 sg13g2_decap_8 FILLER_0_114_136 ();
 sg13g2_decap_8 FILLER_0_114_143 ();
 sg13g2_fill_1 FILLER_0_114_150 ();
 sg13g2_decap_4 FILLER_0_114_190 ();
 sg13g2_fill_2 FILLER_0_114_199 ();
 sg13g2_fill_1 FILLER_0_114_201 ();
 sg13g2_fill_1 FILLER_0_114_211 ();
 sg13g2_decap_8 FILLER_0_114_232 ();
 sg13g2_decap_4 FILLER_0_114_239 ();
 sg13g2_decap_8 FILLER_0_114_247 ();
 sg13g2_decap_8 FILLER_0_114_254 ();
 sg13g2_fill_2 FILLER_0_114_295 ();
 sg13g2_fill_1 FILLER_0_114_307 ();
 sg13g2_fill_2 FILLER_0_114_334 ();
 sg13g2_fill_2 FILLER_0_114_346 ();
 sg13g2_fill_2 FILLER_0_114_379 ();
 sg13g2_fill_2 FILLER_0_114_407 ();
 sg13g2_fill_1 FILLER_0_114_409 ();
 sg13g2_fill_1 FILLER_0_114_414 ();
 sg13g2_fill_2 FILLER_0_114_425 ();
 sg13g2_fill_1 FILLER_0_114_427 ();
 sg13g2_decap_4 FILLER_0_114_433 ();
 sg13g2_fill_2 FILLER_0_114_441 ();
 sg13g2_decap_8 FILLER_0_114_486 ();
 sg13g2_decap_8 FILLER_0_114_493 ();
 sg13g2_decap_8 FILLER_0_114_500 ();
 sg13g2_decap_8 FILLER_0_114_507 ();
 sg13g2_decap_8 FILLER_0_114_514 ();
 sg13g2_decap_8 FILLER_0_114_521 ();
 sg13g2_decap_4 FILLER_0_114_528 ();
 sg13g2_fill_1 FILLER_0_114_532 ();
 sg13g2_decap_8 FILLER_0_114_559 ();
 sg13g2_decap_4 FILLER_0_114_566 ();
 sg13g2_fill_2 FILLER_0_114_570 ();
 sg13g2_decap_4 FILLER_0_114_576 ();
 sg13g2_fill_1 FILLER_0_114_599 ();
 sg13g2_fill_1 FILLER_0_114_626 ();
 sg13g2_decap_8 FILLER_0_114_637 ();
 sg13g2_fill_2 FILLER_0_114_644 ();
 sg13g2_fill_1 FILLER_0_114_646 ();
 sg13g2_decap_8 FILLER_0_114_665 ();
 sg13g2_fill_2 FILLER_0_114_672 ();
 sg13g2_decap_4 FILLER_0_114_704 ();
 sg13g2_fill_1 FILLER_0_114_739 ();
 sg13g2_fill_1 FILLER_0_114_772 ();
 sg13g2_fill_1 FILLER_0_114_782 ();
 sg13g2_fill_2 FILLER_0_114_788 ();
 sg13g2_fill_1 FILLER_0_114_790 ();
 sg13g2_decap_8 FILLER_0_114_817 ();
 sg13g2_decap_4 FILLER_0_114_824 ();
 sg13g2_fill_1 FILLER_0_114_838 ();
 sg13g2_fill_1 FILLER_0_114_849 ();
 sg13g2_decap_8 FILLER_0_114_896 ();
 sg13g2_fill_1 FILLER_0_114_908 ();
 sg13g2_decap_8 FILLER_0_114_913 ();
 sg13g2_fill_1 FILLER_0_114_920 ();
 sg13g2_fill_2 FILLER_0_114_960 ();
 sg13g2_fill_1 FILLER_0_114_962 ();
 sg13g2_fill_1 FILLER_0_114_982 ();
 sg13g2_fill_1 FILLER_0_114_1014 ();
 sg13g2_fill_2 FILLER_0_114_1020 ();
 sg13g2_decap_8 FILLER_0_114_1026 ();
 sg13g2_decap_8 FILLER_0_114_1033 ();
 sg13g2_decap_8 FILLER_0_114_1074 ();
 sg13g2_decap_8 FILLER_0_114_1081 ();
 sg13g2_decap_8 FILLER_0_114_1088 ();
 sg13g2_decap_8 FILLER_0_114_1095 ();
 sg13g2_decap_8 FILLER_0_114_1102 ();
 sg13g2_decap_8 FILLER_0_114_1109 ();
 sg13g2_decap_8 FILLER_0_114_1116 ();
 sg13g2_decap_8 FILLER_0_114_1123 ();
 sg13g2_decap_8 FILLER_0_114_1130 ();
 sg13g2_decap_8 FILLER_0_114_1137 ();
 sg13g2_decap_8 FILLER_0_114_1144 ();
 sg13g2_decap_8 FILLER_0_114_1151 ();
 sg13g2_decap_8 FILLER_0_114_1158 ();
 sg13g2_decap_8 FILLER_0_114_1165 ();
 sg13g2_decap_8 FILLER_0_114_1172 ();
 sg13g2_decap_8 FILLER_0_114_1179 ();
 sg13g2_decap_8 FILLER_0_114_1186 ();
 sg13g2_decap_8 FILLER_0_114_1193 ();
 sg13g2_decap_8 FILLER_0_114_1200 ();
 sg13g2_decap_8 FILLER_0_114_1207 ();
 sg13g2_decap_8 FILLER_0_114_1214 ();
 sg13g2_decap_8 FILLER_0_114_1221 ();
 sg13g2_decap_8 FILLER_0_115_0 ();
 sg13g2_decap_8 FILLER_0_115_7 ();
 sg13g2_decap_8 FILLER_0_115_14 ();
 sg13g2_decap_8 FILLER_0_115_21 ();
 sg13g2_decap_8 FILLER_0_115_28 ();
 sg13g2_decap_8 FILLER_0_115_35 ();
 sg13g2_fill_2 FILLER_0_115_42 ();
 sg13g2_fill_1 FILLER_0_115_53 ();
 sg13g2_decap_8 FILLER_0_115_84 ();
 sg13g2_decap_8 FILLER_0_115_91 ();
 sg13g2_decap_8 FILLER_0_115_98 ();
 sg13g2_decap_8 FILLER_0_115_105 ();
 sg13g2_decap_8 FILLER_0_115_112 ();
 sg13g2_decap_8 FILLER_0_115_119 ();
 sg13g2_decap_8 FILLER_0_115_126 ();
 sg13g2_decap_8 FILLER_0_115_133 ();
 sg13g2_decap_8 FILLER_0_115_140 ();
 sg13g2_decap_8 FILLER_0_115_147 ();
 sg13g2_decap_8 FILLER_0_115_154 ();
 sg13g2_decap_8 FILLER_0_115_187 ();
 sg13g2_fill_2 FILLER_0_115_194 ();
 sg13g2_fill_2 FILLER_0_115_200 ();
 sg13g2_fill_1 FILLER_0_115_202 ();
 sg13g2_decap_8 FILLER_0_115_229 ();
 sg13g2_decap_8 FILLER_0_115_236 ();
 sg13g2_decap_8 FILLER_0_115_243 ();
 sg13g2_decap_8 FILLER_0_115_250 ();
 sg13g2_decap_8 FILLER_0_115_257 ();
 sg13g2_decap_8 FILLER_0_115_264 ();
 sg13g2_decap_8 FILLER_0_115_271 ();
 sg13g2_decap_8 FILLER_0_115_278 ();
 sg13g2_fill_2 FILLER_0_115_285 ();
 sg13g2_fill_1 FILLER_0_115_298 ();
 sg13g2_decap_4 FILLER_0_115_303 ();
 sg13g2_fill_2 FILLER_0_115_307 ();
 sg13g2_fill_2 FILLER_0_115_319 ();
 sg13g2_fill_1 FILLER_0_115_325 ();
 sg13g2_fill_1 FILLER_0_115_336 ();
 sg13g2_fill_1 FILLER_0_115_347 ();
 sg13g2_decap_4 FILLER_0_115_374 ();
 sg13g2_decap_8 FILLER_0_115_418 ();
 sg13g2_fill_2 FILLER_0_115_425 ();
 sg13g2_decap_8 FILLER_0_115_453 ();
 sg13g2_fill_2 FILLER_0_115_508 ();
 sg13g2_fill_1 FILLER_0_115_510 ();
 sg13g2_decap_8 FILLER_0_115_556 ();
 sg13g2_decap_4 FILLER_0_115_563 ();
 sg13g2_fill_1 FILLER_0_115_603 ();
 sg13g2_fill_2 FILLER_0_115_614 ();
 sg13g2_fill_1 FILLER_0_115_642 ();
 sg13g2_fill_2 FILLER_0_115_669 ();
 sg13g2_fill_1 FILLER_0_115_676 ();
 sg13g2_decap_8 FILLER_0_115_702 ();
 sg13g2_fill_1 FILLER_0_115_709 ();
 sg13g2_fill_2 FILLER_0_115_736 ();
 sg13g2_fill_1 FILLER_0_115_743 ();
 sg13g2_fill_1 FILLER_0_115_753 ();
 sg13g2_fill_1 FILLER_0_115_759 ();
 sg13g2_fill_2 FILLER_0_115_764 ();
 sg13g2_fill_1 FILLER_0_115_770 ();
 sg13g2_fill_2 FILLER_0_115_811 ();
 sg13g2_fill_2 FILLER_0_115_817 ();
 sg13g2_fill_2 FILLER_0_115_852 ();
 sg13g2_fill_1 FILLER_0_115_854 ();
 sg13g2_decap_8 FILLER_0_115_863 ();
 sg13g2_decap_8 FILLER_0_115_870 ();
 sg13g2_fill_2 FILLER_0_115_877 ();
 sg13g2_fill_1 FILLER_0_115_879 ();
 sg13g2_fill_2 FILLER_0_115_903 ();
 sg13g2_fill_2 FILLER_0_115_917 ();
 sg13g2_fill_1 FILLER_0_115_919 ();
 sg13g2_decap_4 FILLER_0_115_930 ();
 sg13g2_decap_8 FILLER_0_115_943 ();
 sg13g2_fill_1 FILLER_0_115_950 ();
 sg13g2_fill_2 FILLER_0_115_955 ();
 sg13g2_fill_1 FILLER_0_115_957 ();
 sg13g2_fill_2 FILLER_0_115_975 ();
 sg13g2_decap_8 FILLER_0_115_1013 ();
 sg13g2_decap_8 FILLER_0_115_1020 ();
 sg13g2_decap_8 FILLER_0_115_1027 ();
 sg13g2_decap_8 FILLER_0_115_1034 ();
 sg13g2_fill_1 FILLER_0_115_1041 ();
 sg13g2_decap_8 FILLER_0_115_1080 ();
 sg13g2_decap_8 FILLER_0_115_1087 ();
 sg13g2_decap_8 FILLER_0_115_1094 ();
 sg13g2_decap_8 FILLER_0_115_1101 ();
 sg13g2_decap_8 FILLER_0_115_1108 ();
 sg13g2_decap_8 FILLER_0_115_1115 ();
 sg13g2_decap_8 FILLER_0_115_1122 ();
 sg13g2_decap_8 FILLER_0_115_1129 ();
 sg13g2_decap_8 FILLER_0_115_1136 ();
 sg13g2_decap_8 FILLER_0_115_1143 ();
 sg13g2_decap_8 FILLER_0_115_1150 ();
 sg13g2_decap_8 FILLER_0_115_1157 ();
 sg13g2_decap_8 FILLER_0_115_1164 ();
 sg13g2_decap_8 FILLER_0_115_1171 ();
 sg13g2_decap_8 FILLER_0_115_1178 ();
 sg13g2_decap_8 FILLER_0_115_1185 ();
 sg13g2_decap_8 FILLER_0_115_1192 ();
 sg13g2_decap_8 FILLER_0_115_1199 ();
 sg13g2_decap_8 FILLER_0_115_1206 ();
 sg13g2_decap_8 FILLER_0_115_1213 ();
 sg13g2_decap_8 FILLER_0_115_1220 ();
 sg13g2_fill_1 FILLER_0_115_1227 ();
 sg13g2_decap_8 FILLER_0_116_0 ();
 sg13g2_decap_8 FILLER_0_116_7 ();
 sg13g2_decap_8 FILLER_0_116_14 ();
 sg13g2_decap_8 FILLER_0_116_21 ();
 sg13g2_decap_8 FILLER_0_116_28 ();
 sg13g2_decap_4 FILLER_0_116_35 ();
 sg13g2_fill_1 FILLER_0_116_39 ();
 sg13g2_decap_8 FILLER_0_116_71 ();
 sg13g2_decap_8 FILLER_0_116_78 ();
 sg13g2_decap_8 FILLER_0_116_85 ();
 sg13g2_decap_8 FILLER_0_116_92 ();
 sg13g2_decap_8 FILLER_0_116_99 ();
 sg13g2_decap_8 FILLER_0_116_106 ();
 sg13g2_decap_8 FILLER_0_116_113 ();
 sg13g2_decap_8 FILLER_0_116_120 ();
 sg13g2_decap_8 FILLER_0_116_127 ();
 sg13g2_decap_4 FILLER_0_116_134 ();
 sg13g2_fill_1 FILLER_0_116_138 ();
 sg13g2_decap_8 FILLER_0_116_147 ();
 sg13g2_fill_2 FILLER_0_116_154 ();
 sg13g2_fill_1 FILLER_0_116_156 ();
 sg13g2_decap_8 FILLER_0_116_187 ();
 sg13g2_decap_8 FILLER_0_116_235 ();
 sg13g2_decap_8 FILLER_0_116_242 ();
 sg13g2_decap_8 FILLER_0_116_249 ();
 sg13g2_decap_8 FILLER_0_116_256 ();
 sg13g2_decap_8 FILLER_0_116_263 ();
 sg13g2_decap_8 FILLER_0_116_270 ();
 sg13g2_decap_8 FILLER_0_116_277 ();
 sg13g2_decap_8 FILLER_0_116_284 ();
 sg13g2_decap_8 FILLER_0_116_291 ();
 sg13g2_decap_8 FILLER_0_116_298 ();
 sg13g2_decap_4 FILLER_0_116_305 ();
 sg13g2_fill_2 FILLER_0_116_309 ();
 sg13g2_fill_1 FILLER_0_116_352 ();
 sg13g2_fill_2 FILLER_0_116_379 ();
 sg13g2_fill_2 FILLER_0_116_386 ();
 sg13g2_fill_1 FILLER_0_116_392 ();
 sg13g2_decap_8 FILLER_0_116_401 ();
 sg13g2_decap_8 FILLER_0_116_408 ();
 sg13g2_decap_8 FILLER_0_116_415 ();
 sg13g2_decap_8 FILLER_0_116_422 ();
 sg13g2_decap_4 FILLER_0_116_429 ();
 sg13g2_fill_2 FILLER_0_116_433 ();
 sg13g2_fill_2 FILLER_0_116_439 ();
 sg13g2_fill_1 FILLER_0_116_446 ();
 sg13g2_decap_8 FILLER_0_116_457 ();
 sg13g2_fill_1 FILLER_0_116_464 ();
 sg13g2_decap_4 FILLER_0_116_475 ();
 sg13g2_decap_8 FILLER_0_116_483 ();
 sg13g2_fill_2 FILLER_0_116_490 ();
 sg13g2_fill_1 FILLER_0_116_533 ();
 sg13g2_decap_8 FILLER_0_116_560 ();
 sg13g2_decap_4 FILLER_0_116_567 ();
 sg13g2_fill_2 FILLER_0_116_575 ();
 sg13g2_fill_1 FILLER_0_116_577 ();
 sg13g2_decap_8 FILLER_0_116_582 ();
 sg13g2_fill_1 FILLER_0_116_599 ();
 sg13g2_fill_1 FILLER_0_116_605 ();
 sg13g2_fill_1 FILLER_0_116_610 ();
 sg13g2_fill_1 FILLER_0_116_621 ();
 sg13g2_fill_2 FILLER_0_116_627 ();
 sg13g2_decap_8 FILLER_0_116_633 ();
 sg13g2_decap_8 FILLER_0_116_640 ();
 sg13g2_decap_4 FILLER_0_116_647 ();
 sg13g2_decap_8 FILLER_0_116_660 ();
 sg13g2_fill_2 FILLER_0_116_667 ();
 sg13g2_fill_1 FILLER_0_116_669 ();
 sg13g2_fill_2 FILLER_0_116_700 ();
 sg13g2_fill_1 FILLER_0_116_702 ();
 sg13g2_decap_8 FILLER_0_116_753 ();
 sg13g2_decap_8 FILLER_0_116_760 ();
 sg13g2_decap_8 FILLER_0_116_767 ();
 sg13g2_decap_8 FILLER_0_116_774 ();
 sg13g2_decap_8 FILLER_0_116_781 ();
 sg13g2_fill_1 FILLER_0_116_788 ();
 sg13g2_fill_2 FILLER_0_116_793 ();
 sg13g2_decap_4 FILLER_0_116_804 ();
 sg13g2_decap_4 FILLER_0_116_813 ();
 sg13g2_fill_2 FILLER_0_116_817 ();
 sg13g2_fill_2 FILLER_0_116_823 ();
 sg13g2_fill_1 FILLER_0_116_825 ();
 sg13g2_fill_2 FILLER_0_116_839 ();
 sg13g2_fill_1 FILLER_0_116_841 ();
 sg13g2_fill_2 FILLER_0_116_846 ();
 sg13g2_decap_8 FILLER_0_116_853 ();
 sg13g2_fill_2 FILLER_0_116_865 ();
 sg13g2_fill_1 FILLER_0_116_867 ();
 sg13g2_decap_4 FILLER_0_116_876 ();
 sg13g2_fill_1 FILLER_0_116_880 ();
 sg13g2_decap_4 FILLER_0_116_888 ();
 sg13g2_fill_1 FILLER_0_116_892 ();
 sg13g2_fill_1 FILLER_0_116_913 ();
 sg13g2_fill_2 FILLER_0_116_930 ();
 sg13g2_fill_1 FILLER_0_116_932 ();
 sg13g2_fill_1 FILLER_0_116_943 ();
 sg13g2_fill_2 FILLER_0_116_970 ();
 sg13g2_fill_2 FILLER_0_116_1007 ();
 sg13g2_fill_1 FILLER_0_116_1009 ();
 sg13g2_decap_4 FILLER_0_116_1015 ();
 sg13g2_fill_1 FILLER_0_116_1019 ();
 sg13g2_decap_4 FILLER_0_116_1024 ();
 sg13g2_fill_1 FILLER_0_116_1028 ();
 sg13g2_decap_8 FILLER_0_116_1037 ();
 sg13g2_fill_2 FILLER_0_116_1044 ();
 sg13g2_fill_1 FILLER_0_116_1046 ();
 sg13g2_decap_8 FILLER_0_116_1078 ();
 sg13g2_decap_8 FILLER_0_116_1085 ();
 sg13g2_decap_8 FILLER_0_116_1092 ();
 sg13g2_decap_8 FILLER_0_116_1099 ();
 sg13g2_decap_8 FILLER_0_116_1106 ();
 sg13g2_decap_8 FILLER_0_116_1113 ();
 sg13g2_decap_8 FILLER_0_116_1120 ();
 sg13g2_decap_8 FILLER_0_116_1127 ();
 sg13g2_decap_8 FILLER_0_116_1134 ();
 sg13g2_decap_8 FILLER_0_116_1141 ();
 sg13g2_decap_8 FILLER_0_116_1148 ();
 sg13g2_decap_8 FILLER_0_116_1155 ();
 sg13g2_decap_8 FILLER_0_116_1162 ();
 sg13g2_decap_8 FILLER_0_116_1169 ();
 sg13g2_decap_8 FILLER_0_116_1176 ();
 sg13g2_decap_8 FILLER_0_116_1183 ();
 sg13g2_decap_8 FILLER_0_116_1190 ();
 sg13g2_decap_8 FILLER_0_116_1197 ();
 sg13g2_decap_8 FILLER_0_116_1204 ();
 sg13g2_decap_8 FILLER_0_116_1211 ();
 sg13g2_decap_8 FILLER_0_116_1218 ();
 sg13g2_fill_2 FILLER_0_116_1225 ();
 sg13g2_fill_1 FILLER_0_116_1227 ();
 sg13g2_decap_8 FILLER_0_117_0 ();
 sg13g2_decap_8 FILLER_0_117_7 ();
 sg13g2_decap_8 FILLER_0_117_14 ();
 sg13g2_decap_8 FILLER_0_117_21 ();
 sg13g2_decap_8 FILLER_0_117_28 ();
 sg13g2_decap_4 FILLER_0_117_35 ();
 sg13g2_fill_1 FILLER_0_117_39 ();
 sg13g2_decap_8 FILLER_0_117_76 ();
 sg13g2_decap_8 FILLER_0_117_83 ();
 sg13g2_decap_8 FILLER_0_117_90 ();
 sg13g2_decap_8 FILLER_0_117_97 ();
 sg13g2_decap_8 FILLER_0_117_104 ();
 sg13g2_decap_8 FILLER_0_117_111 ();
 sg13g2_decap_8 FILLER_0_117_118 ();
 sg13g2_decap_8 FILLER_0_117_125 ();
 sg13g2_decap_8 FILLER_0_117_132 ();
 sg13g2_decap_8 FILLER_0_117_139 ();
 sg13g2_decap_8 FILLER_0_117_146 ();
 sg13g2_decap_4 FILLER_0_117_153 ();
 sg13g2_decap_8 FILLER_0_117_188 ();
 sg13g2_fill_2 FILLER_0_117_195 ();
 sg13g2_fill_1 FILLER_0_117_197 ();
 sg13g2_decap_8 FILLER_0_117_224 ();
 sg13g2_decap_8 FILLER_0_117_231 ();
 sg13g2_decap_8 FILLER_0_117_238 ();
 sg13g2_decap_8 FILLER_0_117_245 ();
 sg13g2_decap_8 FILLER_0_117_252 ();
 sg13g2_decap_8 FILLER_0_117_259 ();
 sg13g2_decap_8 FILLER_0_117_266 ();
 sg13g2_decap_8 FILLER_0_117_273 ();
 sg13g2_decap_8 FILLER_0_117_280 ();
 sg13g2_decap_8 FILLER_0_117_287 ();
 sg13g2_decap_8 FILLER_0_117_294 ();
 sg13g2_decap_8 FILLER_0_117_301 ();
 sg13g2_fill_2 FILLER_0_117_308 ();
 sg13g2_fill_1 FILLER_0_117_310 ();
 sg13g2_decap_8 FILLER_0_117_337 ();
 sg13g2_decap_4 FILLER_0_117_344 ();
 sg13g2_fill_1 FILLER_0_117_348 ();
 sg13g2_decap_8 FILLER_0_117_387 ();
 sg13g2_decap_8 FILLER_0_117_394 ();
 sg13g2_decap_8 FILLER_0_117_401 ();
 sg13g2_decap_8 FILLER_0_117_408 ();
 sg13g2_decap_8 FILLER_0_117_415 ();
 sg13g2_fill_1 FILLER_0_117_422 ();
 sg13g2_decap_8 FILLER_0_117_453 ();
 sg13g2_fill_2 FILLER_0_117_460 ();
 sg13g2_fill_1 FILLER_0_117_462 ();
 sg13g2_decap_8 FILLER_0_117_494 ();
 sg13g2_fill_1 FILLER_0_117_537 ();
 sg13g2_decap_8 FILLER_0_117_558 ();
 sg13g2_decap_4 FILLER_0_117_565 ();
 sg13g2_fill_1 FILLER_0_117_569 ();
 sg13g2_decap_8 FILLER_0_117_601 ();
 sg13g2_decap_8 FILLER_0_117_608 ();
 sg13g2_decap_8 FILLER_0_117_615 ();
 sg13g2_decap_8 FILLER_0_117_622 ();
 sg13g2_decap_8 FILLER_0_117_629 ();
 sg13g2_decap_8 FILLER_0_117_636 ();
 sg13g2_decap_8 FILLER_0_117_643 ();
 sg13g2_decap_8 FILLER_0_117_650 ();
 sg13g2_decap_4 FILLER_0_117_657 ();
 sg13g2_fill_1 FILLER_0_117_661 ();
 sg13g2_fill_2 FILLER_0_117_703 ();
 sg13g2_fill_2 FILLER_0_117_768 ();
 sg13g2_decap_8 FILLER_0_117_796 ();
 sg13g2_fill_1 FILLER_0_117_803 ();
 sg13g2_fill_1 FILLER_0_117_820 ();
 sg13g2_fill_1 FILLER_0_117_847 ();
 sg13g2_fill_2 FILLER_0_117_853 ();
 sg13g2_fill_1 FILLER_0_117_855 ();
 sg13g2_fill_1 FILLER_0_117_887 ();
 sg13g2_fill_2 FILLER_0_117_893 ();
 sg13g2_fill_1 FILLER_0_117_895 ();
 sg13g2_fill_1 FILLER_0_117_957 ();
 sg13g2_fill_2 FILLER_0_117_962 ();
 sg13g2_decap_8 FILLER_0_117_972 ();
 sg13g2_decap_4 FILLER_0_117_979 ();
 sg13g2_fill_2 FILLER_0_117_991 ();
 sg13g2_fill_1 FILLER_0_117_993 ();
 sg13g2_decap_8 FILLER_0_117_998 ();
 sg13g2_decap_8 FILLER_0_117_1005 ();
 sg13g2_fill_1 FILLER_0_117_1016 ();
 sg13g2_decap_4 FILLER_0_117_1037 ();
 sg13g2_fill_2 FILLER_0_117_1041 ();
 sg13g2_decap_8 FILLER_0_117_1074 ();
 sg13g2_decap_8 FILLER_0_117_1081 ();
 sg13g2_decap_8 FILLER_0_117_1088 ();
 sg13g2_decap_8 FILLER_0_117_1095 ();
 sg13g2_decap_8 FILLER_0_117_1102 ();
 sg13g2_decap_8 FILLER_0_117_1109 ();
 sg13g2_decap_8 FILLER_0_117_1116 ();
 sg13g2_decap_8 FILLER_0_117_1123 ();
 sg13g2_decap_8 FILLER_0_117_1130 ();
 sg13g2_decap_8 FILLER_0_117_1137 ();
 sg13g2_decap_8 FILLER_0_117_1144 ();
 sg13g2_decap_8 FILLER_0_117_1151 ();
 sg13g2_decap_8 FILLER_0_117_1158 ();
 sg13g2_decap_8 FILLER_0_117_1165 ();
 sg13g2_decap_8 FILLER_0_117_1172 ();
 sg13g2_decap_8 FILLER_0_117_1179 ();
 sg13g2_decap_8 FILLER_0_117_1186 ();
 sg13g2_decap_8 FILLER_0_117_1193 ();
 sg13g2_decap_8 FILLER_0_117_1200 ();
 sg13g2_decap_8 FILLER_0_117_1207 ();
 sg13g2_decap_8 FILLER_0_117_1214 ();
 sg13g2_decap_8 FILLER_0_117_1221 ();
 sg13g2_decap_8 FILLER_0_118_0 ();
 sg13g2_decap_8 FILLER_0_118_7 ();
 sg13g2_decap_8 FILLER_0_118_14 ();
 sg13g2_decap_8 FILLER_0_118_21 ();
 sg13g2_decap_8 FILLER_0_118_28 ();
 sg13g2_decap_8 FILLER_0_118_35 ();
 sg13g2_decap_4 FILLER_0_118_42 ();
 sg13g2_fill_1 FILLER_0_118_46 ();
 sg13g2_decap_4 FILLER_0_118_51 ();
 sg13g2_fill_2 FILLER_0_118_55 ();
 sg13g2_fill_2 FILLER_0_118_81 ();
 sg13g2_decap_8 FILLER_0_118_87 ();
 sg13g2_decap_8 FILLER_0_118_94 ();
 sg13g2_decap_8 FILLER_0_118_101 ();
 sg13g2_decap_8 FILLER_0_118_108 ();
 sg13g2_decap_8 FILLER_0_118_115 ();
 sg13g2_decap_8 FILLER_0_118_122 ();
 sg13g2_decap_8 FILLER_0_118_129 ();
 sg13g2_decap_8 FILLER_0_118_136 ();
 sg13g2_decap_8 FILLER_0_118_143 ();
 sg13g2_decap_8 FILLER_0_118_150 ();
 sg13g2_decap_8 FILLER_0_118_157 ();
 sg13g2_decap_4 FILLER_0_118_172 ();
 sg13g2_fill_2 FILLER_0_118_176 ();
 sg13g2_decap_8 FILLER_0_118_188 ();
 sg13g2_fill_1 FILLER_0_118_195 ();
 sg13g2_fill_2 FILLER_0_118_216 ();
 sg13g2_decap_8 FILLER_0_118_228 ();
 sg13g2_decap_8 FILLER_0_118_235 ();
 sg13g2_decap_8 FILLER_0_118_242 ();
 sg13g2_decap_8 FILLER_0_118_249 ();
 sg13g2_decap_8 FILLER_0_118_256 ();
 sg13g2_decap_8 FILLER_0_118_263 ();
 sg13g2_decap_8 FILLER_0_118_270 ();
 sg13g2_decap_8 FILLER_0_118_277 ();
 sg13g2_decap_8 FILLER_0_118_284 ();
 sg13g2_decap_8 FILLER_0_118_291 ();
 sg13g2_decap_8 FILLER_0_118_298 ();
 sg13g2_decap_8 FILLER_0_118_305 ();
 sg13g2_fill_1 FILLER_0_118_312 ();
 sg13g2_decap_4 FILLER_0_118_322 ();
 sg13g2_decap_8 FILLER_0_118_341 ();
 sg13g2_decap_8 FILLER_0_118_348 ();
 sg13g2_decap_8 FILLER_0_118_355 ();
 sg13g2_fill_2 FILLER_0_118_366 ();
 sg13g2_decap_8 FILLER_0_118_371 ();
 sg13g2_decap_8 FILLER_0_118_378 ();
 sg13g2_decap_8 FILLER_0_118_385 ();
 sg13g2_decap_8 FILLER_0_118_392 ();
 sg13g2_decap_8 FILLER_0_118_399 ();
 sg13g2_decap_8 FILLER_0_118_406 ();
 sg13g2_decap_8 FILLER_0_118_413 ();
 sg13g2_fill_2 FILLER_0_118_420 ();
 sg13g2_fill_2 FILLER_0_118_457 ();
 sg13g2_fill_1 FILLER_0_118_459 ();
 sg13g2_fill_2 FILLER_0_118_482 ();
 sg13g2_decap_8 FILLER_0_118_489 ();
 sg13g2_decap_8 FILLER_0_118_500 ();
 sg13g2_decap_8 FILLER_0_118_511 ();
 sg13g2_decap_8 FILLER_0_118_518 ();
 sg13g2_decap_8 FILLER_0_118_525 ();
 sg13g2_fill_2 FILLER_0_118_532 ();
 sg13g2_fill_1 FILLER_0_118_534 ();
 sg13g2_fill_2 FILLER_0_118_539 ();
 sg13g2_decap_8 FILLER_0_118_545 ();
 sg13g2_decap_8 FILLER_0_118_552 ();
 sg13g2_decap_8 FILLER_0_118_559 ();
 sg13g2_decap_8 FILLER_0_118_566 ();
 sg13g2_decap_8 FILLER_0_118_573 ();
 sg13g2_fill_1 FILLER_0_118_589 ();
 sg13g2_decap_8 FILLER_0_118_605 ();
 sg13g2_decap_8 FILLER_0_118_612 ();
 sg13g2_decap_8 FILLER_0_118_619 ();
 sg13g2_decap_8 FILLER_0_118_626 ();
 sg13g2_decap_8 FILLER_0_118_633 ();
 sg13g2_decap_8 FILLER_0_118_640 ();
 sg13g2_decap_8 FILLER_0_118_647 ();
 sg13g2_decap_8 FILLER_0_118_654 ();
 sg13g2_fill_2 FILLER_0_118_673 ();
 sg13g2_fill_1 FILLER_0_118_675 ();
 sg13g2_decap_8 FILLER_0_118_695 ();
 sg13g2_fill_1 FILLER_0_118_702 ();
 sg13g2_decap_4 FILLER_0_118_707 ();
 sg13g2_fill_1 FILLER_0_118_718 ();
 sg13g2_fill_1 FILLER_0_118_724 ();
 sg13g2_fill_1 FILLER_0_118_730 ();
 sg13g2_decap_4 FILLER_0_118_789 ();
 sg13g2_fill_2 FILLER_0_118_793 ();
 sg13g2_decap_4 FILLER_0_118_807 ();
 sg13g2_fill_2 FILLER_0_118_827 ();
 sg13g2_fill_2 FILLER_0_118_842 ();
 sg13g2_fill_2 FILLER_0_118_870 ();
 sg13g2_decap_4 FILLER_0_118_898 ();
 sg13g2_fill_1 FILLER_0_118_902 ();
 sg13g2_fill_1 FILLER_0_118_908 ();
 sg13g2_fill_2 FILLER_0_118_913 ();
 sg13g2_fill_1 FILLER_0_118_919 ();
 sg13g2_fill_1 FILLER_0_118_925 ();
 sg13g2_fill_1 FILLER_0_118_931 ();
 sg13g2_fill_1 FILLER_0_118_940 ();
 sg13g2_fill_2 FILLER_0_118_947 ();
 sg13g2_fill_1 FILLER_0_118_949 ();
 sg13g2_fill_2 FILLER_0_118_976 ();
 sg13g2_decap_8 FILLER_0_118_988 ();
 sg13g2_decap_8 FILLER_0_118_995 ();
 sg13g2_decap_8 FILLER_0_118_1002 ();
 sg13g2_fill_1 FILLER_0_118_1032 ();
 sg13g2_decap_4 FILLER_0_118_1051 ();
 sg13g2_fill_2 FILLER_0_118_1055 ();
 sg13g2_decap_8 FILLER_0_118_1083 ();
 sg13g2_decap_8 FILLER_0_118_1090 ();
 sg13g2_decap_8 FILLER_0_118_1097 ();
 sg13g2_decap_8 FILLER_0_118_1104 ();
 sg13g2_decap_8 FILLER_0_118_1111 ();
 sg13g2_decap_8 FILLER_0_118_1118 ();
 sg13g2_decap_8 FILLER_0_118_1125 ();
 sg13g2_decap_8 FILLER_0_118_1132 ();
 sg13g2_decap_8 FILLER_0_118_1139 ();
 sg13g2_decap_8 FILLER_0_118_1146 ();
 sg13g2_decap_8 FILLER_0_118_1153 ();
 sg13g2_decap_8 FILLER_0_118_1160 ();
 sg13g2_decap_8 FILLER_0_118_1167 ();
 sg13g2_decap_8 FILLER_0_118_1174 ();
 sg13g2_decap_8 FILLER_0_118_1181 ();
 sg13g2_decap_8 FILLER_0_118_1188 ();
 sg13g2_decap_8 FILLER_0_118_1195 ();
 sg13g2_decap_8 FILLER_0_118_1202 ();
 sg13g2_decap_8 FILLER_0_118_1209 ();
 sg13g2_decap_8 FILLER_0_118_1216 ();
 sg13g2_decap_4 FILLER_0_118_1223 ();
 sg13g2_fill_1 FILLER_0_118_1227 ();
 sg13g2_decap_8 FILLER_0_119_0 ();
 sg13g2_decap_8 FILLER_0_119_7 ();
 sg13g2_decap_8 FILLER_0_119_14 ();
 sg13g2_decap_8 FILLER_0_119_21 ();
 sg13g2_decap_8 FILLER_0_119_28 ();
 sg13g2_decap_4 FILLER_0_119_35 ();
 sg13g2_fill_2 FILLER_0_119_39 ();
 sg13g2_fill_1 FILLER_0_119_67 ();
 sg13g2_decap_8 FILLER_0_119_102 ();
 sg13g2_decap_8 FILLER_0_119_109 ();
 sg13g2_decap_8 FILLER_0_119_116 ();
 sg13g2_decap_8 FILLER_0_119_123 ();
 sg13g2_decap_8 FILLER_0_119_130 ();
 sg13g2_decap_8 FILLER_0_119_137 ();
 sg13g2_decap_8 FILLER_0_119_144 ();
 sg13g2_fill_1 FILLER_0_119_151 ();
 sg13g2_decap_8 FILLER_0_119_224 ();
 sg13g2_decap_8 FILLER_0_119_231 ();
 sg13g2_decap_8 FILLER_0_119_238 ();
 sg13g2_decap_8 FILLER_0_119_245 ();
 sg13g2_decap_8 FILLER_0_119_252 ();
 sg13g2_decap_8 FILLER_0_119_259 ();
 sg13g2_decap_8 FILLER_0_119_266 ();
 sg13g2_decap_8 FILLER_0_119_273 ();
 sg13g2_decap_8 FILLER_0_119_280 ();
 sg13g2_decap_8 FILLER_0_119_287 ();
 sg13g2_decap_8 FILLER_0_119_294 ();
 sg13g2_decap_4 FILLER_0_119_301 ();
 sg13g2_decap_8 FILLER_0_119_345 ();
 sg13g2_fill_1 FILLER_0_119_352 ();
 sg13g2_decap_8 FILLER_0_119_380 ();
 sg13g2_fill_2 FILLER_0_119_387 ();
 sg13g2_fill_1 FILLER_0_119_389 ();
 sg13g2_fill_2 FILLER_0_119_399 ();
 sg13g2_fill_1 FILLER_0_119_401 ();
 sg13g2_decap_8 FILLER_0_119_412 ();
 sg13g2_decap_8 FILLER_0_119_419 ();
 sg13g2_fill_2 FILLER_0_119_426 ();
 sg13g2_decap_8 FILLER_0_119_461 ();
 sg13g2_decap_4 FILLER_0_119_468 ();
 sg13g2_fill_1 FILLER_0_119_522 ();
 sg13g2_decap_8 FILLER_0_119_536 ();
 sg13g2_decap_8 FILLER_0_119_543 ();
 sg13g2_decap_8 FILLER_0_119_550 ();
 sg13g2_decap_8 FILLER_0_119_557 ();
 sg13g2_fill_2 FILLER_0_119_564 ();
 sg13g2_fill_2 FILLER_0_119_597 ();
 sg13g2_fill_2 FILLER_0_119_616 ();
 sg13g2_fill_2 FILLER_0_119_628 ();
 sg13g2_fill_1 FILLER_0_119_630 ();
 sg13g2_decap_8 FILLER_0_119_657 ();
 sg13g2_decap_4 FILLER_0_119_664 ();
 sg13g2_fill_2 FILLER_0_119_694 ();
 sg13g2_fill_2 FILLER_0_119_722 ();
 sg13g2_fill_2 FILLER_0_119_729 ();
 sg13g2_fill_2 FILLER_0_119_751 ();
 sg13g2_decap_8 FILLER_0_119_783 ();
 sg13g2_fill_1 FILLER_0_119_790 ();
 sg13g2_fill_2 FILLER_0_119_799 ();
 sg13g2_fill_1 FILLER_0_119_801 ();
 sg13g2_fill_2 FILLER_0_119_830 ();
 sg13g2_decap_8 FILLER_0_119_837 ();
 sg13g2_decap_4 FILLER_0_119_844 ();
 sg13g2_fill_2 FILLER_0_119_848 ();
 sg13g2_decap_4 FILLER_0_119_854 ();
 sg13g2_fill_1 FILLER_0_119_858 ();
 sg13g2_fill_2 FILLER_0_119_864 ();
 sg13g2_fill_2 FILLER_0_119_875 ();
 sg13g2_fill_1 FILLER_0_119_877 ();
 sg13g2_fill_1 FILLER_0_119_898 ();
 sg13g2_fill_1 FILLER_0_119_904 ();
 sg13g2_fill_1 FILLER_0_119_909 ();
 sg13g2_fill_1 FILLER_0_119_918 ();
 sg13g2_fill_1 FILLER_0_119_929 ();
 sg13g2_fill_1 FILLER_0_119_938 ();
 sg13g2_fill_1 FILLER_0_119_944 ();
 sg13g2_fill_1 FILLER_0_119_950 ();
 sg13g2_fill_1 FILLER_0_119_956 ();
 sg13g2_decap_4 FILLER_0_119_961 ();
 sg13g2_fill_2 FILLER_0_119_965 ();
 sg13g2_fill_2 FILLER_0_119_988 ();
 sg13g2_fill_1 FILLER_0_119_990 ();
 sg13g2_fill_1 FILLER_0_119_995 ();
 sg13g2_fill_2 FILLER_0_119_1037 ();
 sg13g2_fill_2 FILLER_0_119_1047 ();
 sg13g2_fill_2 FILLER_0_119_1054 ();
 sg13g2_decap_8 FILLER_0_119_1075 ();
 sg13g2_decap_8 FILLER_0_119_1082 ();
 sg13g2_decap_8 FILLER_0_119_1089 ();
 sg13g2_decap_8 FILLER_0_119_1096 ();
 sg13g2_decap_8 FILLER_0_119_1103 ();
 sg13g2_decap_8 FILLER_0_119_1110 ();
 sg13g2_decap_8 FILLER_0_119_1117 ();
 sg13g2_decap_8 FILLER_0_119_1124 ();
 sg13g2_decap_8 FILLER_0_119_1131 ();
 sg13g2_decap_8 FILLER_0_119_1138 ();
 sg13g2_decap_8 FILLER_0_119_1145 ();
 sg13g2_decap_8 FILLER_0_119_1152 ();
 sg13g2_decap_8 FILLER_0_119_1159 ();
 sg13g2_decap_8 FILLER_0_119_1166 ();
 sg13g2_decap_8 FILLER_0_119_1173 ();
 sg13g2_decap_8 FILLER_0_119_1180 ();
 sg13g2_decap_8 FILLER_0_119_1187 ();
 sg13g2_decap_8 FILLER_0_119_1194 ();
 sg13g2_decap_8 FILLER_0_119_1201 ();
 sg13g2_decap_8 FILLER_0_119_1208 ();
 sg13g2_decap_8 FILLER_0_119_1215 ();
 sg13g2_decap_4 FILLER_0_119_1222 ();
 sg13g2_fill_2 FILLER_0_119_1226 ();
 sg13g2_decap_8 FILLER_0_120_0 ();
 sg13g2_decap_8 FILLER_0_120_7 ();
 sg13g2_decap_8 FILLER_0_120_14 ();
 sg13g2_decap_8 FILLER_0_120_21 ();
 sg13g2_decap_8 FILLER_0_120_28 ();
 sg13g2_decap_8 FILLER_0_120_35 ();
 sg13g2_decap_8 FILLER_0_120_42 ();
 sg13g2_fill_2 FILLER_0_120_109 ();
 sg13g2_decap_8 FILLER_0_120_116 ();
 sg13g2_decap_8 FILLER_0_120_123 ();
 sg13g2_decap_8 FILLER_0_120_130 ();
 sg13g2_decap_8 FILLER_0_120_137 ();
 sg13g2_decap_8 FILLER_0_120_144 ();
 sg13g2_decap_8 FILLER_0_120_151 ();
 sg13g2_decap_8 FILLER_0_120_158 ();
 sg13g2_fill_2 FILLER_0_120_165 ();
 sg13g2_decap_8 FILLER_0_120_186 ();
 sg13g2_fill_1 FILLER_0_120_198 ();
 sg13g2_decap_8 FILLER_0_120_223 ();
 sg13g2_decap_8 FILLER_0_120_230 ();
 sg13g2_decap_8 FILLER_0_120_237 ();
 sg13g2_decap_8 FILLER_0_120_244 ();
 sg13g2_decap_8 FILLER_0_120_251 ();
 sg13g2_decap_8 FILLER_0_120_258 ();
 sg13g2_decap_8 FILLER_0_120_265 ();
 sg13g2_decap_8 FILLER_0_120_272 ();
 sg13g2_decap_8 FILLER_0_120_279 ();
 sg13g2_decap_8 FILLER_0_120_286 ();
 sg13g2_decap_8 FILLER_0_120_293 ();
 sg13g2_decap_8 FILLER_0_120_300 ();
 sg13g2_decap_8 FILLER_0_120_307 ();
 sg13g2_fill_2 FILLER_0_120_314 ();
 sg13g2_fill_1 FILLER_0_120_316 ();
 sg13g2_decap_4 FILLER_0_120_321 ();
 sg13g2_fill_1 FILLER_0_120_325 ();
 sg13g2_fill_2 FILLER_0_120_336 ();
 sg13g2_fill_1 FILLER_0_120_338 ();
 sg13g2_decap_4 FILLER_0_120_349 ();
 sg13g2_fill_1 FILLER_0_120_353 ();
 sg13g2_decap_8 FILLER_0_120_380 ();
 sg13g2_decap_8 FILLER_0_120_413 ();
 sg13g2_decap_4 FILLER_0_120_420 ();
 sg13g2_fill_1 FILLER_0_120_424 ();
 sg13g2_decap_8 FILLER_0_120_451 ();
 sg13g2_decap_4 FILLER_0_120_458 ();
 sg13g2_fill_1 FILLER_0_120_462 ();
 sg13g2_decap_8 FILLER_0_120_493 ();
 sg13g2_decap_4 FILLER_0_120_500 ();
 sg13g2_fill_2 FILLER_0_120_504 ();
 sg13g2_fill_2 FILLER_0_120_545 ();
 sg13g2_fill_1 FILLER_0_120_547 ();
 sg13g2_fill_1 FILLER_0_120_552 ();
 sg13g2_fill_1 FILLER_0_120_602 ();
 sg13g2_fill_1 FILLER_0_120_639 ();
 sg13g2_fill_2 FILLER_0_120_644 ();
 sg13g2_fill_2 FILLER_0_120_651 ();
 sg13g2_fill_2 FILLER_0_120_663 ();
 sg13g2_fill_1 FILLER_0_120_665 ();
 sg13g2_decap_8 FILLER_0_120_696 ();
 sg13g2_decap_8 FILLER_0_120_703 ();
 sg13g2_fill_2 FILLER_0_120_736 ();
 sg13g2_fill_2 FILLER_0_120_759 ();
 sg13g2_fill_2 FILLER_0_120_765 ();
 sg13g2_decap_4 FILLER_0_120_771 ();
 sg13g2_decap_8 FILLER_0_120_780 ();
 sg13g2_decap_4 FILLER_0_120_787 ();
 sg13g2_decap_8 FILLER_0_120_796 ();
 sg13g2_fill_1 FILLER_0_120_803 ();
 sg13g2_fill_1 FILLER_0_120_818 ();
 sg13g2_decap_8 FILLER_0_120_829 ();
 sg13g2_fill_2 FILLER_0_120_841 ();
 sg13g2_fill_1 FILLER_0_120_843 ();
 sg13g2_fill_2 FILLER_0_120_858 ();
 sg13g2_fill_2 FILLER_0_120_870 ();
 sg13g2_fill_2 FILLER_0_120_875 ();
 sg13g2_fill_1 FILLER_0_120_877 ();
 sg13g2_fill_1 FILLER_0_120_916 ();
 sg13g2_fill_2 FILLER_0_120_921 ();
 sg13g2_fill_1 FILLER_0_120_923 ();
 sg13g2_decap_8 FILLER_0_120_953 ();
 sg13g2_fill_1 FILLER_0_120_960 ();
 sg13g2_fill_1 FILLER_0_120_966 ();
 sg13g2_fill_2 FILLER_0_120_989 ();
 sg13g2_fill_1 FILLER_0_120_995 ();
 sg13g2_fill_1 FILLER_0_120_1005 ();
 sg13g2_fill_2 FILLER_0_120_1011 ();
 sg13g2_decap_8 FILLER_0_120_1048 ();
 sg13g2_decap_8 FILLER_0_120_1055 ();
 sg13g2_decap_4 FILLER_0_120_1062 ();
 sg13g2_fill_1 FILLER_0_120_1066 ();
 sg13g2_decap_8 FILLER_0_120_1097 ();
 sg13g2_decap_8 FILLER_0_120_1104 ();
 sg13g2_decap_8 FILLER_0_120_1111 ();
 sg13g2_decap_8 FILLER_0_120_1118 ();
 sg13g2_decap_8 FILLER_0_120_1125 ();
 sg13g2_decap_8 FILLER_0_120_1132 ();
 sg13g2_decap_8 FILLER_0_120_1139 ();
 sg13g2_decap_8 FILLER_0_120_1146 ();
 sg13g2_decap_8 FILLER_0_120_1153 ();
 sg13g2_decap_8 FILLER_0_120_1160 ();
 sg13g2_decap_8 FILLER_0_120_1167 ();
 sg13g2_decap_8 FILLER_0_120_1174 ();
 sg13g2_decap_8 FILLER_0_120_1181 ();
 sg13g2_decap_8 FILLER_0_120_1188 ();
 sg13g2_decap_8 FILLER_0_120_1195 ();
 sg13g2_decap_8 FILLER_0_120_1202 ();
 sg13g2_decap_8 FILLER_0_120_1209 ();
 sg13g2_decap_8 FILLER_0_120_1216 ();
 sg13g2_decap_4 FILLER_0_120_1223 ();
 sg13g2_fill_1 FILLER_0_120_1227 ();
 sg13g2_decap_8 FILLER_0_121_0 ();
 sg13g2_decap_8 FILLER_0_121_7 ();
 sg13g2_decap_8 FILLER_0_121_14 ();
 sg13g2_decap_8 FILLER_0_121_21 ();
 sg13g2_decap_8 FILLER_0_121_28 ();
 sg13g2_decap_8 FILLER_0_121_35 ();
 sg13g2_decap_8 FILLER_0_121_42 ();
 sg13g2_decap_4 FILLER_0_121_49 ();
 sg13g2_fill_1 FILLER_0_121_68 ();
 sg13g2_decap_8 FILLER_0_121_79 ();
 sg13g2_fill_1 FILLER_0_121_86 ();
 sg13g2_fill_2 FILLER_0_121_101 ();
 sg13g2_fill_1 FILLER_0_121_103 ();
 sg13g2_decap_8 FILLER_0_121_114 ();
 sg13g2_decap_8 FILLER_0_121_121 ();
 sg13g2_decap_8 FILLER_0_121_128 ();
 sg13g2_decap_8 FILLER_0_121_135 ();
 sg13g2_decap_8 FILLER_0_121_142 ();
 sg13g2_decap_4 FILLER_0_121_149 ();
 sg13g2_fill_2 FILLER_0_121_153 ();
 sg13g2_decap_4 FILLER_0_121_160 ();
 sg13g2_fill_1 FILLER_0_121_164 ();
 sg13g2_decap_4 FILLER_0_121_191 ();
 sg13g2_decap_8 FILLER_0_121_225 ();
 sg13g2_decap_8 FILLER_0_121_232 ();
 sg13g2_decap_8 FILLER_0_121_239 ();
 sg13g2_decap_8 FILLER_0_121_246 ();
 sg13g2_decap_8 FILLER_0_121_253 ();
 sg13g2_decap_8 FILLER_0_121_260 ();
 sg13g2_decap_8 FILLER_0_121_267 ();
 sg13g2_decap_8 FILLER_0_121_274 ();
 sg13g2_decap_8 FILLER_0_121_281 ();
 sg13g2_decap_8 FILLER_0_121_288 ();
 sg13g2_fill_2 FILLER_0_121_295 ();
 sg13g2_fill_1 FILLER_0_121_297 ();
 sg13g2_decap_4 FILLER_0_121_346 ();
 sg13g2_fill_1 FILLER_0_121_350 ();
 sg13g2_fill_2 FILLER_0_121_381 ();
 sg13g2_decap_4 FILLER_0_121_419 ();
 sg13g2_fill_2 FILLER_0_121_427 ();
 sg13g2_fill_2 FILLER_0_121_433 ();
 sg13g2_decap_4 FILLER_0_121_445 ();
 sg13g2_decap_8 FILLER_0_121_457 ();
 sg13g2_fill_1 FILLER_0_121_464 ();
 sg13g2_decap_8 FILLER_0_121_490 ();
 sg13g2_decap_8 FILLER_0_121_497 ();
 sg13g2_fill_2 FILLER_0_121_504 ();
 sg13g2_fill_2 FILLER_0_121_532 ();
 sg13g2_fill_2 FILLER_0_121_539 ();
 sg13g2_fill_2 FILLER_0_121_567 ();
 sg13g2_fill_1 FILLER_0_121_569 ();
 sg13g2_fill_2 FILLER_0_121_596 ();
 sg13g2_fill_1 FILLER_0_121_598 ();
 sg13g2_fill_1 FILLER_0_121_625 ();
 sg13g2_fill_2 FILLER_0_121_631 ();
 sg13g2_decap_4 FILLER_0_121_663 ();
 sg13g2_fill_1 FILLER_0_121_667 ();
 sg13g2_decap_8 FILLER_0_121_697 ();
 sg13g2_decap_8 FILLER_0_121_704 ();
 sg13g2_decap_4 FILLER_0_121_711 ();
 sg13g2_fill_1 FILLER_0_121_715 ();
 sg13g2_fill_1 FILLER_0_121_720 ();
 sg13g2_fill_1 FILLER_0_121_751 ();
 sg13g2_decap_4 FILLER_0_121_767 ();
 sg13g2_fill_1 FILLER_0_121_771 ();
 sg13g2_decap_8 FILLER_0_121_807 ();
 sg13g2_decap_8 FILLER_0_121_814 ();
 sg13g2_decap_8 FILLER_0_121_821 ();
 sg13g2_fill_1 FILLER_0_121_828 ();
 sg13g2_decap_4 FILLER_0_121_833 ();
 sg13g2_decap_8 FILLER_0_121_852 ();
 sg13g2_decap_4 FILLER_0_121_859 ();
 sg13g2_fill_2 FILLER_0_121_863 ();
 sg13g2_fill_1 FILLER_0_121_869 ();
 sg13g2_decap_4 FILLER_0_121_873 ();
 sg13g2_fill_1 FILLER_0_121_877 ();
 sg13g2_fill_2 FILLER_0_121_885 ();
 sg13g2_fill_1 FILLER_0_121_887 ();
 sg13g2_decap_4 FILLER_0_121_896 ();
 sg13g2_fill_2 FILLER_0_121_900 ();
 sg13g2_decap_8 FILLER_0_121_907 ();
 sg13g2_decap_4 FILLER_0_121_914 ();
 sg13g2_fill_2 FILLER_0_121_918 ();
 sg13g2_fill_1 FILLER_0_121_932 ();
 sg13g2_fill_1 FILLER_0_121_946 ();
 sg13g2_decap_8 FILLER_0_121_955 ();
 sg13g2_decap_8 FILLER_0_121_962 ();
 sg13g2_fill_2 FILLER_0_121_969 ();
 sg13g2_fill_1 FILLER_0_121_971 ();
 sg13g2_fill_1 FILLER_0_121_1044 ();
 sg13g2_decap_8 FILLER_0_121_1049 ();
 sg13g2_decap_8 FILLER_0_121_1056 ();
 sg13g2_decap_8 FILLER_0_121_1063 ();
 sg13g2_decap_8 FILLER_0_121_1070 ();
 sg13g2_fill_1 FILLER_0_121_1077 ();
 sg13g2_decap_8 FILLER_0_121_1096 ();
 sg13g2_decap_8 FILLER_0_121_1103 ();
 sg13g2_decap_8 FILLER_0_121_1110 ();
 sg13g2_decap_8 FILLER_0_121_1117 ();
 sg13g2_decap_8 FILLER_0_121_1124 ();
 sg13g2_decap_8 FILLER_0_121_1131 ();
 sg13g2_decap_8 FILLER_0_121_1138 ();
 sg13g2_decap_8 FILLER_0_121_1145 ();
 sg13g2_decap_8 FILLER_0_121_1152 ();
 sg13g2_decap_8 FILLER_0_121_1159 ();
 sg13g2_decap_8 FILLER_0_121_1166 ();
 sg13g2_decap_8 FILLER_0_121_1173 ();
 sg13g2_decap_8 FILLER_0_121_1180 ();
 sg13g2_decap_8 FILLER_0_121_1187 ();
 sg13g2_decap_8 FILLER_0_121_1194 ();
 sg13g2_decap_8 FILLER_0_121_1201 ();
 sg13g2_decap_8 FILLER_0_121_1208 ();
 sg13g2_decap_8 FILLER_0_121_1215 ();
 sg13g2_decap_4 FILLER_0_121_1222 ();
 sg13g2_fill_2 FILLER_0_121_1226 ();
 sg13g2_decap_8 FILLER_0_122_0 ();
 sg13g2_decap_8 FILLER_0_122_7 ();
 sg13g2_decap_8 FILLER_0_122_14 ();
 sg13g2_decap_8 FILLER_0_122_21 ();
 sg13g2_decap_8 FILLER_0_122_28 ();
 sg13g2_decap_8 FILLER_0_122_35 ();
 sg13g2_decap_8 FILLER_0_122_42 ();
 sg13g2_decap_8 FILLER_0_122_49 ();
 sg13g2_decap_8 FILLER_0_122_56 ();
 sg13g2_fill_2 FILLER_0_122_63 ();
 sg13g2_fill_1 FILLER_0_122_69 ();
 sg13g2_fill_1 FILLER_0_122_74 ();
 sg13g2_decap_4 FILLER_0_122_83 ();
 sg13g2_fill_1 FILLER_0_122_87 ();
 sg13g2_decap_8 FILLER_0_122_119 ();
 sg13g2_fill_2 FILLER_0_122_126 ();
 sg13g2_decap_8 FILLER_0_122_132 ();
 sg13g2_decap_4 FILLER_0_122_139 ();
 sg13g2_fill_1 FILLER_0_122_143 ();
 sg13g2_fill_1 FILLER_0_122_152 ();
 sg13g2_fill_1 FILLER_0_122_193 ();
 sg13g2_decap_8 FILLER_0_122_225 ();
 sg13g2_decap_8 FILLER_0_122_232 ();
 sg13g2_decap_8 FILLER_0_122_239 ();
 sg13g2_decap_8 FILLER_0_122_246 ();
 sg13g2_decap_8 FILLER_0_122_253 ();
 sg13g2_decap_8 FILLER_0_122_260 ();
 sg13g2_decap_8 FILLER_0_122_267 ();
 sg13g2_decap_8 FILLER_0_122_274 ();
 sg13g2_decap_8 FILLER_0_122_281 ();
 sg13g2_decap_8 FILLER_0_122_288 ();
 sg13g2_decap_4 FILLER_0_122_295 ();
 sg13g2_fill_2 FILLER_0_122_299 ();
 sg13g2_decap_4 FILLER_0_122_305 ();
 sg13g2_fill_1 FILLER_0_122_340 ();
 sg13g2_fill_2 FILLER_0_122_382 ();
 sg13g2_fill_1 FILLER_0_122_389 ();
 sg13g2_fill_1 FILLER_0_122_416 ();
 sg13g2_fill_2 FILLER_0_122_443 ();
 sg13g2_decap_4 FILLER_0_122_453 ();
 sg13g2_fill_2 FILLER_0_122_457 ();
 sg13g2_fill_2 FILLER_0_122_498 ();
 sg13g2_fill_1 FILLER_0_122_509 ();
 sg13g2_fill_2 FILLER_0_122_514 ();
 sg13g2_fill_1 FILLER_0_122_526 ();
 sg13g2_decap_8 FILLER_0_122_537 ();
 sg13g2_fill_1 FILLER_0_122_544 ();
 sg13g2_fill_2 FILLER_0_122_571 ();
 sg13g2_fill_1 FILLER_0_122_573 ();
 sg13g2_fill_2 FILLER_0_122_578 ();
 sg13g2_fill_1 FILLER_0_122_580 ();
 sg13g2_decap_8 FILLER_0_122_591 ();
 sg13g2_decap_4 FILLER_0_122_598 ();
 sg13g2_fill_1 FILLER_0_122_602 ();
 sg13g2_fill_2 FILLER_0_122_612 ();
 sg13g2_fill_1 FILLER_0_122_614 ();
 sg13g2_decap_8 FILLER_0_122_625 ();
 sg13g2_fill_1 FILLER_0_122_658 ();
 sg13g2_fill_1 FILLER_0_122_669 ();
 sg13g2_fill_1 FILLER_0_122_675 ();
 sg13g2_fill_1 FILLER_0_122_707 ();
 sg13g2_decap_8 FILLER_0_122_712 ();
 sg13g2_decap_8 FILLER_0_122_719 ();
 sg13g2_decap_4 FILLER_0_122_726 ();
 sg13g2_fill_1 FILLER_0_122_730 ();
 sg13g2_fill_1 FILLER_0_122_735 ();
 sg13g2_decap_4 FILLER_0_122_740 ();
 sg13g2_fill_1 FILLER_0_122_744 ();
 sg13g2_decap_4 FILLER_0_122_759 ();
 sg13g2_decap_8 FILLER_0_122_766 ();
 sg13g2_fill_1 FILLER_0_122_773 ();
 sg13g2_fill_2 FILLER_0_122_784 ();
 sg13g2_fill_2 FILLER_0_122_790 ();
 sg13g2_fill_1 FILLER_0_122_792 ();
 sg13g2_fill_2 FILLER_0_122_798 ();
 sg13g2_fill_1 FILLER_0_122_800 ();
 sg13g2_fill_2 FILLER_0_122_809 ();
 sg13g2_fill_2 FILLER_0_122_841 ();
 sg13g2_decap_8 FILLER_0_122_853 ();
 sg13g2_fill_1 FILLER_0_122_860 ();
 sg13g2_fill_2 FILLER_0_122_871 ();
 sg13g2_fill_1 FILLER_0_122_887 ();
 sg13g2_fill_1 FILLER_0_122_897 ();
 sg13g2_fill_1 FILLER_0_122_924 ();
 sg13g2_fill_1 FILLER_0_122_934 ();
 sg13g2_decap_4 FILLER_0_122_966 ();
 sg13g2_fill_2 FILLER_0_122_984 ();
 sg13g2_fill_2 FILLER_0_122_994 ();
 sg13g2_fill_1 FILLER_0_122_996 ();
 sg13g2_decap_8 FILLER_0_122_1043 ();
 sg13g2_decap_8 FILLER_0_122_1050 ();
 sg13g2_decap_8 FILLER_0_122_1057 ();
 sg13g2_fill_2 FILLER_0_122_1064 ();
 sg13g2_decap_8 FILLER_0_122_1097 ();
 sg13g2_decap_8 FILLER_0_122_1104 ();
 sg13g2_decap_8 FILLER_0_122_1111 ();
 sg13g2_decap_8 FILLER_0_122_1118 ();
 sg13g2_decap_8 FILLER_0_122_1125 ();
 sg13g2_decap_8 FILLER_0_122_1132 ();
 sg13g2_decap_8 FILLER_0_122_1139 ();
 sg13g2_decap_8 FILLER_0_122_1146 ();
 sg13g2_decap_8 FILLER_0_122_1153 ();
 sg13g2_decap_8 FILLER_0_122_1160 ();
 sg13g2_decap_8 FILLER_0_122_1167 ();
 sg13g2_decap_8 FILLER_0_122_1174 ();
 sg13g2_decap_8 FILLER_0_122_1181 ();
 sg13g2_decap_8 FILLER_0_122_1188 ();
 sg13g2_decap_8 FILLER_0_122_1195 ();
 sg13g2_decap_8 FILLER_0_122_1202 ();
 sg13g2_decap_8 FILLER_0_122_1209 ();
 sg13g2_decap_8 FILLER_0_122_1216 ();
 sg13g2_decap_4 FILLER_0_122_1223 ();
 sg13g2_fill_1 FILLER_0_122_1227 ();
 sg13g2_decap_8 FILLER_0_123_0 ();
 sg13g2_decap_8 FILLER_0_123_7 ();
 sg13g2_decap_8 FILLER_0_123_14 ();
 sg13g2_decap_8 FILLER_0_123_21 ();
 sg13g2_decap_8 FILLER_0_123_28 ();
 sg13g2_decap_8 FILLER_0_123_35 ();
 sg13g2_fill_1 FILLER_0_123_42 ();
 sg13g2_fill_2 FILLER_0_123_79 ();
 sg13g2_decap_4 FILLER_0_123_111 ();
 sg13g2_fill_2 FILLER_0_123_115 ();
 sg13g2_fill_1 FILLER_0_123_188 ();
 sg13g2_fill_1 FILLER_0_123_197 ();
 sg13g2_fill_1 FILLER_0_123_207 ();
 sg13g2_fill_1 FILLER_0_123_212 ();
 sg13g2_decap_8 FILLER_0_123_223 ();
 sg13g2_decap_8 FILLER_0_123_230 ();
 sg13g2_decap_8 FILLER_0_123_237 ();
 sg13g2_decap_8 FILLER_0_123_244 ();
 sg13g2_decap_8 FILLER_0_123_251 ();
 sg13g2_decap_8 FILLER_0_123_258 ();
 sg13g2_decap_8 FILLER_0_123_265 ();
 sg13g2_decap_8 FILLER_0_123_272 ();
 sg13g2_decap_8 FILLER_0_123_279 ();
 sg13g2_decap_8 FILLER_0_123_286 ();
 sg13g2_decap_8 FILLER_0_123_293 ();
 sg13g2_decap_8 FILLER_0_123_300 ();
 sg13g2_decap_8 FILLER_0_123_307 ();
 sg13g2_fill_2 FILLER_0_123_314 ();
 sg13g2_fill_1 FILLER_0_123_325 ();
 sg13g2_fill_1 FILLER_0_123_344 ();
 sg13g2_decap_4 FILLER_0_123_349 ();
 sg13g2_decap_8 FILLER_0_123_357 ();
 sg13g2_decap_4 FILLER_0_123_368 ();
 sg13g2_fill_1 FILLER_0_123_372 ();
 sg13g2_decap_4 FILLER_0_123_377 ();
 sg13g2_fill_2 FILLER_0_123_389 ();
 sg13g2_fill_2 FILLER_0_123_395 ();
 sg13g2_fill_2 FILLER_0_123_401 ();
 sg13g2_fill_2 FILLER_0_123_408 ();
 sg13g2_fill_1 FILLER_0_123_410 ();
 sg13g2_fill_1 FILLER_0_123_421 ();
 sg13g2_fill_2 FILLER_0_123_427 ();
 sg13g2_fill_1 FILLER_0_123_429 ();
 sg13g2_fill_2 FILLER_0_123_456 ();
 sg13g2_decap_8 FILLER_0_123_484 ();
 sg13g2_decap_8 FILLER_0_123_491 ();
 sg13g2_decap_4 FILLER_0_123_524 ();
 sg13g2_fill_2 FILLER_0_123_541 ();
 sg13g2_fill_1 FILLER_0_123_548 ();
 sg13g2_decap_8 FILLER_0_123_563 ();
 sg13g2_fill_2 FILLER_0_123_570 ();
 sg13g2_decap_4 FILLER_0_123_576 ();
 sg13g2_decap_4 FILLER_0_123_592 ();
 sg13g2_fill_1 FILLER_0_123_596 ();
 sg13g2_fill_2 FILLER_0_123_611 ();
 sg13g2_fill_1 FILLER_0_123_613 ();
 sg13g2_decap_4 FILLER_0_123_628 ();
 sg13g2_decap_8 FILLER_0_123_655 ();
 sg13g2_fill_2 FILLER_0_123_662 ();
 sg13g2_fill_1 FILLER_0_123_664 ();
 sg13g2_decap_4 FILLER_0_123_670 ();
 sg13g2_fill_1 FILLER_0_123_674 ();
 sg13g2_decap_8 FILLER_0_123_694 ();
 sg13g2_fill_1 FILLER_0_123_701 ();
 sg13g2_decap_8 FILLER_0_123_728 ();
 sg13g2_fill_1 FILLER_0_123_735 ();
 sg13g2_fill_1 FILLER_0_123_739 ();
 sg13g2_fill_2 FILLER_0_123_745 ();
 sg13g2_fill_1 FILLER_0_123_747 ();
 sg13g2_fill_2 FILLER_0_123_769 ();
 sg13g2_fill_1 FILLER_0_123_771 ();
 sg13g2_fill_2 FILLER_0_123_777 ();
 sg13g2_fill_1 FILLER_0_123_784 ();
 sg13g2_fill_2 FILLER_0_123_789 ();
 sg13g2_fill_2 FILLER_0_123_796 ();
 sg13g2_decap_8 FILLER_0_123_837 ();
 sg13g2_fill_1 FILLER_0_123_848 ();
 sg13g2_fill_1 FILLER_0_123_861 ();
 sg13g2_fill_1 FILLER_0_123_910 ();
 sg13g2_fill_2 FILLER_0_123_914 ();
 sg13g2_fill_2 FILLER_0_123_928 ();
 sg13g2_fill_1 FILLER_0_123_930 ();
 sg13g2_fill_2 FILLER_0_123_940 ();
 sg13g2_fill_1 FILLER_0_123_942 ();
 sg13g2_fill_1 FILLER_0_123_999 ();
 sg13g2_fill_2 FILLER_0_123_1035 ();
 sg13g2_decap_8 FILLER_0_123_1042 ();
 sg13g2_fill_1 FILLER_0_123_1049 ();
 sg13g2_decap_8 FILLER_0_123_1059 ();
 sg13g2_decap_8 FILLER_0_123_1066 ();
 sg13g2_fill_1 FILLER_0_123_1073 ();
 sg13g2_decap_8 FILLER_0_123_1123 ();
 sg13g2_decap_8 FILLER_0_123_1130 ();
 sg13g2_decap_8 FILLER_0_123_1137 ();
 sg13g2_decap_8 FILLER_0_123_1144 ();
 sg13g2_decap_8 FILLER_0_123_1151 ();
 sg13g2_decap_8 FILLER_0_123_1158 ();
 sg13g2_decap_8 FILLER_0_123_1165 ();
 sg13g2_decap_8 FILLER_0_123_1172 ();
 sg13g2_decap_8 FILLER_0_123_1179 ();
 sg13g2_decap_8 FILLER_0_123_1186 ();
 sg13g2_decap_8 FILLER_0_123_1193 ();
 sg13g2_decap_8 FILLER_0_123_1200 ();
 sg13g2_decap_8 FILLER_0_123_1207 ();
 sg13g2_decap_8 FILLER_0_123_1214 ();
 sg13g2_decap_8 FILLER_0_123_1221 ();
 sg13g2_decap_8 FILLER_0_124_0 ();
 sg13g2_decap_8 FILLER_0_124_7 ();
 sg13g2_decap_8 FILLER_0_124_14 ();
 sg13g2_decap_8 FILLER_0_124_21 ();
 sg13g2_decap_8 FILLER_0_124_28 ();
 sg13g2_decap_8 FILLER_0_124_35 ();
 sg13g2_fill_2 FILLER_0_124_42 ();
 sg13g2_decap_4 FILLER_0_124_84 ();
 sg13g2_fill_1 FILLER_0_124_88 ();
 sg13g2_decap_4 FILLER_0_124_108 ();
 sg13g2_fill_1 FILLER_0_124_112 ();
 sg13g2_decap_4 FILLER_0_124_124 ();
 sg13g2_fill_1 FILLER_0_124_128 ();
 sg13g2_fill_2 FILLER_0_124_173 ();
 sg13g2_fill_1 FILLER_0_124_175 ();
 sg13g2_fill_2 FILLER_0_124_186 ();
 sg13g2_decap_8 FILLER_0_124_228 ();
 sg13g2_decap_8 FILLER_0_124_235 ();
 sg13g2_decap_8 FILLER_0_124_242 ();
 sg13g2_decap_8 FILLER_0_124_249 ();
 sg13g2_decap_8 FILLER_0_124_256 ();
 sg13g2_decap_8 FILLER_0_124_263 ();
 sg13g2_decap_8 FILLER_0_124_270 ();
 sg13g2_decap_8 FILLER_0_124_277 ();
 sg13g2_decap_8 FILLER_0_124_284 ();
 sg13g2_decap_8 FILLER_0_124_291 ();
 sg13g2_decap_8 FILLER_0_124_298 ();
 sg13g2_decap_8 FILLER_0_124_305 ();
 sg13g2_decap_8 FILLER_0_124_312 ();
 sg13g2_decap_8 FILLER_0_124_319 ();
 sg13g2_decap_8 FILLER_0_124_326 ();
 sg13g2_decap_8 FILLER_0_124_340 ();
 sg13g2_decap_8 FILLER_0_124_347 ();
 sg13g2_fill_2 FILLER_0_124_354 ();
 sg13g2_decap_4 FILLER_0_124_364 ();
 sg13g2_decap_4 FILLER_0_124_390 ();
 sg13g2_fill_1 FILLER_0_124_394 ();
 sg13g2_decap_8 FILLER_0_124_417 ();
 sg13g2_decap_8 FILLER_0_124_424 ();
 sg13g2_decap_8 FILLER_0_124_431 ();
 sg13g2_decap_4 FILLER_0_124_438 ();
 sg13g2_fill_2 FILLER_0_124_442 ();
 sg13g2_decap_8 FILLER_0_124_480 ();
 sg13g2_decap_8 FILLER_0_124_487 ();
 sg13g2_fill_1 FILLER_0_124_494 ();
 sg13g2_decap_4 FILLER_0_124_504 ();
 sg13g2_decap_8 FILLER_0_124_518 ();
 sg13g2_fill_2 FILLER_0_124_525 ();
 sg13g2_fill_1 FILLER_0_124_527 ();
 sg13g2_decap_8 FILLER_0_124_546 ();
 sg13g2_decap_8 FILLER_0_124_563 ();
 sg13g2_decap_8 FILLER_0_124_570 ();
 sg13g2_decap_8 FILLER_0_124_577 ();
 sg13g2_decap_4 FILLER_0_124_629 ();
 sg13g2_fill_2 FILLER_0_124_663 ();
 sg13g2_fill_1 FILLER_0_124_665 ();
 sg13g2_decap_8 FILLER_0_124_700 ();
 sg13g2_fill_1 FILLER_0_124_707 ();
 sg13g2_fill_2 FILLER_0_124_734 ();
 sg13g2_fill_1 FILLER_0_124_736 ();
 sg13g2_fill_1 FILLER_0_124_767 ();
 sg13g2_fill_1 FILLER_0_124_777 ();
 sg13g2_fill_1 FILLER_0_124_791 ();
 sg13g2_fill_1 FILLER_0_124_816 ();
 sg13g2_decap_4 FILLER_0_124_822 ();
 sg13g2_fill_1 FILLER_0_124_826 ();
 sg13g2_fill_2 FILLER_0_124_832 ();
 sg13g2_fill_1 FILLER_0_124_834 ();
 sg13g2_fill_2 FILLER_0_124_864 ();
 sg13g2_fill_2 FILLER_0_124_873 ();
 sg13g2_fill_1 FILLER_0_124_898 ();
 sg13g2_fill_2 FILLER_0_124_904 ();
 sg13g2_fill_1 FILLER_0_124_926 ();
 sg13g2_fill_1 FILLER_0_124_936 ();
 sg13g2_fill_1 FILLER_0_124_977 ();
 sg13g2_fill_1 FILLER_0_124_988 ();
 sg13g2_fill_1 FILLER_0_124_992 ();
 sg13g2_fill_2 FILLER_0_124_998 ();
 sg13g2_fill_1 FILLER_0_124_1005 ();
 sg13g2_fill_1 FILLER_0_124_1011 ();
 sg13g2_decap_4 FILLER_0_124_1026 ();
 sg13g2_fill_2 FILLER_0_124_1030 ();
 sg13g2_decap_4 FILLER_0_124_1037 ();
 sg13g2_decap_8 FILLER_0_124_1067 ();
 sg13g2_fill_2 FILLER_0_124_1074 ();
 sg13g2_fill_1 FILLER_0_124_1076 ();
 sg13g2_decap_8 FILLER_0_124_1109 ();
 sg13g2_decap_8 FILLER_0_124_1116 ();
 sg13g2_decap_8 FILLER_0_124_1123 ();
 sg13g2_decap_8 FILLER_0_124_1130 ();
 sg13g2_decap_8 FILLER_0_124_1137 ();
 sg13g2_decap_8 FILLER_0_124_1144 ();
 sg13g2_decap_8 FILLER_0_124_1151 ();
 sg13g2_decap_8 FILLER_0_124_1158 ();
 sg13g2_decap_8 FILLER_0_124_1165 ();
 sg13g2_decap_8 FILLER_0_124_1172 ();
 sg13g2_decap_8 FILLER_0_124_1179 ();
 sg13g2_decap_8 FILLER_0_124_1186 ();
 sg13g2_decap_8 FILLER_0_124_1193 ();
 sg13g2_decap_8 FILLER_0_124_1200 ();
 sg13g2_decap_8 FILLER_0_124_1207 ();
 sg13g2_decap_8 FILLER_0_124_1214 ();
 sg13g2_decap_8 FILLER_0_124_1221 ();
 sg13g2_decap_8 FILLER_0_125_0 ();
 sg13g2_decap_8 FILLER_0_125_7 ();
 sg13g2_decap_8 FILLER_0_125_14 ();
 sg13g2_decap_8 FILLER_0_125_21 ();
 sg13g2_decap_8 FILLER_0_125_28 ();
 sg13g2_decap_4 FILLER_0_125_35 ();
 sg13g2_fill_1 FILLER_0_125_39 ();
 sg13g2_decap_4 FILLER_0_125_45 ();
 sg13g2_fill_1 FILLER_0_125_49 ();
 sg13g2_decap_8 FILLER_0_125_79 ();
 sg13g2_decap_8 FILLER_0_125_86 ();
 sg13g2_decap_8 FILLER_0_125_93 ();
 sg13g2_decap_8 FILLER_0_125_100 ();
 sg13g2_decap_8 FILLER_0_125_107 ();
 sg13g2_decap_4 FILLER_0_125_114 ();
 sg13g2_fill_2 FILLER_0_125_149 ();
 sg13g2_decap_4 FILLER_0_125_159 ();
 sg13g2_fill_1 FILLER_0_125_168 ();
 sg13g2_decap_8 FILLER_0_125_231 ();
 sg13g2_decap_8 FILLER_0_125_238 ();
 sg13g2_decap_8 FILLER_0_125_245 ();
 sg13g2_decap_8 FILLER_0_125_252 ();
 sg13g2_decap_8 FILLER_0_125_259 ();
 sg13g2_decap_8 FILLER_0_125_266 ();
 sg13g2_decap_8 FILLER_0_125_273 ();
 sg13g2_decap_8 FILLER_0_125_280 ();
 sg13g2_decap_8 FILLER_0_125_287 ();
 sg13g2_decap_8 FILLER_0_125_294 ();
 sg13g2_decap_8 FILLER_0_125_301 ();
 sg13g2_decap_8 FILLER_0_125_308 ();
 sg13g2_decap_8 FILLER_0_125_315 ();
 sg13g2_decap_8 FILLER_0_125_322 ();
 sg13g2_decap_8 FILLER_0_125_329 ();
 sg13g2_decap_8 FILLER_0_125_336 ();
 sg13g2_fill_2 FILLER_0_125_343 ();
 sg13g2_fill_1 FILLER_0_125_345 ();
 sg13g2_fill_2 FILLER_0_125_376 ();
 sg13g2_fill_1 FILLER_0_125_378 ();
 sg13g2_fill_2 FILLER_0_125_415 ();
 sg13g2_decap_8 FILLER_0_125_421 ();
 sg13g2_decap_4 FILLER_0_125_428 ();
 sg13g2_fill_1 FILLER_0_125_432 ();
 sg13g2_fill_1 FILLER_0_125_442 ();
 sg13g2_fill_2 FILLER_0_125_452 ();
 sg13g2_fill_2 FILLER_0_125_464 ();
 sg13g2_fill_1 FILLER_0_125_466 ();
 sg13g2_decap_8 FILLER_0_125_479 ();
 sg13g2_fill_1 FILLER_0_125_486 ();
 sg13g2_decap_4 FILLER_0_125_624 ();
 sg13g2_decap_8 FILLER_0_125_658 ();
 sg13g2_decap_4 FILLER_0_125_665 ();
 sg13g2_fill_1 FILLER_0_125_669 ();
 sg13g2_decap_8 FILLER_0_125_700 ();
 sg13g2_fill_2 FILLER_0_125_707 ();
 sg13g2_fill_1 FILLER_0_125_733 ();
 sg13g2_fill_1 FILLER_0_125_765 ();
 sg13g2_fill_1 FILLER_0_125_777 ();
 sg13g2_decap_4 FILLER_0_125_796 ();
 sg13g2_fill_2 FILLER_0_125_803 ();
 sg13g2_fill_1 FILLER_0_125_823 ();
 sg13g2_fill_1 FILLER_0_125_830 ();
 sg13g2_fill_1 FILLER_0_125_835 ();
 sg13g2_fill_1 FILLER_0_125_848 ();
 sg13g2_fill_2 FILLER_0_125_857 ();
 sg13g2_fill_1 FILLER_0_125_859 ();
 sg13g2_decap_4 FILLER_0_125_869 ();
 sg13g2_fill_2 FILLER_0_125_873 ();
 sg13g2_decap_4 FILLER_0_125_880 ();
 sg13g2_fill_2 FILLER_0_125_889 ();
 sg13g2_fill_1 FILLER_0_125_891 ();
 sg13g2_fill_1 FILLER_0_125_935 ();
 sg13g2_fill_1 FILLER_0_125_961 ();
 sg13g2_fill_2 FILLER_0_125_971 ();
 sg13g2_fill_2 FILLER_0_125_1014 ();
 sg13g2_fill_2 FILLER_0_125_1029 ();
 sg13g2_fill_1 FILLER_0_125_1049 ();
 sg13g2_fill_1 FILLER_0_125_1054 ();
 sg13g2_fill_1 FILLER_0_125_1076 ();
 sg13g2_decap_8 FILLER_0_125_1111 ();
 sg13g2_decap_8 FILLER_0_125_1118 ();
 sg13g2_decap_8 FILLER_0_125_1125 ();
 sg13g2_decap_8 FILLER_0_125_1132 ();
 sg13g2_decap_8 FILLER_0_125_1139 ();
 sg13g2_decap_8 FILLER_0_125_1146 ();
 sg13g2_decap_8 FILLER_0_125_1153 ();
 sg13g2_decap_8 FILLER_0_125_1160 ();
 sg13g2_decap_8 FILLER_0_125_1167 ();
 sg13g2_decap_8 FILLER_0_125_1174 ();
 sg13g2_decap_8 FILLER_0_125_1181 ();
 sg13g2_decap_8 FILLER_0_125_1188 ();
 sg13g2_decap_8 FILLER_0_125_1195 ();
 sg13g2_decap_8 FILLER_0_125_1202 ();
 sg13g2_decap_8 FILLER_0_125_1209 ();
 sg13g2_decap_8 FILLER_0_125_1216 ();
 sg13g2_decap_4 FILLER_0_125_1223 ();
 sg13g2_fill_1 FILLER_0_125_1227 ();
 sg13g2_decap_8 FILLER_0_126_0 ();
 sg13g2_decap_8 FILLER_0_126_7 ();
 sg13g2_decap_8 FILLER_0_126_14 ();
 sg13g2_decap_8 FILLER_0_126_21 ();
 sg13g2_decap_8 FILLER_0_126_28 ();
 sg13g2_decap_8 FILLER_0_126_35 ();
 sg13g2_decap_8 FILLER_0_126_92 ();
 sg13g2_decap_8 FILLER_0_126_99 ();
 sg13g2_decap_8 FILLER_0_126_106 ();
 sg13g2_decap_8 FILLER_0_126_113 ();
 sg13g2_decap_8 FILLER_0_126_120 ();
 sg13g2_decap_4 FILLER_0_126_127 ();
 sg13g2_fill_1 FILLER_0_126_131 ();
 sg13g2_fill_1 FILLER_0_126_136 ();
 sg13g2_fill_1 FILLER_0_126_163 ();
 sg13g2_decap_8 FILLER_0_126_225 ();
 sg13g2_decap_8 FILLER_0_126_232 ();
 sg13g2_decap_8 FILLER_0_126_239 ();
 sg13g2_decap_4 FILLER_0_126_246 ();
 sg13g2_decap_8 FILLER_0_126_256 ();
 sg13g2_decap_8 FILLER_0_126_263 ();
 sg13g2_decap_8 FILLER_0_126_270 ();
 sg13g2_decap_8 FILLER_0_126_277 ();
 sg13g2_decap_8 FILLER_0_126_284 ();
 sg13g2_decap_8 FILLER_0_126_291 ();
 sg13g2_decap_8 FILLER_0_126_298 ();
 sg13g2_decap_8 FILLER_0_126_305 ();
 sg13g2_decap_8 FILLER_0_126_312 ();
 sg13g2_decap_8 FILLER_0_126_319 ();
 sg13g2_decap_8 FILLER_0_126_326 ();
 sg13g2_decap_8 FILLER_0_126_333 ();
 sg13g2_decap_8 FILLER_0_126_340 ();
 sg13g2_decap_4 FILLER_0_126_347 ();
 sg13g2_fill_1 FILLER_0_126_433 ();
 sg13g2_decap_4 FILLER_0_126_444 ();
 sg13g2_fill_1 FILLER_0_126_448 ();
 sg13g2_decap_4 FILLER_0_126_459 ();
 sg13g2_fill_1 FILLER_0_126_463 ();
 sg13g2_decap_8 FILLER_0_126_469 ();
 sg13g2_fill_1 FILLER_0_126_476 ();
 sg13g2_fill_1 FILLER_0_126_523 ();
 sg13g2_decap_4 FILLER_0_126_528 ();
 sg13g2_decap_4 FILLER_0_126_562 ();
 sg13g2_fill_1 FILLER_0_126_566 ();
 sg13g2_fill_2 FILLER_0_126_597 ();
 sg13g2_fill_1 FILLER_0_126_599 ();
 sg13g2_decap_8 FILLER_0_126_626 ();
 sg13g2_decap_8 FILLER_0_126_659 ();
 sg13g2_fill_2 FILLER_0_126_666 ();
 sg13g2_fill_1 FILLER_0_126_668 ();
 sg13g2_decap_8 FILLER_0_126_702 ();
 sg13g2_decap_8 FILLER_0_126_709 ();
 sg13g2_fill_2 FILLER_0_126_734 ();
 sg13g2_fill_1 FILLER_0_126_748 ();
 sg13g2_fill_1 FILLER_0_126_767 ();
 sg13g2_fill_1 FILLER_0_126_772 ();
 sg13g2_decap_4 FILLER_0_126_779 ();
 sg13g2_fill_1 FILLER_0_126_809 ();
 sg13g2_fill_2 FILLER_0_126_851 ();
 sg13g2_fill_2 FILLER_0_126_858 ();
 sg13g2_fill_1 FILLER_0_126_875 ();
 sg13g2_fill_2 FILLER_0_126_894 ();
 sg13g2_fill_1 FILLER_0_126_917 ();
 sg13g2_fill_1 FILLER_0_126_925 ();
 sg13g2_fill_2 FILLER_0_126_965 ();
 sg13g2_fill_2 FILLER_0_126_972 ();
 sg13g2_fill_1 FILLER_0_126_974 ();
 sg13g2_fill_2 FILLER_0_126_1000 ();
 sg13g2_decap_8 FILLER_0_126_1022 ();
 sg13g2_decap_8 FILLER_0_126_1029 ();
 sg13g2_fill_1 FILLER_0_126_1036 ();
 sg13g2_fill_2 FILLER_0_126_1062 ();
 sg13g2_fill_1 FILLER_0_126_1064 ();
 sg13g2_fill_1 FILLER_0_126_1070 ();
 sg13g2_decap_4 FILLER_0_126_1079 ();
 sg13g2_decap_4 FILLER_0_126_1088 ();
 sg13g2_fill_2 FILLER_0_126_1092 ();
 sg13g2_decap_8 FILLER_0_126_1104 ();
 sg13g2_decap_8 FILLER_0_126_1111 ();
 sg13g2_decap_8 FILLER_0_126_1118 ();
 sg13g2_decap_8 FILLER_0_126_1125 ();
 sg13g2_decap_8 FILLER_0_126_1132 ();
 sg13g2_decap_8 FILLER_0_126_1139 ();
 sg13g2_decap_8 FILLER_0_126_1146 ();
 sg13g2_decap_8 FILLER_0_126_1153 ();
 sg13g2_decap_8 FILLER_0_126_1160 ();
 sg13g2_decap_8 FILLER_0_126_1167 ();
 sg13g2_decap_8 FILLER_0_126_1174 ();
 sg13g2_decap_8 FILLER_0_126_1181 ();
 sg13g2_decap_8 FILLER_0_126_1188 ();
 sg13g2_decap_8 FILLER_0_126_1195 ();
 sg13g2_decap_8 FILLER_0_126_1202 ();
 sg13g2_decap_8 FILLER_0_126_1209 ();
 sg13g2_decap_8 FILLER_0_126_1216 ();
 sg13g2_decap_4 FILLER_0_126_1223 ();
 sg13g2_fill_1 FILLER_0_126_1227 ();
 sg13g2_decap_8 FILLER_0_127_0 ();
 sg13g2_decap_8 FILLER_0_127_7 ();
 sg13g2_decap_8 FILLER_0_127_14 ();
 sg13g2_decap_8 FILLER_0_127_21 ();
 sg13g2_decap_8 FILLER_0_127_28 ();
 sg13g2_fill_1 FILLER_0_127_35 ();
 sg13g2_fill_1 FILLER_0_127_61 ();
 sg13g2_decap_8 FILLER_0_127_79 ();
 sg13g2_decap_8 FILLER_0_127_86 ();
 sg13g2_decap_8 FILLER_0_127_93 ();
 sg13g2_decap_8 FILLER_0_127_100 ();
 sg13g2_decap_8 FILLER_0_127_107 ();
 sg13g2_decap_8 FILLER_0_127_114 ();
 sg13g2_decap_8 FILLER_0_127_121 ();
 sg13g2_decap_4 FILLER_0_127_128 ();
 sg13g2_fill_2 FILLER_0_127_132 ();
 sg13g2_decap_4 FILLER_0_127_139 ();
 sg13g2_fill_1 FILLER_0_127_143 ();
 sg13g2_fill_2 FILLER_0_127_148 ();
 sg13g2_fill_1 FILLER_0_127_186 ();
 sg13g2_fill_1 FILLER_0_127_192 ();
 sg13g2_decap_4 FILLER_0_127_208 ();
 sg13g2_fill_1 FILLER_0_127_212 ();
 sg13g2_decap_8 FILLER_0_127_217 ();
 sg13g2_decap_8 FILLER_0_127_224 ();
 sg13g2_decap_8 FILLER_0_127_231 ();
 sg13g2_decap_8 FILLER_0_127_238 ();
 sg13g2_decap_8 FILLER_0_127_245 ();
 sg13g2_decap_8 FILLER_0_127_252 ();
 sg13g2_decap_8 FILLER_0_127_259 ();
 sg13g2_decap_8 FILLER_0_127_266 ();
 sg13g2_decap_8 FILLER_0_127_273 ();
 sg13g2_decap_8 FILLER_0_127_280 ();
 sg13g2_decap_8 FILLER_0_127_287 ();
 sg13g2_decap_8 FILLER_0_127_294 ();
 sg13g2_decap_8 FILLER_0_127_301 ();
 sg13g2_decap_8 FILLER_0_127_308 ();
 sg13g2_decap_8 FILLER_0_127_315 ();
 sg13g2_decap_8 FILLER_0_127_322 ();
 sg13g2_decap_8 FILLER_0_127_329 ();
 sg13g2_decap_4 FILLER_0_127_336 ();
 sg13g2_fill_2 FILLER_0_127_340 ();
 sg13g2_fill_1 FILLER_0_127_368 ();
 sg13g2_fill_2 FILLER_0_127_393 ();
 sg13g2_fill_2 FILLER_0_127_400 ();
 sg13g2_fill_1 FILLER_0_127_402 ();
 sg13g2_fill_2 FILLER_0_127_429 ();
 sg13g2_fill_1 FILLER_0_127_431 ();
 sg13g2_fill_2 FILLER_0_127_477 ();
 sg13g2_decap_8 FILLER_0_127_505 ();
 sg13g2_decap_8 FILLER_0_127_512 ();
 sg13g2_fill_2 FILLER_0_127_519 ();
 sg13g2_fill_1 FILLER_0_127_526 ();
 sg13g2_decap_8 FILLER_0_127_546 ();
 sg13g2_decap_8 FILLER_0_127_553 ();
 sg13g2_fill_2 FILLER_0_127_560 ();
 sg13g2_fill_1 FILLER_0_127_588 ();
 sg13g2_decap_8 FILLER_0_127_620 ();
 sg13g2_decap_8 FILLER_0_127_627 ();
 sg13g2_fill_2 FILLER_0_127_634 ();
 sg13g2_fill_1 FILLER_0_127_636 ();
 sg13g2_decap_8 FILLER_0_127_699 ();
 sg13g2_decap_8 FILLER_0_127_706 ();
 sg13g2_fill_2 FILLER_0_127_713 ();
 sg13g2_fill_2 FILLER_0_127_741 ();
 sg13g2_fill_1 FILLER_0_127_743 ();
 sg13g2_fill_2 FILLER_0_127_753 ();
 sg13g2_fill_1 FILLER_0_127_755 ();
 sg13g2_decap_4 FILLER_0_127_760 ();
 sg13g2_fill_1 FILLER_0_127_764 ();
 sg13g2_fill_1 FILLER_0_127_770 ();
 sg13g2_fill_2 FILLER_0_127_775 ();
 sg13g2_fill_1 FILLER_0_127_777 ();
 sg13g2_decap_8 FILLER_0_127_797 ();
 sg13g2_fill_2 FILLER_0_127_809 ();
 sg13g2_fill_2 FILLER_0_127_816 ();
 sg13g2_fill_2 FILLER_0_127_826 ();
 sg13g2_fill_1 FILLER_0_127_828 ();
 sg13g2_fill_2 FILLER_0_127_834 ();
 sg13g2_fill_1 FILLER_0_127_836 ();
 sg13g2_fill_2 FILLER_0_127_842 ();
 sg13g2_decap_8 FILLER_0_127_851 ();
 sg13g2_decap_8 FILLER_0_127_858 ();
 sg13g2_decap_8 FILLER_0_127_865 ();
 sg13g2_decap_8 FILLER_0_127_872 ();
 sg13g2_fill_2 FILLER_0_127_879 ();
 sg13g2_fill_1 FILLER_0_127_881 ();
 sg13g2_decap_8 FILLER_0_127_886 ();
 sg13g2_decap_8 FILLER_0_127_893 ();
 sg13g2_fill_2 FILLER_0_127_900 ();
 sg13g2_fill_1 FILLER_0_127_902 ();
 sg13g2_fill_2 FILLER_0_127_907 ();
 sg13g2_fill_2 FILLER_0_127_922 ();
 sg13g2_fill_1 FILLER_0_127_924 ();
 sg13g2_fill_2 FILLER_0_127_943 ();
 sg13g2_fill_1 FILLER_0_127_949 ();
 sg13g2_fill_1 FILLER_0_127_970 ();
 sg13g2_decap_4 FILLER_0_127_976 ();
 sg13g2_fill_2 FILLER_0_127_980 ();
 sg13g2_decap_4 FILLER_0_127_987 ();
 sg13g2_fill_1 FILLER_0_127_991 ();
 sg13g2_decap_4 FILLER_0_127_1004 ();
 sg13g2_fill_1 FILLER_0_127_1008 ();
 sg13g2_decap_4 FILLER_0_127_1022 ();
 sg13g2_fill_2 FILLER_0_127_1036 ();
 sg13g2_fill_1 FILLER_0_127_1043 ();
 sg13g2_decap_4 FILLER_0_127_1067 ();
 sg13g2_fill_1 FILLER_0_127_1081 ();
 sg13g2_decap_8 FILLER_0_127_1112 ();
 sg13g2_decap_8 FILLER_0_127_1119 ();
 sg13g2_decap_8 FILLER_0_127_1126 ();
 sg13g2_decap_8 FILLER_0_127_1133 ();
 sg13g2_decap_8 FILLER_0_127_1140 ();
 sg13g2_decap_8 FILLER_0_127_1147 ();
 sg13g2_decap_8 FILLER_0_127_1154 ();
 sg13g2_decap_8 FILLER_0_127_1161 ();
 sg13g2_decap_8 FILLER_0_127_1168 ();
 sg13g2_decap_8 FILLER_0_127_1175 ();
 sg13g2_decap_8 FILLER_0_127_1182 ();
 sg13g2_decap_8 FILLER_0_127_1189 ();
 sg13g2_decap_8 FILLER_0_127_1196 ();
 sg13g2_decap_8 FILLER_0_127_1203 ();
 sg13g2_decap_8 FILLER_0_127_1210 ();
 sg13g2_decap_8 FILLER_0_127_1217 ();
 sg13g2_decap_4 FILLER_0_127_1224 ();
 sg13g2_decap_8 FILLER_0_128_0 ();
 sg13g2_decap_8 FILLER_0_128_7 ();
 sg13g2_decap_8 FILLER_0_128_14 ();
 sg13g2_decap_8 FILLER_0_128_21 ();
 sg13g2_decap_8 FILLER_0_128_28 ();
 sg13g2_decap_8 FILLER_0_128_35 ();
 sg13g2_decap_8 FILLER_0_128_73 ();
 sg13g2_decap_8 FILLER_0_128_80 ();
 sg13g2_decap_8 FILLER_0_128_87 ();
 sg13g2_decap_8 FILLER_0_128_94 ();
 sg13g2_decap_8 FILLER_0_128_105 ();
 sg13g2_decap_8 FILLER_0_128_112 ();
 sg13g2_decap_8 FILLER_0_128_119 ();
 sg13g2_decap_4 FILLER_0_128_126 ();
 sg13g2_fill_2 FILLER_0_128_130 ();
 sg13g2_decap_8 FILLER_0_128_151 ();
 sg13g2_fill_2 FILLER_0_128_158 ();
 sg13g2_fill_2 FILLER_0_128_170 ();
 sg13g2_fill_1 FILLER_0_128_172 ();
 sg13g2_fill_1 FILLER_0_128_182 ();
 sg13g2_decap_8 FILLER_0_128_187 ();
 sg13g2_fill_2 FILLER_0_128_194 ();
 sg13g2_decap_8 FILLER_0_128_200 ();
 sg13g2_decap_8 FILLER_0_128_207 ();
 sg13g2_decap_8 FILLER_0_128_214 ();
 sg13g2_decap_8 FILLER_0_128_221 ();
 sg13g2_decap_8 FILLER_0_128_228 ();
 sg13g2_decap_8 FILLER_0_128_235 ();
 sg13g2_decap_8 FILLER_0_128_242 ();
 sg13g2_decap_8 FILLER_0_128_249 ();
 sg13g2_decap_8 FILLER_0_128_256 ();
 sg13g2_decap_8 FILLER_0_128_263 ();
 sg13g2_decap_8 FILLER_0_128_270 ();
 sg13g2_decap_8 FILLER_0_128_277 ();
 sg13g2_decap_8 FILLER_0_128_284 ();
 sg13g2_decap_8 FILLER_0_128_291 ();
 sg13g2_decap_8 FILLER_0_128_298 ();
 sg13g2_decap_8 FILLER_0_128_305 ();
 sg13g2_decap_8 FILLER_0_128_312 ();
 sg13g2_decap_8 FILLER_0_128_319 ();
 sg13g2_decap_8 FILLER_0_128_326 ();
 sg13g2_decap_8 FILLER_0_128_333 ();
 sg13g2_fill_2 FILLER_0_128_340 ();
 sg13g2_fill_1 FILLER_0_128_342 ();
 sg13g2_fill_1 FILLER_0_128_352 ();
 sg13g2_decap_8 FILLER_0_128_373 ();
 sg13g2_decap_8 FILLER_0_128_380 ();
 sg13g2_decap_8 FILLER_0_128_387 ();
 sg13g2_decap_8 FILLER_0_128_394 ();
 sg13g2_decap_4 FILLER_0_128_405 ();
 sg13g2_fill_2 FILLER_0_128_419 ();
 sg13g2_fill_1 FILLER_0_128_421 ();
 sg13g2_decap_4 FILLER_0_128_427 ();
 sg13g2_fill_2 FILLER_0_128_431 ();
 sg13g2_fill_2 FILLER_0_128_438 ();
 sg13g2_fill_2 FILLER_0_128_444 ();
 sg13g2_fill_1 FILLER_0_128_446 ();
 sg13g2_fill_2 FILLER_0_128_492 ();
 sg13g2_decap_8 FILLER_0_128_498 ();
 sg13g2_decap_8 FILLER_0_128_505 ();
 sg13g2_decap_4 FILLER_0_128_512 ();
 sg13g2_fill_2 FILLER_0_128_516 ();
 sg13g2_decap_8 FILLER_0_128_537 ();
 sg13g2_decap_8 FILLER_0_128_544 ();
 sg13g2_decap_8 FILLER_0_128_551 ();
 sg13g2_decap_8 FILLER_0_128_558 ();
 sg13g2_decap_4 FILLER_0_128_565 ();
 sg13g2_fill_1 FILLER_0_128_569 ();
 sg13g2_decap_4 FILLER_0_128_575 ();
 sg13g2_fill_2 FILLER_0_128_579 ();
 sg13g2_decap_8 FILLER_0_128_591 ();
 sg13g2_decap_4 FILLER_0_128_598 ();
 sg13g2_fill_2 FILLER_0_128_602 ();
 sg13g2_fill_2 FILLER_0_128_642 ();
 sg13g2_fill_1 FILLER_0_128_644 ();
 sg13g2_decap_4 FILLER_0_128_650 ();
 sg13g2_fill_1 FILLER_0_128_654 ();
 sg13g2_fill_2 FILLER_0_128_659 ();
 sg13g2_fill_1 FILLER_0_128_661 ();
 sg13g2_decap_8 FILLER_0_128_666 ();
 sg13g2_fill_1 FILLER_0_128_678 ();
 sg13g2_decap_8 FILLER_0_128_691 ();
 sg13g2_decap_8 FILLER_0_128_698 ();
 sg13g2_decap_8 FILLER_0_128_705 ();
 sg13g2_decap_8 FILLER_0_128_712 ();
 sg13g2_fill_2 FILLER_0_128_719 ();
 sg13g2_decap_8 FILLER_0_128_725 ();
 sg13g2_decap_4 FILLER_0_128_732 ();
 sg13g2_fill_1 FILLER_0_128_740 ();
 sg13g2_fill_1 FILLER_0_128_755 ();
 sg13g2_decap_4 FILLER_0_128_771 ();
 sg13g2_fill_1 FILLER_0_128_775 ();
 sg13g2_fill_2 FILLER_0_128_786 ();
 sg13g2_decap_8 FILLER_0_128_796 ();
 sg13g2_decap_8 FILLER_0_128_803 ();
 sg13g2_decap_8 FILLER_0_128_810 ();
 sg13g2_decap_8 FILLER_0_128_817 ();
 sg13g2_fill_2 FILLER_0_128_824 ();
 sg13g2_fill_1 FILLER_0_128_826 ();
 sg13g2_decap_4 FILLER_0_128_851 ();
 sg13g2_decap_8 FILLER_0_128_863 ();
 sg13g2_fill_1 FILLER_0_128_870 ();
 sg13g2_decap_4 FILLER_0_128_880 ();
 sg13g2_decap_8 FILLER_0_128_892 ();
 sg13g2_fill_2 FILLER_0_128_899 ();
 sg13g2_decap_8 FILLER_0_128_916 ();
 sg13g2_fill_1 FILLER_0_128_923 ();
 sg13g2_fill_2 FILLER_0_128_928 ();
 sg13g2_fill_1 FILLER_0_128_939 ();
 sg13g2_decap_8 FILLER_0_128_954 ();
 sg13g2_fill_2 FILLER_0_128_961 ();
 sg13g2_fill_1 FILLER_0_128_963 ();
 sg13g2_decap_8 FILLER_0_128_968 ();
 sg13g2_decap_8 FILLER_0_128_975 ();
 sg13g2_decap_4 FILLER_0_128_982 ();
 sg13g2_fill_2 FILLER_0_128_986 ();
 sg13g2_fill_1 FILLER_0_128_1003 ();
 sg13g2_decap_8 FILLER_0_128_1022 ();
 sg13g2_decap_4 FILLER_0_128_1029 ();
 sg13g2_decap_4 FILLER_0_128_1043 ();
 sg13g2_fill_2 FILLER_0_128_1055 ();
 sg13g2_fill_2 FILLER_0_128_1073 ();
 sg13g2_fill_1 FILLER_0_128_1075 ();
 sg13g2_decap_4 FILLER_0_128_1081 ();
 sg13g2_fill_2 FILLER_0_128_1090 ();
 sg13g2_fill_1 FILLER_0_128_1092 ();
 sg13g2_decap_8 FILLER_0_128_1103 ();
 sg13g2_decap_8 FILLER_0_128_1110 ();
 sg13g2_decap_8 FILLER_0_128_1117 ();
 sg13g2_decap_8 FILLER_0_128_1124 ();
 sg13g2_decap_8 FILLER_0_128_1131 ();
 sg13g2_decap_8 FILLER_0_128_1138 ();
 sg13g2_decap_8 FILLER_0_128_1145 ();
 sg13g2_decap_8 FILLER_0_128_1152 ();
 sg13g2_decap_8 FILLER_0_128_1159 ();
 sg13g2_decap_8 FILLER_0_128_1166 ();
 sg13g2_decap_8 FILLER_0_128_1173 ();
 sg13g2_decap_8 FILLER_0_128_1180 ();
 sg13g2_decap_8 FILLER_0_128_1187 ();
 sg13g2_decap_8 FILLER_0_128_1194 ();
 sg13g2_decap_8 FILLER_0_128_1201 ();
 sg13g2_decap_8 FILLER_0_128_1208 ();
 sg13g2_decap_8 FILLER_0_128_1215 ();
 sg13g2_decap_4 FILLER_0_128_1222 ();
 sg13g2_fill_2 FILLER_0_128_1226 ();
 sg13g2_decap_8 FILLER_0_129_0 ();
 sg13g2_decap_8 FILLER_0_129_7 ();
 sg13g2_decap_8 FILLER_0_129_14 ();
 sg13g2_decap_8 FILLER_0_129_21 ();
 sg13g2_decap_8 FILLER_0_129_28 ();
 sg13g2_fill_1 FILLER_0_129_35 ();
 sg13g2_decap_8 FILLER_0_129_77 ();
 sg13g2_decap_8 FILLER_0_129_84 ();
 sg13g2_decap_8 FILLER_0_129_91 ();
 sg13g2_decap_8 FILLER_0_129_98 ();
 sg13g2_decap_8 FILLER_0_129_105 ();
 sg13g2_decap_4 FILLER_0_129_112 ();
 sg13g2_fill_2 FILLER_0_129_161 ();
 sg13g2_decap_8 FILLER_0_129_173 ();
 sg13g2_decap_8 FILLER_0_129_180 ();
 sg13g2_decap_8 FILLER_0_129_187 ();
 sg13g2_decap_8 FILLER_0_129_194 ();
 sg13g2_decap_8 FILLER_0_129_201 ();
 sg13g2_decap_8 FILLER_0_129_208 ();
 sg13g2_decap_8 FILLER_0_129_215 ();
 sg13g2_decap_8 FILLER_0_129_222 ();
 sg13g2_decap_8 FILLER_0_129_229 ();
 sg13g2_decap_8 FILLER_0_129_236 ();
 sg13g2_decap_8 FILLER_0_129_243 ();
 sg13g2_decap_8 FILLER_0_129_250 ();
 sg13g2_decap_8 FILLER_0_129_257 ();
 sg13g2_decap_8 FILLER_0_129_264 ();
 sg13g2_decap_8 FILLER_0_129_271 ();
 sg13g2_decap_8 FILLER_0_129_278 ();
 sg13g2_decap_8 FILLER_0_129_285 ();
 sg13g2_decap_8 FILLER_0_129_292 ();
 sg13g2_decap_8 FILLER_0_129_299 ();
 sg13g2_decap_8 FILLER_0_129_306 ();
 sg13g2_decap_8 FILLER_0_129_313 ();
 sg13g2_decap_8 FILLER_0_129_320 ();
 sg13g2_decap_8 FILLER_0_129_327 ();
 sg13g2_decap_8 FILLER_0_129_334 ();
 sg13g2_fill_1 FILLER_0_129_341 ();
 sg13g2_decap_8 FILLER_0_129_373 ();
 sg13g2_decap_8 FILLER_0_129_380 ();
 sg13g2_fill_2 FILLER_0_129_387 ();
 sg13g2_fill_1 FILLER_0_129_389 ();
 sg13g2_decap_8 FILLER_0_129_434 ();
 sg13g2_decap_8 FILLER_0_129_441 ();
 sg13g2_decap_8 FILLER_0_129_448 ();
 sg13g2_fill_1 FILLER_0_129_455 ();
 sg13g2_decap_8 FILLER_0_129_482 ();
 sg13g2_decap_8 FILLER_0_129_489 ();
 sg13g2_decap_8 FILLER_0_129_496 ();
 sg13g2_fill_1 FILLER_0_129_503 ();
 sg13g2_decap_4 FILLER_0_129_508 ();
 sg13g2_fill_1 FILLER_0_129_512 ();
 sg13g2_fill_2 FILLER_0_129_518 ();
 sg13g2_fill_1 FILLER_0_129_520 ();
 sg13g2_decap_4 FILLER_0_129_547 ();
 sg13g2_fill_1 FILLER_0_129_551 ();
 sg13g2_decap_8 FILLER_0_129_578 ();
 sg13g2_decap_8 FILLER_0_129_585 ();
 sg13g2_decap_8 FILLER_0_129_592 ();
 sg13g2_decap_8 FILLER_0_129_599 ();
 sg13g2_decap_8 FILLER_0_129_708 ();
 sg13g2_decap_4 FILLER_0_129_715 ();
 sg13g2_fill_2 FILLER_0_129_719 ();
 sg13g2_decap_4 FILLER_0_129_725 ();
 sg13g2_fill_2 FILLER_0_129_729 ();
 sg13g2_decap_8 FILLER_0_129_741 ();
 sg13g2_fill_2 FILLER_0_129_748 ();
 sg13g2_fill_1 FILLER_0_129_754 ();
 sg13g2_fill_1 FILLER_0_129_758 ();
 sg13g2_fill_1 FILLER_0_129_764 ();
 sg13g2_fill_2 FILLER_0_129_780 ();
 sg13g2_fill_1 FILLER_0_129_782 ();
 sg13g2_fill_1 FILLER_0_129_787 ();
 sg13g2_decap_4 FILLER_0_129_792 ();
 sg13g2_fill_2 FILLER_0_129_796 ();
 sg13g2_fill_2 FILLER_0_129_806 ();
 sg13g2_decap_4 FILLER_0_129_818 ();
 sg13g2_fill_1 FILLER_0_129_822 ();
 sg13g2_fill_2 FILLER_0_129_833 ();
 sg13g2_fill_1 FILLER_0_129_835 ();
 sg13g2_decap_8 FILLER_0_129_846 ();
 sg13g2_fill_1 FILLER_0_129_869 ();
 sg13g2_fill_2 FILLER_0_129_880 ();
 sg13g2_fill_2 FILLER_0_129_889 ();
 sg13g2_fill_1 FILLER_0_129_891 ();
 sg13g2_fill_2 FILLER_0_129_896 ();
 sg13g2_fill_1 FILLER_0_129_898 ();
 sg13g2_decap_4 FILLER_0_129_904 ();
 sg13g2_fill_2 FILLER_0_129_908 ();
 sg13g2_fill_2 FILLER_0_129_924 ();
 sg13g2_fill_1 FILLER_0_129_926 ();
 sg13g2_fill_1 FILLER_0_129_937 ();
 sg13g2_fill_1 FILLER_0_129_942 ();
 sg13g2_fill_1 FILLER_0_129_952 ();
 sg13g2_fill_1 FILLER_0_129_964 ();
 sg13g2_fill_1 FILLER_0_129_970 ();
 sg13g2_fill_2 FILLER_0_129_992 ();
 sg13g2_fill_1 FILLER_0_129_1000 ();
 sg13g2_fill_1 FILLER_0_129_1006 ();
 sg13g2_fill_1 FILLER_0_129_1012 ();
 sg13g2_fill_1 FILLER_0_129_1018 ();
 sg13g2_decap_8 FILLER_0_129_1025 ();
 sg13g2_fill_2 FILLER_0_129_1058 ();
 sg13g2_decap_8 FILLER_0_129_1065 ();
 sg13g2_decap_8 FILLER_0_129_1072 ();
 sg13g2_fill_2 FILLER_0_129_1079 ();
 sg13g2_fill_1 FILLER_0_129_1081 ();
 sg13g2_decap_8 FILLER_0_129_1112 ();
 sg13g2_decap_8 FILLER_0_129_1119 ();
 sg13g2_decap_8 FILLER_0_129_1126 ();
 sg13g2_decap_8 FILLER_0_129_1133 ();
 sg13g2_decap_8 FILLER_0_129_1140 ();
 sg13g2_decap_8 FILLER_0_129_1147 ();
 sg13g2_decap_8 FILLER_0_129_1154 ();
 sg13g2_decap_8 FILLER_0_129_1161 ();
 sg13g2_decap_8 FILLER_0_129_1168 ();
 sg13g2_decap_8 FILLER_0_129_1175 ();
 sg13g2_decap_8 FILLER_0_129_1182 ();
 sg13g2_decap_8 FILLER_0_129_1189 ();
 sg13g2_decap_8 FILLER_0_129_1196 ();
 sg13g2_decap_8 FILLER_0_129_1203 ();
 sg13g2_decap_8 FILLER_0_129_1210 ();
 sg13g2_decap_8 FILLER_0_129_1217 ();
 sg13g2_decap_4 FILLER_0_129_1224 ();
 sg13g2_decap_8 FILLER_0_130_0 ();
 sg13g2_decap_8 FILLER_0_130_7 ();
 sg13g2_decap_8 FILLER_0_130_14 ();
 sg13g2_decap_8 FILLER_0_130_21 ();
 sg13g2_decap_8 FILLER_0_130_28 ();
 sg13g2_decap_8 FILLER_0_130_35 ();
 sg13g2_decap_8 FILLER_0_130_42 ();
 sg13g2_fill_2 FILLER_0_130_49 ();
 sg13g2_fill_1 FILLER_0_130_51 ();
 sg13g2_decap_4 FILLER_0_130_56 ();
 sg13g2_fill_2 FILLER_0_130_60 ();
 sg13g2_decap_8 FILLER_0_130_72 ();
 sg13g2_decap_8 FILLER_0_130_79 ();
 sg13g2_decap_8 FILLER_0_130_86 ();
 sg13g2_decap_8 FILLER_0_130_93 ();
 sg13g2_decap_8 FILLER_0_130_100 ();
 sg13g2_decap_8 FILLER_0_130_107 ();
 sg13g2_fill_1 FILLER_0_130_114 ();
 sg13g2_decap_8 FILLER_0_130_177 ();
 sg13g2_decap_8 FILLER_0_130_184 ();
 sg13g2_decap_8 FILLER_0_130_191 ();
 sg13g2_decap_8 FILLER_0_130_198 ();
 sg13g2_decap_8 FILLER_0_130_205 ();
 sg13g2_decap_8 FILLER_0_130_212 ();
 sg13g2_decap_8 FILLER_0_130_219 ();
 sg13g2_decap_8 FILLER_0_130_226 ();
 sg13g2_decap_8 FILLER_0_130_233 ();
 sg13g2_decap_8 FILLER_0_130_240 ();
 sg13g2_decap_8 FILLER_0_130_247 ();
 sg13g2_decap_8 FILLER_0_130_254 ();
 sg13g2_decap_8 FILLER_0_130_261 ();
 sg13g2_decap_8 FILLER_0_130_268 ();
 sg13g2_decap_8 FILLER_0_130_275 ();
 sg13g2_decap_8 FILLER_0_130_282 ();
 sg13g2_decap_8 FILLER_0_130_289 ();
 sg13g2_decap_8 FILLER_0_130_296 ();
 sg13g2_decap_8 FILLER_0_130_303 ();
 sg13g2_decap_8 FILLER_0_130_310 ();
 sg13g2_decap_8 FILLER_0_130_317 ();
 sg13g2_decap_8 FILLER_0_130_324 ();
 sg13g2_decap_8 FILLER_0_130_331 ();
 sg13g2_decap_4 FILLER_0_130_338 ();
 sg13g2_fill_1 FILLER_0_130_347 ();
 sg13g2_fill_1 FILLER_0_130_374 ();
 sg13g2_fill_1 FILLER_0_130_379 ();
 sg13g2_fill_2 FILLER_0_130_415 ();
 sg13g2_decap_8 FILLER_0_130_421 ();
 sg13g2_decap_8 FILLER_0_130_428 ();
 sg13g2_decap_8 FILLER_0_130_435 ();
 sg13g2_decap_4 FILLER_0_130_442 ();
 sg13g2_fill_1 FILLER_0_130_446 ();
 sg13g2_fill_2 FILLER_0_130_465 ();
 sg13g2_fill_1 FILLER_0_130_467 ();
 sg13g2_fill_1 FILLER_0_130_472 ();
 sg13g2_fill_1 FILLER_0_130_493 ();
 sg13g2_decap_4 FILLER_0_130_543 ();
 sg13g2_fill_2 FILLER_0_130_547 ();
 sg13g2_decap_8 FILLER_0_130_594 ();
 sg13g2_decap_4 FILLER_0_130_601 ();
 sg13g2_decap_8 FILLER_0_130_636 ();
 sg13g2_decap_8 FILLER_0_130_643 ();
 sg13g2_decap_8 FILLER_0_130_650 ();
 sg13g2_fill_1 FILLER_0_130_657 ();
 sg13g2_decap_4 FILLER_0_130_663 ();
 sg13g2_fill_2 FILLER_0_130_667 ();
 sg13g2_decap_8 FILLER_0_130_694 ();
 sg13g2_decap_8 FILLER_0_130_701 ();
 sg13g2_decap_4 FILLER_0_130_708 ();
 sg13g2_fill_1 FILLER_0_130_779 ();
 sg13g2_fill_1 FILLER_0_130_785 ();
 sg13g2_decap_4 FILLER_0_130_790 ();
 sg13g2_fill_1 FILLER_0_130_794 ();
 sg13g2_fill_1 FILLER_0_130_804 ();
 sg13g2_fill_2 FILLER_0_130_810 ();
 sg13g2_fill_2 FILLER_0_130_824 ();
 sg13g2_fill_1 FILLER_0_130_826 ();
 sg13g2_fill_1 FILLER_0_130_839 ();
 sg13g2_fill_2 FILLER_0_130_844 ();
 sg13g2_fill_2 FILLER_0_130_883 ();
 sg13g2_fill_2 FILLER_0_130_890 ();
 sg13g2_fill_1 FILLER_0_130_892 ();
 sg13g2_fill_1 FILLER_0_130_920 ();
 sg13g2_fill_2 FILLER_0_130_969 ();
 sg13g2_fill_1 FILLER_0_130_971 ();
 sg13g2_fill_1 FILLER_0_130_1000 ();
 sg13g2_fill_2 FILLER_0_130_1005 ();
 sg13g2_fill_1 FILLER_0_130_1007 ();
 sg13g2_fill_2 FILLER_0_130_1013 ();
 sg13g2_fill_1 FILLER_0_130_1015 ();
 sg13g2_decap_8 FILLER_0_130_1025 ();
 sg13g2_fill_2 FILLER_0_130_1032 ();
 sg13g2_fill_2 FILLER_0_130_1043 ();
 sg13g2_fill_1 FILLER_0_130_1053 ();
 sg13g2_decap_8 FILLER_0_130_1058 ();
 sg13g2_decap_8 FILLER_0_130_1065 ();
 sg13g2_decap_4 FILLER_0_130_1072 ();
 sg13g2_fill_1 FILLER_0_130_1076 ();
 sg13g2_fill_1 FILLER_0_130_1086 ();
 sg13g2_decap_8 FILLER_0_130_1101 ();
 sg13g2_decap_8 FILLER_0_130_1108 ();
 sg13g2_decap_8 FILLER_0_130_1115 ();
 sg13g2_decap_8 FILLER_0_130_1122 ();
 sg13g2_decap_8 FILLER_0_130_1129 ();
 sg13g2_decap_8 FILLER_0_130_1136 ();
 sg13g2_decap_8 FILLER_0_130_1143 ();
 sg13g2_decap_8 FILLER_0_130_1150 ();
 sg13g2_decap_8 FILLER_0_130_1157 ();
 sg13g2_decap_8 FILLER_0_130_1164 ();
 sg13g2_decap_8 FILLER_0_130_1171 ();
 sg13g2_decap_8 FILLER_0_130_1178 ();
 sg13g2_decap_8 FILLER_0_130_1185 ();
 sg13g2_decap_8 FILLER_0_130_1192 ();
 sg13g2_decap_8 FILLER_0_130_1199 ();
 sg13g2_decap_8 FILLER_0_130_1206 ();
 sg13g2_decap_8 FILLER_0_130_1213 ();
 sg13g2_decap_8 FILLER_0_130_1220 ();
 sg13g2_fill_1 FILLER_0_130_1227 ();
 sg13g2_decap_8 FILLER_0_131_0 ();
 sg13g2_decap_8 FILLER_0_131_7 ();
 sg13g2_decap_8 FILLER_0_131_14 ();
 sg13g2_decap_8 FILLER_0_131_21 ();
 sg13g2_decap_8 FILLER_0_131_28 ();
 sg13g2_fill_2 FILLER_0_131_35 ();
 sg13g2_fill_1 FILLER_0_131_37 ();
 sg13g2_decap_8 FILLER_0_131_73 ();
 sg13g2_decap_8 FILLER_0_131_80 ();
 sg13g2_fill_1 FILLER_0_131_87 ();
 sg13g2_fill_2 FILLER_0_131_114 ();
 sg13g2_fill_2 FILLER_0_131_150 ();
 sg13g2_fill_1 FILLER_0_131_152 ();
 sg13g2_fill_2 FILLER_0_131_157 ();
 sg13g2_decap_8 FILLER_0_131_199 ();
 sg13g2_decap_8 FILLER_0_131_206 ();
 sg13g2_decap_8 FILLER_0_131_213 ();
 sg13g2_decap_8 FILLER_0_131_220 ();
 sg13g2_decap_8 FILLER_0_131_227 ();
 sg13g2_decap_8 FILLER_0_131_234 ();
 sg13g2_decap_8 FILLER_0_131_241 ();
 sg13g2_decap_8 FILLER_0_131_248 ();
 sg13g2_decap_8 FILLER_0_131_255 ();
 sg13g2_decap_8 FILLER_0_131_262 ();
 sg13g2_decap_8 FILLER_0_131_269 ();
 sg13g2_decap_8 FILLER_0_131_276 ();
 sg13g2_decap_8 FILLER_0_131_283 ();
 sg13g2_decap_8 FILLER_0_131_290 ();
 sg13g2_decap_8 FILLER_0_131_297 ();
 sg13g2_decap_8 FILLER_0_131_304 ();
 sg13g2_decap_8 FILLER_0_131_311 ();
 sg13g2_decap_8 FILLER_0_131_318 ();
 sg13g2_fill_1 FILLER_0_131_325 ();
 sg13g2_decap_4 FILLER_0_131_331 ();
 sg13g2_fill_1 FILLER_0_131_335 ();
 sg13g2_fill_1 FILLER_0_131_390 ();
 sg13g2_decap_8 FILLER_0_131_430 ();
 sg13g2_decap_8 FILLER_0_131_437 ();
 sg13g2_decap_8 FILLER_0_131_444 ();
 sg13g2_fill_1 FILLER_0_131_451 ();
 sg13g2_fill_2 FILLER_0_131_486 ();
 sg13g2_fill_1 FILLER_0_131_488 ();
 sg13g2_fill_2 FILLER_0_131_530 ();
 sg13g2_fill_1 FILLER_0_131_532 ();
 sg13g2_decap_4 FILLER_0_131_576 ();
 sg13g2_fill_2 FILLER_0_131_580 ();
 sg13g2_decap_8 FILLER_0_131_592 ();
 sg13g2_decap_8 FILLER_0_131_599 ();
 sg13g2_decap_8 FILLER_0_131_606 ();
 sg13g2_fill_1 FILLER_0_131_613 ();
 sg13g2_fill_1 FILLER_0_131_618 ();
 sg13g2_fill_2 FILLER_0_131_628 ();
 sg13g2_decap_8 FILLER_0_131_640 ();
 sg13g2_decap_8 FILLER_0_131_647 ();
 sg13g2_decap_8 FILLER_0_131_654 ();
 sg13g2_decap_8 FILLER_0_131_661 ();
 sg13g2_fill_2 FILLER_0_131_668 ();
 sg13g2_fill_1 FILLER_0_131_670 ();
 sg13g2_decap_8 FILLER_0_131_697 ();
 sg13g2_decap_8 FILLER_0_131_704 ();
 sg13g2_decap_8 FILLER_0_131_711 ();
 sg13g2_fill_1 FILLER_0_131_776 ();
 sg13g2_fill_1 FILLER_0_131_781 ();
 sg13g2_fill_1 FILLER_0_131_786 ();
 sg13g2_fill_1 FILLER_0_131_800 ();
 sg13g2_fill_2 FILLER_0_131_811 ();
 sg13g2_fill_1 FILLER_0_131_817 ();
 sg13g2_fill_1 FILLER_0_131_832 ();
 sg13g2_decap_4 FILLER_0_131_845 ();
 sg13g2_fill_1 FILLER_0_131_849 ();
 sg13g2_fill_2 FILLER_0_131_855 ();
 sg13g2_fill_1 FILLER_0_131_857 ();
 sg13g2_fill_1 FILLER_0_131_872 ();
 sg13g2_fill_2 FILLER_0_131_890 ();
 sg13g2_fill_2 FILLER_0_131_953 ();
 sg13g2_fill_1 FILLER_0_131_955 ();
 sg13g2_fill_2 FILLER_0_131_970 ();
 sg13g2_fill_1 FILLER_0_131_976 ();
 sg13g2_fill_1 FILLER_0_131_981 ();
 sg13g2_fill_1 FILLER_0_131_987 ();
 sg13g2_fill_1 FILLER_0_131_998 ();
 sg13g2_fill_2 FILLER_0_131_1014 ();
 sg13g2_fill_2 FILLER_0_131_1020 ();
 sg13g2_fill_1 FILLER_0_131_1022 ();
 sg13g2_decap_8 FILLER_0_131_1038 ();
 sg13g2_fill_1 FILLER_0_131_1045 ();
 sg13g2_fill_2 FILLER_0_131_1059 ();
 sg13g2_decap_8 FILLER_0_131_1065 ();
 sg13g2_decap_8 FILLER_0_131_1072 ();
 sg13g2_fill_1 FILLER_0_131_1079 ();
 sg13g2_decap_8 FILLER_0_131_1114 ();
 sg13g2_decap_8 FILLER_0_131_1121 ();
 sg13g2_decap_8 FILLER_0_131_1128 ();
 sg13g2_decap_8 FILLER_0_131_1135 ();
 sg13g2_decap_8 FILLER_0_131_1142 ();
 sg13g2_decap_8 FILLER_0_131_1149 ();
 sg13g2_decap_8 FILLER_0_131_1156 ();
 sg13g2_decap_8 FILLER_0_131_1163 ();
 sg13g2_decap_8 FILLER_0_131_1170 ();
 sg13g2_decap_8 FILLER_0_131_1177 ();
 sg13g2_decap_8 FILLER_0_131_1184 ();
 sg13g2_decap_8 FILLER_0_131_1191 ();
 sg13g2_decap_8 FILLER_0_131_1198 ();
 sg13g2_decap_8 FILLER_0_131_1205 ();
 sg13g2_decap_8 FILLER_0_131_1212 ();
 sg13g2_decap_8 FILLER_0_131_1219 ();
 sg13g2_fill_2 FILLER_0_131_1226 ();
 sg13g2_decap_8 FILLER_0_132_0 ();
 sg13g2_decap_8 FILLER_0_132_7 ();
 sg13g2_decap_8 FILLER_0_132_14 ();
 sg13g2_decap_8 FILLER_0_132_21 ();
 sg13g2_decap_8 FILLER_0_132_28 ();
 sg13g2_decap_8 FILLER_0_132_35 ();
 sg13g2_fill_2 FILLER_0_132_42 ();
 sg13g2_fill_1 FILLER_0_132_44 ();
 sg13g2_fill_1 FILLER_0_132_55 ();
 sg13g2_fill_1 FILLER_0_132_82 ();
 sg13g2_fill_1 FILLER_0_132_93 ();
 sg13g2_decap_8 FILLER_0_132_142 ();
 sg13g2_decap_8 FILLER_0_132_149 ();
 sg13g2_fill_2 FILLER_0_132_156 ();
 sg13g2_fill_1 FILLER_0_132_158 ();
 sg13g2_decap_8 FILLER_0_132_208 ();
 sg13g2_decap_8 FILLER_0_132_220 ();
 sg13g2_decap_8 FILLER_0_132_227 ();
 sg13g2_decap_8 FILLER_0_132_234 ();
 sg13g2_decap_8 FILLER_0_132_241 ();
 sg13g2_decap_8 FILLER_0_132_248 ();
 sg13g2_decap_8 FILLER_0_132_255 ();
 sg13g2_decap_8 FILLER_0_132_262 ();
 sg13g2_decap_8 FILLER_0_132_269 ();
 sg13g2_decap_8 FILLER_0_132_276 ();
 sg13g2_decap_8 FILLER_0_132_283 ();
 sg13g2_decap_8 FILLER_0_132_290 ();
 sg13g2_decap_8 FILLER_0_132_297 ();
 sg13g2_decap_8 FILLER_0_132_304 ();
 sg13g2_decap_4 FILLER_0_132_311 ();
 sg13g2_fill_1 FILLER_0_132_315 ();
 sg13g2_decap_4 FILLER_0_132_320 ();
 sg13g2_decap_8 FILLER_0_132_354 ();
 sg13g2_decap_8 FILLER_0_132_361 ();
 sg13g2_fill_2 FILLER_0_132_368 ();
 sg13g2_fill_1 FILLER_0_132_374 ();
 sg13g2_fill_1 FILLER_0_132_385 ();
 sg13g2_fill_1 FILLER_0_132_396 ();
 sg13g2_fill_1 FILLER_0_132_401 ();
 sg13g2_fill_1 FILLER_0_132_412 ();
 sg13g2_decap_8 FILLER_0_132_416 ();
 sg13g2_decap_8 FILLER_0_132_423 ();
 sg13g2_decap_8 FILLER_0_132_430 ();
 sg13g2_decap_8 FILLER_0_132_437 ();
 sg13g2_decap_8 FILLER_0_132_444 ();
 sg13g2_decap_8 FILLER_0_132_451 ();
 sg13g2_fill_1 FILLER_0_132_499 ();
 sg13g2_decap_8 FILLER_0_132_504 ();
 sg13g2_decap_4 FILLER_0_132_511 ();
 sg13g2_fill_1 FILLER_0_132_515 ();
 sg13g2_decap_4 FILLER_0_132_526 ();
 sg13g2_fill_2 FILLER_0_132_535 ();
 sg13g2_fill_2 FILLER_0_132_541 ();
 sg13g2_fill_1 FILLER_0_132_543 ();
 sg13g2_decap_8 FILLER_0_132_554 ();
 sg13g2_decap_8 FILLER_0_132_561 ();
 sg13g2_decap_8 FILLER_0_132_568 ();
 sg13g2_decap_8 FILLER_0_132_575 ();
 sg13g2_decap_8 FILLER_0_132_582 ();
 sg13g2_decap_8 FILLER_0_132_589 ();
 sg13g2_decap_8 FILLER_0_132_596 ();
 sg13g2_decap_8 FILLER_0_132_603 ();
 sg13g2_decap_8 FILLER_0_132_610 ();
 sg13g2_decap_8 FILLER_0_132_617 ();
 sg13g2_decap_8 FILLER_0_132_665 ();
 sg13g2_decap_4 FILLER_0_132_672 ();
 sg13g2_fill_1 FILLER_0_132_676 ();
 sg13g2_decap_8 FILLER_0_132_711 ();
 sg13g2_fill_1 FILLER_0_132_718 ();
 sg13g2_fill_1 FILLER_0_132_742 ();
 sg13g2_decap_4 FILLER_0_132_747 ();
 sg13g2_fill_1 FILLER_0_132_751 ();
 sg13g2_fill_1 FILLER_0_132_772 ();
 sg13g2_fill_2 FILLER_0_132_781 ();
 sg13g2_fill_2 FILLER_0_132_805 ();
 sg13g2_fill_1 FILLER_0_132_807 ();
 sg13g2_fill_1 FILLER_0_132_811 ();
 sg13g2_fill_1 FILLER_0_132_829 ();
 sg13g2_fill_2 FILLER_0_132_844 ();
 sg13g2_fill_1 FILLER_0_132_846 ();
 sg13g2_fill_1 FILLER_0_132_856 ();
 sg13g2_decap_4 FILLER_0_132_862 ();
 sg13g2_fill_1 FILLER_0_132_866 ();
 sg13g2_fill_1 FILLER_0_132_885 ();
 sg13g2_fill_2 FILLER_0_132_898 ();
 sg13g2_fill_1 FILLER_0_132_905 ();
 sg13g2_fill_1 FILLER_0_132_941 ();
 sg13g2_fill_2 FILLER_0_132_951 ();
 sg13g2_fill_1 FILLER_0_132_953 ();
 sg13g2_fill_1 FILLER_0_132_958 ();
 sg13g2_fill_1 FILLER_0_132_968 ();
 sg13g2_decap_8 FILLER_0_132_978 ();
 sg13g2_decap_8 FILLER_0_132_985 ();
 sg13g2_decap_8 FILLER_0_132_992 ();
 sg13g2_decap_8 FILLER_0_132_999 ();
 sg13g2_decap_8 FILLER_0_132_1006 ();
 sg13g2_decap_8 FILLER_0_132_1013 ();
 sg13g2_decap_4 FILLER_0_132_1020 ();
 sg13g2_fill_1 FILLER_0_132_1024 ();
 sg13g2_decap_8 FILLER_0_132_1065 ();
 sg13g2_decap_8 FILLER_0_132_1072 ();
 sg13g2_fill_2 FILLER_0_132_1079 ();
 sg13g2_fill_1 FILLER_0_132_1086 ();
 sg13g2_decap_8 FILLER_0_132_1101 ();
 sg13g2_decap_8 FILLER_0_132_1108 ();
 sg13g2_decap_8 FILLER_0_132_1115 ();
 sg13g2_decap_8 FILLER_0_132_1122 ();
 sg13g2_decap_8 FILLER_0_132_1129 ();
 sg13g2_decap_8 FILLER_0_132_1136 ();
 sg13g2_decap_8 FILLER_0_132_1143 ();
 sg13g2_decap_8 FILLER_0_132_1150 ();
 sg13g2_decap_8 FILLER_0_132_1157 ();
 sg13g2_decap_8 FILLER_0_132_1164 ();
 sg13g2_decap_8 FILLER_0_132_1171 ();
 sg13g2_decap_8 FILLER_0_132_1178 ();
 sg13g2_decap_8 FILLER_0_132_1185 ();
 sg13g2_decap_8 FILLER_0_132_1192 ();
 sg13g2_decap_8 FILLER_0_132_1199 ();
 sg13g2_decap_8 FILLER_0_132_1206 ();
 sg13g2_decap_8 FILLER_0_132_1213 ();
 sg13g2_decap_8 FILLER_0_132_1220 ();
 sg13g2_fill_1 FILLER_0_132_1227 ();
 sg13g2_decap_8 FILLER_0_133_0 ();
 sg13g2_decap_8 FILLER_0_133_7 ();
 sg13g2_decap_8 FILLER_0_133_14 ();
 sg13g2_decap_8 FILLER_0_133_21 ();
 sg13g2_decap_8 FILLER_0_133_28 ();
 sg13g2_decap_8 FILLER_0_133_35 ();
 sg13g2_decap_8 FILLER_0_133_42 ();
 sg13g2_decap_8 FILLER_0_133_135 ();
 sg13g2_decap_8 FILLER_0_133_147 ();
 sg13g2_decap_8 FILLER_0_133_154 ();
 sg13g2_fill_2 FILLER_0_133_161 ();
 sg13g2_fill_1 FILLER_0_133_163 ();
 sg13g2_fill_1 FILLER_0_133_176 ();
 sg13g2_decap_4 FILLER_0_133_203 ();
 sg13g2_fill_2 FILLER_0_133_207 ();
 sg13g2_decap_4 FILLER_0_133_245 ();
 sg13g2_fill_2 FILLER_0_133_249 ();
 sg13g2_decap_8 FILLER_0_133_255 ();
 sg13g2_decap_8 FILLER_0_133_262 ();
 sg13g2_decap_8 FILLER_0_133_269 ();
 sg13g2_decap_8 FILLER_0_133_276 ();
 sg13g2_decap_8 FILLER_0_133_283 ();
 sg13g2_decap_8 FILLER_0_133_290 ();
 sg13g2_decap_8 FILLER_0_133_297 ();
 sg13g2_decap_8 FILLER_0_133_304 ();
 sg13g2_fill_2 FILLER_0_133_311 ();
 sg13g2_decap_8 FILLER_0_133_354 ();
 sg13g2_decap_8 FILLER_0_133_361 ();
 sg13g2_decap_8 FILLER_0_133_368 ();
 sg13g2_decap_8 FILLER_0_133_375 ();
 sg13g2_decap_8 FILLER_0_133_382 ();
 sg13g2_decap_8 FILLER_0_133_389 ();
 sg13g2_decap_8 FILLER_0_133_396 ();
 sg13g2_decap_8 FILLER_0_133_413 ();
 sg13g2_decap_8 FILLER_0_133_420 ();
 sg13g2_decap_8 FILLER_0_133_427 ();
 sg13g2_decap_8 FILLER_0_133_434 ();
 sg13g2_decap_8 FILLER_0_133_441 ();
 sg13g2_decap_8 FILLER_0_133_448 ();
 sg13g2_decap_8 FILLER_0_133_455 ();
 sg13g2_decap_4 FILLER_0_133_467 ();
 sg13g2_decap_4 FILLER_0_133_475 ();
 sg13g2_decap_8 FILLER_0_133_489 ();
 sg13g2_fill_2 FILLER_0_133_527 ();
 sg13g2_decap_4 FILLER_0_133_539 ();
 sg13g2_decap_8 FILLER_0_133_553 ();
 sg13g2_decap_8 FILLER_0_133_560 ();
 sg13g2_decap_8 FILLER_0_133_567 ();
 sg13g2_decap_8 FILLER_0_133_574 ();
 sg13g2_decap_8 FILLER_0_133_581 ();
 sg13g2_decap_8 FILLER_0_133_588 ();
 sg13g2_decap_8 FILLER_0_133_595 ();
 sg13g2_decap_8 FILLER_0_133_602 ();
 sg13g2_decap_8 FILLER_0_133_609 ();
 sg13g2_decap_8 FILLER_0_133_616 ();
 sg13g2_decap_4 FILLER_0_133_623 ();
 sg13g2_fill_2 FILLER_0_133_627 ();
 sg13g2_fill_2 FILLER_0_133_659 ();
 sg13g2_decap_8 FILLER_0_133_669 ();
 sg13g2_decap_8 FILLER_0_133_676 ();
 sg13g2_fill_2 FILLER_0_133_683 ();
 sg13g2_decap_8 FILLER_0_133_708 ();
 sg13g2_decap_8 FILLER_0_133_715 ();
 sg13g2_decap_4 FILLER_0_133_722 ();
 sg13g2_decap_4 FILLER_0_133_744 ();
 sg13g2_fill_1 FILLER_0_133_748 ();
 sg13g2_fill_1 FILLER_0_133_753 ();
 sg13g2_fill_2 FILLER_0_133_759 ();
 sg13g2_fill_2 FILLER_0_133_785 ();
 sg13g2_fill_1 FILLER_0_133_787 ();
 sg13g2_fill_2 FILLER_0_133_833 ();
 sg13g2_fill_1 FILLER_0_133_835 ();
 sg13g2_fill_1 FILLER_0_133_860 ();
 sg13g2_fill_2 FILLER_0_133_867 ();
 sg13g2_fill_1 FILLER_0_133_869 ();
 sg13g2_fill_2 FILLER_0_133_878 ();
 sg13g2_decap_8 FILLER_0_133_911 ();
 sg13g2_fill_1 FILLER_0_133_924 ();
 sg13g2_fill_2 FILLER_0_133_934 ();
 sg13g2_fill_2 FILLER_0_133_944 ();
 sg13g2_fill_1 FILLER_0_133_951 ();
 sg13g2_fill_2 FILLER_0_133_972 ();
 sg13g2_fill_2 FILLER_0_133_984 ();
 sg13g2_decap_4 FILLER_0_133_990 ();
 sg13g2_decap_4 FILLER_0_133_999 ();
 sg13g2_fill_2 FILLER_0_133_1007 ();
 sg13g2_fill_1 FILLER_0_133_1009 ();
 sg13g2_decap_4 FILLER_0_133_1020 ();
 sg13g2_fill_2 FILLER_0_133_1024 ();
 sg13g2_fill_2 FILLER_0_133_1040 ();
 sg13g2_fill_1 FILLER_0_133_1042 ();
 sg13g2_fill_2 FILLER_0_133_1059 ();
 sg13g2_decap_8 FILLER_0_133_1065 ();
 sg13g2_decap_8 FILLER_0_133_1072 ();
 sg13g2_fill_2 FILLER_0_133_1079 ();
 sg13g2_fill_1 FILLER_0_133_1081 ();
 sg13g2_decap_8 FILLER_0_133_1108 ();
 sg13g2_decap_8 FILLER_0_133_1115 ();
 sg13g2_decap_8 FILLER_0_133_1122 ();
 sg13g2_decap_8 FILLER_0_133_1129 ();
 sg13g2_decap_8 FILLER_0_133_1136 ();
 sg13g2_decap_8 FILLER_0_133_1143 ();
 sg13g2_decap_8 FILLER_0_133_1150 ();
 sg13g2_decap_8 FILLER_0_133_1157 ();
 sg13g2_decap_8 FILLER_0_133_1164 ();
 sg13g2_decap_8 FILLER_0_133_1171 ();
 sg13g2_decap_8 FILLER_0_133_1178 ();
 sg13g2_decap_8 FILLER_0_133_1185 ();
 sg13g2_decap_8 FILLER_0_133_1192 ();
 sg13g2_decap_8 FILLER_0_133_1199 ();
 sg13g2_decap_8 FILLER_0_133_1206 ();
 sg13g2_decap_8 FILLER_0_133_1213 ();
 sg13g2_decap_8 FILLER_0_133_1220 ();
 sg13g2_fill_1 FILLER_0_133_1227 ();
 sg13g2_decap_8 FILLER_0_134_0 ();
 sg13g2_decap_8 FILLER_0_134_7 ();
 sg13g2_decap_8 FILLER_0_134_14 ();
 sg13g2_decap_8 FILLER_0_134_21 ();
 sg13g2_decap_8 FILLER_0_134_28 ();
 sg13g2_decap_4 FILLER_0_134_35 ();
 sg13g2_fill_2 FILLER_0_134_39 ();
 sg13g2_fill_1 FILLER_0_134_56 ();
 sg13g2_fill_1 FILLER_0_134_62 ();
 sg13g2_fill_1 FILLER_0_134_67 ();
 sg13g2_fill_2 FILLER_0_134_78 ();
 sg13g2_fill_1 FILLER_0_134_98 ();
 sg13g2_decap_8 FILLER_0_134_103 ();
 sg13g2_decap_8 FILLER_0_134_110 ();
 sg13g2_decap_8 FILLER_0_134_117 ();
 sg13g2_decap_8 FILLER_0_134_159 ();
 sg13g2_decap_8 FILLER_0_134_166 ();
 sg13g2_fill_2 FILLER_0_134_173 ();
 sg13g2_decap_8 FILLER_0_134_184 ();
 sg13g2_fill_1 FILLER_0_134_191 ();
 sg13g2_fill_1 FILLER_0_134_197 ();
 sg13g2_decap_8 FILLER_0_134_208 ();
 sg13g2_fill_1 FILLER_0_134_215 ();
 sg13g2_decap_8 FILLER_0_134_255 ();
 sg13g2_decap_8 FILLER_0_134_262 ();
 sg13g2_decap_8 FILLER_0_134_269 ();
 sg13g2_decap_8 FILLER_0_134_276 ();
 sg13g2_decap_8 FILLER_0_134_283 ();
 sg13g2_decap_8 FILLER_0_134_290 ();
 sg13g2_decap_8 FILLER_0_134_297 ();
 sg13g2_decap_8 FILLER_0_134_304 ();
 sg13g2_decap_4 FILLER_0_134_311 ();
 sg13g2_fill_1 FILLER_0_134_315 ();
 sg13g2_decap_8 FILLER_0_134_345 ();
 sg13g2_decap_8 FILLER_0_134_352 ();
 sg13g2_fill_2 FILLER_0_134_359 ();
 sg13g2_decap_8 FILLER_0_134_365 ();
 sg13g2_fill_2 FILLER_0_134_372 ();
 sg13g2_fill_1 FILLER_0_134_374 ();
 sg13g2_decap_8 FILLER_0_134_395 ();
 sg13g2_fill_1 FILLER_0_134_402 ();
 sg13g2_decap_8 FILLER_0_134_434 ();
 sg13g2_decap_4 FILLER_0_134_441 ();
 sg13g2_decap_4 FILLER_0_134_455 ();
 sg13g2_decap_8 FILLER_0_134_489 ();
 sg13g2_decap_4 FILLER_0_134_496 ();
 sg13g2_fill_2 FILLER_0_134_536 ();
 sg13g2_fill_1 FILLER_0_134_538 ();
 sg13g2_decap_8 FILLER_0_134_565 ();
 sg13g2_decap_8 FILLER_0_134_572 ();
 sg13g2_decap_8 FILLER_0_134_579 ();
 sg13g2_decap_8 FILLER_0_134_586 ();
 sg13g2_decap_8 FILLER_0_134_593 ();
 sg13g2_decap_8 FILLER_0_134_600 ();
 sg13g2_decap_8 FILLER_0_134_607 ();
 sg13g2_decap_8 FILLER_0_134_614 ();
 sg13g2_decap_8 FILLER_0_134_621 ();
 sg13g2_decap_8 FILLER_0_134_628 ();
 sg13g2_decap_4 FILLER_0_134_635 ();
 sg13g2_fill_1 FILLER_0_134_643 ();
 sg13g2_decap_4 FILLER_0_134_679 ();
 sg13g2_fill_2 FILLER_0_134_709 ();
 sg13g2_fill_1 FILLER_0_134_772 ();
 sg13g2_fill_1 FILLER_0_134_778 ();
 sg13g2_fill_1 FILLER_0_134_783 ();
 sg13g2_fill_2 FILLER_0_134_792 ();
 sg13g2_fill_1 FILLER_0_134_815 ();
 sg13g2_decap_8 FILLER_0_134_831 ();
 sg13g2_decap_4 FILLER_0_134_838 ();
 sg13g2_fill_1 FILLER_0_134_842 ();
 sg13g2_fill_1 FILLER_0_134_849 ();
 sg13g2_fill_2 FILLER_0_134_854 ();
 sg13g2_decap_8 FILLER_0_134_861 ();
 sg13g2_decap_4 FILLER_0_134_868 ();
 sg13g2_decap_4 FILLER_0_134_877 ();
 sg13g2_fill_1 FILLER_0_134_881 ();
 sg13g2_decap_8 FILLER_0_134_927 ();
 sg13g2_decap_8 FILLER_0_134_934 ();
 sg13g2_fill_2 FILLER_0_134_941 ();
 sg13g2_fill_2 FILLER_0_134_947 ();
 sg13g2_fill_1 FILLER_0_134_949 ();
 sg13g2_fill_2 FILLER_0_134_954 ();
 sg13g2_fill_1 FILLER_0_134_956 ();
 sg13g2_fill_1 FILLER_0_134_987 ();
 sg13g2_fill_2 FILLER_0_134_1018 ();
 sg13g2_fill_1 FILLER_0_134_1020 ();
 sg13g2_fill_1 FILLER_0_134_1025 ();
 sg13g2_decap_8 FILLER_0_134_1034 ();
 sg13g2_decap_4 FILLER_0_134_1041 ();
 sg13g2_fill_1 FILLER_0_134_1045 ();
 sg13g2_decap_8 FILLER_0_134_1073 ();
 sg13g2_fill_1 FILLER_0_134_1080 ();
 sg13g2_decap_8 FILLER_0_134_1112 ();
 sg13g2_decap_8 FILLER_0_134_1119 ();
 sg13g2_decap_8 FILLER_0_134_1126 ();
 sg13g2_decap_8 FILLER_0_134_1133 ();
 sg13g2_decap_8 FILLER_0_134_1140 ();
 sg13g2_decap_8 FILLER_0_134_1147 ();
 sg13g2_decap_8 FILLER_0_134_1154 ();
 sg13g2_decap_8 FILLER_0_134_1161 ();
 sg13g2_decap_8 FILLER_0_134_1168 ();
 sg13g2_decap_8 FILLER_0_134_1175 ();
 sg13g2_decap_8 FILLER_0_134_1182 ();
 sg13g2_decap_8 FILLER_0_134_1189 ();
 sg13g2_decap_8 FILLER_0_134_1196 ();
 sg13g2_decap_8 FILLER_0_134_1203 ();
 sg13g2_decap_8 FILLER_0_134_1210 ();
 sg13g2_decap_8 FILLER_0_134_1217 ();
 sg13g2_decap_4 FILLER_0_134_1224 ();
 sg13g2_decap_8 FILLER_0_135_0 ();
 sg13g2_decap_8 FILLER_0_135_7 ();
 sg13g2_decap_8 FILLER_0_135_14 ();
 sg13g2_decap_8 FILLER_0_135_21 ();
 sg13g2_decap_4 FILLER_0_135_28 ();
 sg13g2_fill_1 FILLER_0_135_32 ();
 sg13g2_decap_8 FILLER_0_135_75 ();
 sg13g2_decap_8 FILLER_0_135_82 ();
 sg13g2_decap_8 FILLER_0_135_89 ();
 sg13g2_decap_8 FILLER_0_135_96 ();
 sg13g2_decap_8 FILLER_0_135_103 ();
 sg13g2_decap_8 FILLER_0_135_110 ();
 sg13g2_fill_2 FILLER_0_135_132 ();
 sg13g2_fill_1 FILLER_0_135_134 ();
 sg13g2_decap_4 FILLER_0_135_171 ();
 sg13g2_decap_4 FILLER_0_135_221 ();
 sg13g2_fill_1 FILLER_0_135_230 ();
 sg13g2_decap_8 FILLER_0_135_261 ();
 sg13g2_decap_8 FILLER_0_135_268 ();
 sg13g2_decap_8 FILLER_0_135_275 ();
 sg13g2_decap_8 FILLER_0_135_282 ();
 sg13g2_decap_8 FILLER_0_135_289 ();
 sg13g2_decap_8 FILLER_0_135_296 ();
 sg13g2_decap_8 FILLER_0_135_303 ();
 sg13g2_decap_4 FILLER_0_135_310 ();
 sg13g2_decap_8 FILLER_0_135_345 ();
 sg13g2_decap_4 FILLER_0_135_352 ();
 sg13g2_fill_1 FILLER_0_135_356 ();
 sg13g2_fill_1 FILLER_0_135_383 ();
 sg13g2_fill_2 FILLER_0_135_389 ();
 sg13g2_fill_1 FILLER_0_135_391 ();
 sg13g2_decap_4 FILLER_0_135_422 ();
 sg13g2_fill_1 FILLER_0_135_426 ();
 sg13g2_decap_4 FILLER_0_135_458 ();
 sg13g2_fill_1 FILLER_0_135_462 ();
 sg13g2_decap_4 FILLER_0_135_468 ();
 sg13g2_fill_2 FILLER_0_135_472 ();
 sg13g2_decap_4 FILLER_0_135_478 ();
 sg13g2_fill_2 FILLER_0_135_482 ();
 sg13g2_fill_2 FILLER_0_135_494 ();
 sg13g2_decap_8 FILLER_0_135_561 ();
 sg13g2_decap_8 FILLER_0_135_568 ();
 sg13g2_decap_8 FILLER_0_135_575 ();
 sg13g2_decap_8 FILLER_0_135_582 ();
 sg13g2_decap_8 FILLER_0_135_589 ();
 sg13g2_decap_8 FILLER_0_135_596 ();
 sg13g2_decap_8 FILLER_0_135_603 ();
 sg13g2_decap_8 FILLER_0_135_610 ();
 sg13g2_decap_8 FILLER_0_135_617 ();
 sg13g2_decap_8 FILLER_0_135_624 ();
 sg13g2_decap_8 FILLER_0_135_631 ();
 sg13g2_decap_4 FILLER_0_135_638 ();
 sg13g2_fill_1 FILLER_0_135_688 ();
 sg13g2_fill_2 FILLER_0_135_707 ();
 sg13g2_fill_1 FILLER_0_135_709 ();
 sg13g2_fill_1 FILLER_0_135_743 ();
 sg13g2_fill_2 FILLER_0_135_767 ();
 sg13g2_fill_1 FILLER_0_135_769 ();
 sg13g2_fill_2 FILLER_0_135_775 ();
 sg13g2_decap_4 FILLER_0_135_781 ();
 sg13g2_fill_2 FILLER_0_135_785 ();
 sg13g2_decap_4 FILLER_0_135_795 ();
 sg13g2_fill_1 FILLER_0_135_799 ();
 sg13g2_fill_1 FILLER_0_135_825 ();
 sg13g2_decap_8 FILLER_0_135_831 ();
 sg13g2_decap_8 FILLER_0_135_838 ();
 sg13g2_decap_4 FILLER_0_135_845 ();
 sg13g2_fill_2 FILLER_0_135_849 ();
 sg13g2_fill_1 FILLER_0_135_859 ();
 sg13g2_decap_8 FILLER_0_135_865 ();
 sg13g2_fill_1 FILLER_0_135_872 ();
 sg13g2_decap_4 FILLER_0_135_878 ();
 sg13g2_fill_1 FILLER_0_135_882 ();
 sg13g2_decap_4 FILLER_0_135_888 ();
 sg13g2_fill_2 FILLER_0_135_907 ();
 sg13g2_fill_1 FILLER_0_135_909 ();
 sg13g2_fill_1 FILLER_0_135_922 ();
 sg13g2_fill_2 FILLER_0_135_932 ();
 sg13g2_decap_4 FILLER_0_135_938 ();
 sg13g2_decap_8 FILLER_0_135_957 ();
 sg13g2_fill_2 FILLER_0_135_964 ();
 sg13g2_decap_8 FILLER_0_135_979 ();
 sg13g2_fill_1 FILLER_0_135_986 ();
 sg13g2_fill_2 FILLER_0_135_992 ();
 sg13g2_fill_1 FILLER_0_135_994 ();
 sg13g2_fill_2 FILLER_0_135_999 ();
 sg13g2_decap_8 FILLER_0_135_1031 ();
 sg13g2_fill_2 FILLER_0_135_1038 ();
 sg13g2_fill_1 FILLER_0_135_1040 ();
 sg13g2_fill_1 FILLER_0_135_1046 ();
 sg13g2_fill_2 FILLER_0_135_1060 ();
 sg13g2_decap_8 FILLER_0_135_1072 ();
 sg13g2_decap_8 FILLER_0_135_1079 ();
 sg13g2_decap_4 FILLER_0_135_1086 ();
 sg13g2_decap_8 FILLER_0_135_1104 ();
 sg13g2_decap_8 FILLER_0_135_1111 ();
 sg13g2_decap_8 FILLER_0_135_1118 ();
 sg13g2_decap_8 FILLER_0_135_1125 ();
 sg13g2_decap_8 FILLER_0_135_1132 ();
 sg13g2_decap_8 FILLER_0_135_1139 ();
 sg13g2_decap_8 FILLER_0_135_1146 ();
 sg13g2_decap_8 FILLER_0_135_1153 ();
 sg13g2_decap_8 FILLER_0_135_1160 ();
 sg13g2_decap_8 FILLER_0_135_1167 ();
 sg13g2_decap_8 FILLER_0_135_1174 ();
 sg13g2_decap_8 FILLER_0_135_1181 ();
 sg13g2_decap_8 FILLER_0_135_1188 ();
 sg13g2_decap_8 FILLER_0_135_1195 ();
 sg13g2_decap_8 FILLER_0_135_1202 ();
 sg13g2_decap_8 FILLER_0_135_1209 ();
 sg13g2_decap_8 FILLER_0_135_1216 ();
 sg13g2_decap_4 FILLER_0_135_1223 ();
 sg13g2_fill_1 FILLER_0_135_1227 ();
 sg13g2_decap_8 FILLER_0_136_0 ();
 sg13g2_decap_8 FILLER_0_136_7 ();
 sg13g2_decap_8 FILLER_0_136_14 ();
 sg13g2_decap_8 FILLER_0_136_21 ();
 sg13g2_fill_2 FILLER_0_136_61 ();
 sg13g2_decap_8 FILLER_0_136_78 ();
 sg13g2_decap_8 FILLER_0_136_85 ();
 sg13g2_decap_8 FILLER_0_136_92 ();
 sg13g2_fill_2 FILLER_0_136_99 ();
 sg13g2_fill_2 FILLER_0_136_109 ();
 sg13g2_fill_1 FILLER_0_136_111 ();
 sg13g2_decap_4 FILLER_0_136_117 ();
 sg13g2_fill_2 FILLER_0_136_147 ();
 sg13g2_fill_1 FILLER_0_136_149 ();
 sg13g2_fill_2 FILLER_0_136_164 ();
 sg13g2_fill_1 FILLER_0_136_166 ();
 sg13g2_fill_2 FILLER_0_136_193 ();
 sg13g2_fill_1 FILLER_0_136_195 ();
 sg13g2_decap_8 FILLER_0_136_200 ();
 sg13g2_decap_4 FILLER_0_136_207 ();
 sg13g2_fill_1 FILLER_0_136_211 ();
 sg13g2_decap_8 FILLER_0_136_222 ();
 sg13g2_decap_4 FILLER_0_136_229 ();
 sg13g2_fill_1 FILLER_0_136_233 ();
 sg13g2_decap_8 FILLER_0_136_251 ();
 sg13g2_decap_8 FILLER_0_136_258 ();
 sg13g2_decap_8 FILLER_0_136_265 ();
 sg13g2_decap_8 FILLER_0_136_272 ();
 sg13g2_decap_8 FILLER_0_136_279 ();
 sg13g2_decap_8 FILLER_0_136_286 ();
 sg13g2_decap_8 FILLER_0_136_293 ();
 sg13g2_decap_8 FILLER_0_136_300 ();
 sg13g2_decap_8 FILLER_0_136_307 ();
 sg13g2_decap_4 FILLER_0_136_314 ();
 sg13g2_fill_1 FILLER_0_136_349 ();
 sg13g2_fill_2 FILLER_0_136_388 ();
 sg13g2_fill_1 FILLER_0_136_390 ();
 sg13g2_fill_2 FILLER_0_136_405 ();
 sg13g2_decap_8 FILLER_0_136_417 ();
 sg13g2_decap_4 FILLER_0_136_459 ();
 sg13g2_fill_2 FILLER_0_136_463 ();
 sg13g2_decap_8 FILLER_0_136_491 ();
 sg13g2_decap_8 FILLER_0_136_498 ();
 sg13g2_decap_4 FILLER_0_136_505 ();
 sg13g2_decap_8 FILLER_0_136_550 ();
 sg13g2_decap_8 FILLER_0_136_557 ();
 sg13g2_decap_8 FILLER_0_136_564 ();
 sg13g2_decap_8 FILLER_0_136_571 ();
 sg13g2_decap_8 FILLER_0_136_578 ();
 sg13g2_decap_8 FILLER_0_136_585 ();
 sg13g2_decap_8 FILLER_0_136_592 ();
 sg13g2_decap_8 FILLER_0_136_599 ();
 sg13g2_decap_8 FILLER_0_136_606 ();
 sg13g2_decap_8 FILLER_0_136_613 ();
 sg13g2_decap_8 FILLER_0_136_620 ();
 sg13g2_decap_8 FILLER_0_136_627 ();
 sg13g2_decap_8 FILLER_0_136_634 ();
 sg13g2_decap_8 FILLER_0_136_641 ();
 sg13g2_fill_2 FILLER_0_136_648 ();
 sg13g2_fill_1 FILLER_0_136_680 ();
 sg13g2_decap_8 FILLER_0_136_712 ();
 sg13g2_fill_2 FILLER_0_136_758 ();
 sg13g2_decap_8 FILLER_0_136_795 ();
 sg13g2_decap_8 FILLER_0_136_802 ();
 sg13g2_decap_8 FILLER_0_136_809 ();
 sg13g2_fill_1 FILLER_0_136_816 ();
 sg13g2_decap_8 FILLER_0_136_836 ();
 sg13g2_fill_1 FILLER_0_136_843 ();
 sg13g2_fill_1 FILLER_0_136_849 ();
 sg13g2_fill_2 FILLER_0_136_860 ();
 sg13g2_fill_1 FILLER_0_136_862 ();
 sg13g2_decap_4 FILLER_0_136_871 ();
 sg13g2_fill_1 FILLER_0_136_875 ();
 sg13g2_fill_2 FILLER_0_136_897 ();
 sg13g2_fill_1 FILLER_0_136_899 ();
 sg13g2_fill_1 FILLER_0_136_905 ();
 sg13g2_decap_8 FILLER_0_136_944 ();
 sg13g2_decap_8 FILLER_0_136_951 ();
 sg13g2_fill_1 FILLER_0_136_958 ();
 sg13g2_decap_8 FILLER_0_136_963 ();
 sg13g2_decap_8 FILLER_0_136_970 ();
 sg13g2_fill_1 FILLER_0_136_977 ();
 sg13g2_fill_2 FILLER_0_136_982 ();
 sg13g2_fill_2 FILLER_0_136_988 ();
 sg13g2_decap_8 FILLER_0_136_995 ();
 sg13g2_fill_2 FILLER_0_136_1002 ();
 sg13g2_fill_1 FILLER_0_136_1004 ();
 sg13g2_fill_1 FILLER_0_136_1017 ();
 sg13g2_decap_4 FILLER_0_136_1031 ();
 sg13g2_fill_2 FILLER_0_136_1053 ();
 sg13g2_fill_1 FILLER_0_136_1055 ();
 sg13g2_decap_8 FILLER_0_136_1086 ();
 sg13g2_decap_8 FILLER_0_136_1093 ();
 sg13g2_decap_8 FILLER_0_136_1100 ();
 sg13g2_decap_8 FILLER_0_136_1107 ();
 sg13g2_decap_8 FILLER_0_136_1114 ();
 sg13g2_decap_8 FILLER_0_136_1121 ();
 sg13g2_decap_8 FILLER_0_136_1128 ();
 sg13g2_decap_8 FILLER_0_136_1135 ();
 sg13g2_decap_8 FILLER_0_136_1142 ();
 sg13g2_decap_8 FILLER_0_136_1149 ();
 sg13g2_decap_8 FILLER_0_136_1156 ();
 sg13g2_decap_8 FILLER_0_136_1163 ();
 sg13g2_decap_8 FILLER_0_136_1170 ();
 sg13g2_decap_8 FILLER_0_136_1177 ();
 sg13g2_decap_8 FILLER_0_136_1184 ();
 sg13g2_decap_8 FILLER_0_136_1191 ();
 sg13g2_decap_8 FILLER_0_136_1198 ();
 sg13g2_decap_8 FILLER_0_136_1205 ();
 sg13g2_decap_8 FILLER_0_136_1212 ();
 sg13g2_decap_8 FILLER_0_136_1219 ();
 sg13g2_fill_2 FILLER_0_136_1226 ();
 sg13g2_decap_8 FILLER_0_137_0 ();
 sg13g2_decap_8 FILLER_0_137_7 ();
 sg13g2_decap_8 FILLER_0_137_14 ();
 sg13g2_decap_8 FILLER_0_137_21 ();
 sg13g2_decap_8 FILLER_0_137_28 ();
 sg13g2_fill_2 FILLER_0_137_35 ();
 sg13g2_fill_1 FILLER_0_137_105 ();
 sg13g2_decap_8 FILLER_0_137_142 ();
 sg13g2_fill_2 FILLER_0_137_149 ();
 sg13g2_fill_1 FILLER_0_137_151 ();
 sg13g2_fill_2 FILLER_0_137_171 ();
 sg13g2_fill_1 FILLER_0_137_173 ();
 sg13g2_fill_2 FILLER_0_137_178 ();
 sg13g2_fill_1 FILLER_0_137_180 ();
 sg13g2_fill_2 FILLER_0_137_202 ();
 sg13g2_fill_1 FILLER_0_137_204 ();
 sg13g2_decap_8 FILLER_0_137_250 ();
 sg13g2_decap_8 FILLER_0_137_257 ();
 sg13g2_decap_8 FILLER_0_137_264 ();
 sg13g2_decap_8 FILLER_0_137_271 ();
 sg13g2_decap_8 FILLER_0_137_278 ();
 sg13g2_decap_8 FILLER_0_137_285 ();
 sg13g2_decap_8 FILLER_0_137_292 ();
 sg13g2_decap_8 FILLER_0_137_299 ();
 sg13g2_decap_8 FILLER_0_137_306 ();
 sg13g2_decap_8 FILLER_0_137_313 ();
 sg13g2_decap_4 FILLER_0_137_320 ();
 sg13g2_fill_1 FILLER_0_137_324 ();
 sg13g2_decap_8 FILLER_0_137_329 ();
 sg13g2_decap_4 FILLER_0_137_346 ();
 sg13g2_fill_2 FILLER_0_137_350 ();
 sg13g2_decap_8 FILLER_0_137_360 ();
 sg13g2_fill_2 FILLER_0_137_367 ();
 sg13g2_decap_8 FILLER_0_137_383 ();
 sg13g2_decap_8 FILLER_0_137_390 ();
 sg13g2_decap_8 FILLER_0_137_397 ();
 sg13g2_decap_8 FILLER_0_137_404 ();
 sg13g2_decap_8 FILLER_0_137_411 ();
 sg13g2_decap_8 FILLER_0_137_418 ();
 sg13g2_decap_8 FILLER_0_137_425 ();
 sg13g2_decap_8 FILLER_0_137_436 ();
 sg13g2_decap_8 FILLER_0_137_443 ();
 sg13g2_fill_1 FILLER_0_137_450 ();
 sg13g2_decap_8 FILLER_0_137_461 ();
 sg13g2_decap_4 FILLER_0_137_468 ();
 sg13g2_fill_1 FILLER_0_137_472 ();
 sg13g2_fill_2 FILLER_0_137_477 ();
 sg13g2_fill_1 FILLER_0_137_479 ();
 sg13g2_decap_8 FILLER_0_137_495 ();
 sg13g2_decap_8 FILLER_0_137_502 ();
 sg13g2_decap_8 FILLER_0_137_509 ();
 sg13g2_decap_4 FILLER_0_137_516 ();
 sg13g2_fill_1 FILLER_0_137_520 ();
 sg13g2_decap_8 FILLER_0_137_525 ();
 sg13g2_decap_8 FILLER_0_137_532 ();
 sg13g2_decap_8 FILLER_0_137_539 ();
 sg13g2_decap_8 FILLER_0_137_546 ();
 sg13g2_decap_8 FILLER_0_137_553 ();
 sg13g2_decap_8 FILLER_0_137_560 ();
 sg13g2_decap_8 FILLER_0_137_567 ();
 sg13g2_decap_8 FILLER_0_137_574 ();
 sg13g2_decap_8 FILLER_0_137_581 ();
 sg13g2_decap_4 FILLER_0_137_588 ();
 sg13g2_fill_1 FILLER_0_137_592 ();
 sg13g2_decap_8 FILLER_0_137_598 ();
 sg13g2_fill_1 FILLER_0_137_605 ();
 sg13g2_decap_8 FILLER_0_137_642 ();
 sg13g2_decap_8 FILLER_0_137_682 ();
 sg13g2_fill_2 FILLER_0_137_689 ();
 sg13g2_decap_8 FILLER_0_137_705 ();
 sg13g2_decap_8 FILLER_0_137_712 ();
 sg13g2_fill_1 FILLER_0_137_719 ();
 sg13g2_fill_2 FILLER_0_137_767 ();
 sg13g2_fill_1 FILLER_0_137_769 ();
 sg13g2_fill_1 FILLER_0_137_775 ();
 sg13g2_fill_1 FILLER_0_137_793 ();
 sg13g2_fill_2 FILLER_0_137_800 ();
 sg13g2_fill_1 FILLER_0_137_806 ();
 sg13g2_fill_2 FILLER_0_137_817 ();
 sg13g2_fill_1 FILLER_0_137_819 ();
 sg13g2_fill_2 FILLER_0_137_833 ();
 sg13g2_fill_1 FILLER_0_137_842 ();
 sg13g2_fill_1 FILLER_0_137_853 ();
 sg13g2_fill_1 FILLER_0_137_859 ();
 sg13g2_fill_1 FILLER_0_137_868 ();
 sg13g2_fill_2 FILLER_0_137_885 ();
 sg13g2_fill_2 FILLER_0_137_892 ();
 sg13g2_fill_1 FILLER_0_137_899 ();
 sg13g2_fill_2 FILLER_0_137_915 ();
 sg13g2_fill_2 FILLER_0_137_928 ();
 sg13g2_fill_1 FILLER_0_137_953 ();
 sg13g2_fill_1 FILLER_0_137_959 ();
 sg13g2_fill_2 FILLER_0_137_979 ();
 sg13g2_fill_1 FILLER_0_137_981 ();
 sg13g2_decap_8 FILLER_0_137_986 ();
 sg13g2_decap_8 FILLER_0_137_993 ();
 sg13g2_fill_2 FILLER_0_137_1000 ();
 sg13g2_fill_2 FILLER_0_137_1032 ();
 sg13g2_fill_1 FILLER_0_137_1078 ();
 sg13g2_decap_8 FILLER_0_137_1084 ();
 sg13g2_decap_8 FILLER_0_137_1091 ();
 sg13g2_decap_8 FILLER_0_137_1098 ();
 sg13g2_fill_2 FILLER_0_137_1105 ();
 sg13g2_decap_8 FILLER_0_137_1117 ();
 sg13g2_decap_8 FILLER_0_137_1124 ();
 sg13g2_decap_8 FILLER_0_137_1131 ();
 sg13g2_decap_8 FILLER_0_137_1138 ();
 sg13g2_decap_8 FILLER_0_137_1145 ();
 sg13g2_decap_8 FILLER_0_137_1152 ();
 sg13g2_decap_8 FILLER_0_137_1159 ();
 sg13g2_decap_8 FILLER_0_137_1166 ();
 sg13g2_decap_8 FILLER_0_137_1173 ();
 sg13g2_decap_8 FILLER_0_137_1180 ();
 sg13g2_decap_8 FILLER_0_137_1187 ();
 sg13g2_decap_8 FILLER_0_137_1194 ();
 sg13g2_decap_8 FILLER_0_137_1201 ();
 sg13g2_decap_8 FILLER_0_137_1208 ();
 sg13g2_decap_8 FILLER_0_137_1215 ();
 sg13g2_decap_4 FILLER_0_137_1222 ();
 sg13g2_fill_2 FILLER_0_137_1226 ();
 sg13g2_decap_8 FILLER_0_138_0 ();
 sg13g2_decap_8 FILLER_0_138_7 ();
 sg13g2_decap_8 FILLER_0_138_14 ();
 sg13g2_decap_8 FILLER_0_138_21 ();
 sg13g2_fill_1 FILLER_0_138_28 ();
 sg13g2_fill_1 FILLER_0_138_64 ();
 sg13g2_decap_8 FILLER_0_138_130 ();
 sg13g2_decap_8 FILLER_0_138_137 ();
 sg13g2_decap_8 FILLER_0_138_144 ();
 sg13g2_decap_8 FILLER_0_138_151 ();
 sg13g2_decap_4 FILLER_0_138_158 ();
 sg13g2_fill_1 FILLER_0_138_162 ();
 sg13g2_fill_2 FILLER_0_138_194 ();
 sg13g2_decap_8 FILLER_0_138_222 ();
 sg13g2_fill_2 FILLER_0_138_229 ();
 sg13g2_decap_8 FILLER_0_138_235 ();
 sg13g2_decap_8 FILLER_0_138_242 ();
 sg13g2_decap_8 FILLER_0_138_249 ();
 sg13g2_decap_8 FILLER_0_138_256 ();
 sg13g2_decap_8 FILLER_0_138_263 ();
 sg13g2_decap_8 FILLER_0_138_270 ();
 sg13g2_decap_8 FILLER_0_138_277 ();
 sg13g2_decap_8 FILLER_0_138_284 ();
 sg13g2_decap_8 FILLER_0_138_291 ();
 sg13g2_decap_8 FILLER_0_138_298 ();
 sg13g2_decap_8 FILLER_0_138_305 ();
 sg13g2_fill_1 FILLER_0_138_312 ();
 sg13g2_decap_4 FILLER_0_138_348 ();
 sg13g2_decap_8 FILLER_0_138_383 ();
 sg13g2_decap_8 FILLER_0_138_390 ();
 sg13g2_decap_8 FILLER_0_138_397 ();
 sg13g2_decap_8 FILLER_0_138_404 ();
 sg13g2_decap_8 FILLER_0_138_411 ();
 sg13g2_decap_4 FILLER_0_138_418 ();
 sg13g2_fill_1 FILLER_0_138_422 ();
 sg13g2_decap_8 FILLER_0_138_453 ();
 sg13g2_fill_2 FILLER_0_138_460 ();
 sg13g2_fill_1 FILLER_0_138_462 ();
 sg13g2_decap_8 FILLER_0_138_494 ();
 sg13g2_decap_8 FILLER_0_138_501 ();
 sg13g2_decap_8 FILLER_0_138_508 ();
 sg13g2_decap_8 FILLER_0_138_515 ();
 sg13g2_decap_8 FILLER_0_138_522 ();
 sg13g2_decap_8 FILLER_0_138_529 ();
 sg13g2_decap_8 FILLER_0_138_536 ();
 sg13g2_decap_8 FILLER_0_138_543 ();
 sg13g2_decap_8 FILLER_0_138_550 ();
 sg13g2_decap_8 FILLER_0_138_557 ();
 sg13g2_decap_8 FILLER_0_138_564 ();
 sg13g2_decap_8 FILLER_0_138_571 ();
 sg13g2_fill_2 FILLER_0_138_578 ();
 sg13g2_fill_1 FILLER_0_138_585 ();
 sg13g2_decap_4 FILLER_0_138_612 ();
 sg13g2_decap_8 FILLER_0_138_621 ();
 sg13g2_decap_8 FILLER_0_138_628 ();
 sg13g2_decap_4 FILLER_0_138_635 ();
 sg13g2_fill_2 FILLER_0_138_682 ();
 sg13g2_fill_1 FILLER_0_138_684 ();
 sg13g2_fill_2 FILLER_0_138_690 ();
 sg13g2_fill_1 FILLER_0_138_692 ();
 sg13g2_fill_2 FILLER_0_138_712 ();
 sg13g2_decap_4 FILLER_0_138_719 ();
 sg13g2_fill_1 FILLER_0_138_723 ();
 sg13g2_fill_1 FILLER_0_138_737 ();
 sg13g2_decap_4 FILLER_0_138_794 ();
 sg13g2_fill_2 FILLER_0_138_798 ();
 sg13g2_fill_2 FILLER_0_138_804 ();
 sg13g2_fill_1 FILLER_0_138_806 ();
 sg13g2_decap_4 FILLER_0_138_812 ();
 sg13g2_fill_2 FILLER_0_138_816 ();
 sg13g2_fill_1 FILLER_0_138_823 ();
 sg13g2_fill_1 FILLER_0_138_829 ();
 sg13g2_fill_1 FILLER_0_138_835 ();
 sg13g2_fill_1 FILLER_0_138_842 ();
 sg13g2_fill_2 FILLER_0_138_847 ();
 sg13g2_fill_1 FILLER_0_138_854 ();
 sg13g2_fill_2 FILLER_0_138_860 ();
 sg13g2_decap_8 FILLER_0_138_867 ();
 sg13g2_decap_4 FILLER_0_138_874 ();
 sg13g2_fill_2 FILLER_0_138_886 ();
 sg13g2_fill_1 FILLER_0_138_896 ();
 sg13g2_fill_2 FILLER_0_138_902 ();
 sg13g2_fill_2 FILLER_0_138_909 ();
 sg13g2_fill_1 FILLER_0_138_916 ();
 sg13g2_fill_1 FILLER_0_138_923 ();
 sg13g2_fill_1 FILLER_0_138_930 ();
 sg13g2_decap_4 FILLER_0_138_968 ();
 sg13g2_fill_1 FILLER_0_138_980 ();
 sg13g2_fill_2 FILLER_0_138_991 ();
 sg13g2_fill_1 FILLER_0_138_993 ();
 sg13g2_fill_2 FILLER_0_138_1004 ();
 sg13g2_fill_1 FILLER_0_138_1079 ();
 sg13g2_fill_2 FILLER_0_138_1085 ();
 sg13g2_fill_1 FILLER_0_138_1087 ();
 sg13g2_decap_8 FILLER_0_138_1119 ();
 sg13g2_decap_8 FILLER_0_138_1126 ();
 sg13g2_decap_8 FILLER_0_138_1133 ();
 sg13g2_decap_8 FILLER_0_138_1140 ();
 sg13g2_decap_8 FILLER_0_138_1147 ();
 sg13g2_decap_8 FILLER_0_138_1154 ();
 sg13g2_decap_8 FILLER_0_138_1161 ();
 sg13g2_decap_8 FILLER_0_138_1168 ();
 sg13g2_decap_8 FILLER_0_138_1175 ();
 sg13g2_decap_8 FILLER_0_138_1182 ();
 sg13g2_decap_8 FILLER_0_138_1189 ();
 sg13g2_decap_8 FILLER_0_138_1196 ();
 sg13g2_decap_8 FILLER_0_138_1203 ();
 sg13g2_decap_8 FILLER_0_138_1210 ();
 sg13g2_decap_8 FILLER_0_138_1217 ();
 sg13g2_decap_4 FILLER_0_138_1224 ();
 sg13g2_decap_8 FILLER_0_139_0 ();
 sg13g2_decap_8 FILLER_0_139_7 ();
 sg13g2_decap_8 FILLER_0_139_14 ();
 sg13g2_decap_8 FILLER_0_139_21 ();
 sg13g2_fill_2 FILLER_0_139_28 ();
 sg13g2_fill_1 FILLER_0_139_30 ();
 sg13g2_fill_1 FILLER_0_139_36 ();
 sg13g2_decap_8 FILLER_0_139_47 ();
 sg13g2_decap_4 FILLER_0_139_54 ();
 sg13g2_fill_2 FILLER_0_139_58 ();
 sg13g2_fill_1 FILLER_0_139_79 ();
 sg13g2_decap_8 FILLER_0_139_124 ();
 sg13g2_decap_8 FILLER_0_139_131 ();
 sg13g2_decap_8 FILLER_0_139_138 ();
 sg13g2_decap_8 FILLER_0_139_145 ();
 sg13g2_decap_8 FILLER_0_139_152 ();
 sg13g2_decap_8 FILLER_0_139_159 ();
 sg13g2_decap_8 FILLER_0_139_166 ();
 sg13g2_fill_1 FILLER_0_139_173 ();
 sg13g2_fill_1 FILLER_0_139_178 ();
 sg13g2_fill_1 FILLER_0_139_210 ();
 sg13g2_decap_8 FILLER_0_139_237 ();
 sg13g2_decap_8 FILLER_0_139_244 ();
 sg13g2_decap_8 FILLER_0_139_251 ();
 sg13g2_decap_8 FILLER_0_139_258 ();
 sg13g2_decap_8 FILLER_0_139_265 ();
 sg13g2_decap_8 FILLER_0_139_272 ();
 sg13g2_decap_8 FILLER_0_139_279 ();
 sg13g2_decap_8 FILLER_0_139_286 ();
 sg13g2_decap_8 FILLER_0_139_293 ();
 sg13g2_decap_8 FILLER_0_139_300 ();
 sg13g2_decap_8 FILLER_0_139_307 ();
 sg13g2_fill_2 FILLER_0_139_314 ();
 sg13g2_decap_8 FILLER_0_139_321 ();
 sg13g2_decap_8 FILLER_0_139_328 ();
 sg13g2_decap_4 FILLER_0_139_335 ();
 sg13g2_fill_1 FILLER_0_139_339 ();
 sg13g2_fill_2 FILLER_0_139_350 ();
 sg13g2_fill_1 FILLER_0_139_357 ();
 sg13g2_decap_8 FILLER_0_139_372 ();
 sg13g2_decap_8 FILLER_0_139_379 ();
 sg13g2_decap_8 FILLER_0_139_386 ();
 sg13g2_decap_8 FILLER_0_139_393 ();
 sg13g2_decap_8 FILLER_0_139_400 ();
 sg13g2_decap_8 FILLER_0_139_407 ();
 sg13g2_decap_8 FILLER_0_139_414 ();
 sg13g2_fill_1 FILLER_0_139_421 ();
 sg13g2_fill_2 FILLER_0_139_453 ();
 sg13g2_fill_1 FILLER_0_139_455 ();
 sg13g2_decap_8 FILLER_0_139_500 ();
 sg13g2_decap_8 FILLER_0_139_507 ();
 sg13g2_decap_8 FILLER_0_139_514 ();
 sg13g2_decap_8 FILLER_0_139_521 ();
 sg13g2_decap_8 FILLER_0_139_528 ();
 sg13g2_decap_8 FILLER_0_139_535 ();
 sg13g2_decap_8 FILLER_0_139_542 ();
 sg13g2_decap_8 FILLER_0_139_549 ();
 sg13g2_decap_8 FILLER_0_139_556 ();
 sg13g2_decap_4 FILLER_0_139_563 ();
 sg13g2_fill_2 FILLER_0_139_567 ();
 sg13g2_fill_2 FILLER_0_139_628 ();
 sg13g2_fill_1 FILLER_0_139_712 ();
 sg13g2_fill_1 FILLER_0_139_750 ();
 sg13g2_fill_2 FILLER_0_139_769 ();
 sg13g2_fill_2 FILLER_0_139_780 ();
 sg13g2_fill_1 FILLER_0_139_782 ();
 sg13g2_fill_1 FILLER_0_139_806 ();
 sg13g2_decap_8 FILLER_0_139_821 ();
 sg13g2_decap_8 FILLER_0_139_828 ();
 sg13g2_decap_8 FILLER_0_139_835 ();
 sg13g2_decap_4 FILLER_0_139_842 ();
 sg13g2_fill_1 FILLER_0_139_846 ();
 sg13g2_decap_8 FILLER_0_139_852 ();
 sg13g2_decap_4 FILLER_0_139_859 ();
 sg13g2_fill_1 FILLER_0_139_863 ();
 sg13g2_decap_4 FILLER_0_139_872 ();
 sg13g2_fill_2 FILLER_0_139_895 ();
 sg13g2_fill_1 FILLER_0_139_897 ();
 sg13g2_decap_8 FILLER_0_139_908 ();
 sg13g2_decap_4 FILLER_0_139_915 ();
 sg13g2_fill_2 FILLER_0_139_919 ();
 sg13g2_fill_1 FILLER_0_139_925 ();
 sg13g2_fill_2 FILLER_0_139_940 ();
 sg13g2_fill_1 FILLER_0_139_942 ();
 sg13g2_fill_2 FILLER_0_139_953 ();
 sg13g2_fill_2 FILLER_0_139_989 ();
 sg13g2_fill_1 FILLER_0_139_1010 ();
 sg13g2_decap_4 FILLER_0_139_1038 ();
 sg13g2_fill_2 FILLER_0_139_1042 ();
 sg13g2_fill_1 FILLER_0_139_1048 ();
 sg13g2_fill_1 FILLER_0_139_1054 ();
 sg13g2_fill_1 FILLER_0_139_1059 ();
 sg13g2_fill_2 FILLER_0_139_1064 ();
 sg13g2_decap_8 FILLER_0_139_1072 ();
 sg13g2_decap_8 FILLER_0_139_1079 ();
 sg13g2_decap_4 FILLER_0_139_1086 ();
 sg13g2_fill_2 FILLER_0_139_1090 ();
 sg13g2_decap_8 FILLER_0_139_1096 ();
 sg13g2_decap_8 FILLER_0_139_1103 ();
 sg13g2_decap_8 FILLER_0_139_1110 ();
 sg13g2_decap_8 FILLER_0_139_1117 ();
 sg13g2_decap_8 FILLER_0_139_1124 ();
 sg13g2_decap_8 FILLER_0_139_1131 ();
 sg13g2_decap_8 FILLER_0_139_1138 ();
 sg13g2_decap_8 FILLER_0_139_1145 ();
 sg13g2_decap_8 FILLER_0_139_1152 ();
 sg13g2_decap_8 FILLER_0_139_1159 ();
 sg13g2_decap_8 FILLER_0_139_1166 ();
 sg13g2_decap_8 FILLER_0_139_1173 ();
 sg13g2_decap_8 FILLER_0_139_1180 ();
 sg13g2_decap_8 FILLER_0_139_1187 ();
 sg13g2_decap_8 FILLER_0_139_1194 ();
 sg13g2_decap_8 FILLER_0_139_1201 ();
 sg13g2_decap_8 FILLER_0_139_1208 ();
 sg13g2_decap_8 FILLER_0_139_1215 ();
 sg13g2_decap_4 FILLER_0_139_1222 ();
 sg13g2_fill_2 FILLER_0_139_1226 ();
 sg13g2_decap_8 FILLER_0_140_0 ();
 sg13g2_decap_8 FILLER_0_140_7 ();
 sg13g2_decap_8 FILLER_0_140_14 ();
 sg13g2_decap_8 FILLER_0_140_21 ();
 sg13g2_fill_1 FILLER_0_140_28 ();
 sg13g2_decap_8 FILLER_0_140_64 ();
 sg13g2_decap_8 FILLER_0_140_71 ();
 sg13g2_decap_8 FILLER_0_140_78 ();
 sg13g2_decap_8 FILLER_0_140_85 ();
 sg13g2_decap_8 FILLER_0_140_92 ();
 sg13g2_fill_2 FILLER_0_140_99 ();
 sg13g2_decap_8 FILLER_0_140_104 ();
 sg13g2_decap_8 FILLER_0_140_111 ();
 sg13g2_decap_8 FILLER_0_140_118 ();
 sg13g2_decap_8 FILLER_0_140_125 ();
 sg13g2_decap_8 FILLER_0_140_132 ();
 sg13g2_decap_8 FILLER_0_140_139 ();
 sg13g2_decap_8 FILLER_0_140_146 ();
 sg13g2_decap_8 FILLER_0_140_153 ();
 sg13g2_decap_8 FILLER_0_140_160 ();
 sg13g2_decap_8 FILLER_0_140_167 ();
 sg13g2_decap_4 FILLER_0_140_174 ();
 sg13g2_fill_1 FILLER_0_140_187 ();
 sg13g2_fill_1 FILLER_0_140_223 ();
 sg13g2_decap_8 FILLER_0_140_228 ();
 sg13g2_decap_8 FILLER_0_140_235 ();
 sg13g2_decap_8 FILLER_0_140_242 ();
 sg13g2_decap_8 FILLER_0_140_249 ();
 sg13g2_decap_8 FILLER_0_140_256 ();
 sg13g2_decap_8 FILLER_0_140_263 ();
 sg13g2_decap_8 FILLER_0_140_270 ();
 sg13g2_decap_8 FILLER_0_140_277 ();
 sg13g2_decap_8 FILLER_0_140_284 ();
 sg13g2_decap_8 FILLER_0_140_291 ();
 sg13g2_decap_8 FILLER_0_140_298 ();
 sg13g2_decap_4 FILLER_0_140_305 ();
 sg13g2_decap_8 FILLER_0_140_388 ();
 sg13g2_decap_8 FILLER_0_140_395 ();
 sg13g2_decap_8 FILLER_0_140_402 ();
 sg13g2_decap_8 FILLER_0_140_409 ();
 sg13g2_decap_8 FILLER_0_140_416 ();
 sg13g2_decap_4 FILLER_0_140_423 ();
 sg13g2_fill_2 FILLER_0_140_442 ();
 sg13g2_decap_4 FILLER_0_140_459 ();
 sg13g2_decap_8 FILLER_0_140_499 ();
 sg13g2_decap_8 FILLER_0_140_506 ();
 sg13g2_decap_8 FILLER_0_140_513 ();
 sg13g2_decap_8 FILLER_0_140_520 ();
 sg13g2_decap_8 FILLER_0_140_527 ();
 sg13g2_decap_8 FILLER_0_140_534 ();
 sg13g2_decap_8 FILLER_0_140_541 ();
 sg13g2_decap_8 FILLER_0_140_548 ();
 sg13g2_decap_8 FILLER_0_140_555 ();
 sg13g2_decap_8 FILLER_0_140_562 ();
 sg13g2_decap_4 FILLER_0_140_569 ();
 sg13g2_fill_1 FILLER_0_140_582 ();
 sg13g2_fill_1 FILLER_0_140_593 ();
 sg13g2_decap_8 FILLER_0_140_623 ();
 sg13g2_decap_8 FILLER_0_140_630 ();
 sg13g2_decap_8 FILLER_0_140_637 ();
 sg13g2_fill_2 FILLER_0_140_644 ();
 sg13g2_fill_2 FILLER_0_140_656 ();
 sg13g2_fill_1 FILLER_0_140_658 ();
 sg13g2_decap_8 FILLER_0_140_681 ();
 sg13g2_decap_8 FILLER_0_140_717 ();
 sg13g2_fill_2 FILLER_0_140_733 ();
 sg13g2_fill_2 FILLER_0_140_759 ();
 sg13g2_fill_1 FILLER_0_140_766 ();
 sg13g2_fill_2 FILLER_0_140_787 ();
 sg13g2_fill_2 FILLER_0_140_801 ();
 sg13g2_fill_2 FILLER_0_140_807 ();
 sg13g2_fill_1 FILLER_0_140_817 ();
 sg13g2_fill_1 FILLER_0_140_823 ();
 sg13g2_decap_4 FILLER_0_140_834 ();
 sg13g2_fill_2 FILLER_0_140_842 ();
 sg13g2_fill_1 FILLER_0_140_848 ();
 sg13g2_decap_8 FILLER_0_140_863 ();
 sg13g2_decap_4 FILLER_0_140_870 ();
 sg13g2_fill_2 FILLER_0_140_874 ();
 sg13g2_fill_2 FILLER_0_140_884 ();
 sg13g2_fill_2 FILLER_0_140_896 ();
 sg13g2_decap_8 FILLER_0_140_903 ();
 sg13g2_fill_2 FILLER_0_140_910 ();
 sg13g2_fill_1 FILLER_0_140_912 ();
 sg13g2_decap_4 FILLER_0_140_918 ();
 sg13g2_fill_1 FILLER_0_140_922 ();
 sg13g2_decap_4 FILLER_0_140_939 ();
 sg13g2_decap_4 FILLER_0_140_947 ();
 sg13g2_fill_2 FILLER_0_140_958 ();
 sg13g2_decap_4 FILLER_0_140_975 ();
 sg13g2_decap_4 FILLER_0_140_1000 ();
 sg13g2_fill_2 FILLER_0_140_1004 ();
 sg13g2_decap_4 FILLER_0_140_1014 ();
 sg13g2_decap_8 FILLER_0_140_1022 ();
 sg13g2_decap_8 FILLER_0_140_1029 ();
 sg13g2_fill_2 FILLER_0_140_1036 ();
 sg13g2_decap_4 FILLER_0_140_1042 ();
 sg13g2_decap_4 FILLER_0_140_1054 ();
 sg13g2_fill_2 FILLER_0_140_1062 ();
 sg13g2_decap_8 FILLER_0_140_1069 ();
 sg13g2_decap_8 FILLER_0_140_1076 ();
 sg13g2_decap_8 FILLER_0_140_1083 ();
 sg13g2_fill_2 FILLER_0_140_1090 ();
 sg13g2_fill_1 FILLER_0_140_1092 ();
 sg13g2_decap_8 FILLER_0_140_1098 ();
 sg13g2_fill_2 FILLER_0_140_1105 ();
 sg13g2_fill_1 FILLER_0_140_1107 ();
 sg13g2_decap_8 FILLER_0_140_1118 ();
 sg13g2_decap_8 FILLER_0_140_1125 ();
 sg13g2_decap_8 FILLER_0_140_1132 ();
 sg13g2_decap_8 FILLER_0_140_1139 ();
 sg13g2_decap_8 FILLER_0_140_1146 ();
 sg13g2_decap_8 FILLER_0_140_1153 ();
 sg13g2_decap_8 FILLER_0_140_1160 ();
 sg13g2_decap_8 FILLER_0_140_1167 ();
 sg13g2_decap_8 FILLER_0_140_1174 ();
 sg13g2_decap_8 FILLER_0_140_1181 ();
 sg13g2_decap_8 FILLER_0_140_1188 ();
 sg13g2_decap_8 FILLER_0_140_1195 ();
 sg13g2_decap_8 FILLER_0_140_1202 ();
 sg13g2_decap_8 FILLER_0_140_1209 ();
 sg13g2_decap_8 FILLER_0_140_1216 ();
 sg13g2_decap_4 FILLER_0_140_1223 ();
 sg13g2_fill_1 FILLER_0_140_1227 ();
 sg13g2_decap_8 FILLER_0_141_0 ();
 sg13g2_decap_8 FILLER_0_141_7 ();
 sg13g2_decap_4 FILLER_0_141_14 ();
 sg13g2_fill_1 FILLER_0_141_18 ();
 sg13g2_fill_2 FILLER_0_141_34 ();
 sg13g2_decap_8 FILLER_0_141_51 ();
 sg13g2_decap_8 FILLER_0_141_58 ();
 sg13g2_decap_4 FILLER_0_141_65 ();
 sg13g2_fill_1 FILLER_0_141_69 ();
 sg13g2_decap_8 FILLER_0_141_104 ();
 sg13g2_decap_8 FILLER_0_141_111 ();
 sg13g2_decap_8 FILLER_0_141_118 ();
 sg13g2_decap_8 FILLER_0_141_125 ();
 sg13g2_decap_8 FILLER_0_141_132 ();
 sg13g2_decap_8 FILLER_0_141_139 ();
 sg13g2_decap_8 FILLER_0_141_146 ();
 sg13g2_decap_8 FILLER_0_141_153 ();
 sg13g2_decap_8 FILLER_0_141_160 ();
 sg13g2_decap_8 FILLER_0_141_167 ();
 sg13g2_decap_8 FILLER_0_141_174 ();
 sg13g2_decap_8 FILLER_0_141_181 ();
 sg13g2_decap_8 FILLER_0_141_188 ();
 sg13g2_decap_8 FILLER_0_141_195 ();
 sg13g2_decap_8 FILLER_0_141_202 ();
 sg13g2_decap_8 FILLER_0_141_209 ();
 sg13g2_decap_8 FILLER_0_141_216 ();
 sg13g2_decap_8 FILLER_0_141_223 ();
 sg13g2_decap_8 FILLER_0_141_230 ();
 sg13g2_decap_8 FILLER_0_141_237 ();
 sg13g2_decap_8 FILLER_0_141_244 ();
 sg13g2_decap_8 FILLER_0_141_251 ();
 sg13g2_decap_8 FILLER_0_141_258 ();
 sg13g2_decap_8 FILLER_0_141_265 ();
 sg13g2_decap_8 FILLER_0_141_272 ();
 sg13g2_decap_8 FILLER_0_141_279 ();
 sg13g2_decap_8 FILLER_0_141_286 ();
 sg13g2_decap_8 FILLER_0_141_293 ();
 sg13g2_decap_8 FILLER_0_141_300 ();
 sg13g2_decap_8 FILLER_0_141_307 ();
 sg13g2_decap_8 FILLER_0_141_327 ();
 sg13g2_fill_1 FILLER_0_141_334 ();
 sg13g2_fill_1 FILLER_0_141_345 ();
 sg13g2_fill_2 FILLER_0_141_354 ();
 sg13g2_decap_8 FILLER_0_141_395 ();
 sg13g2_decap_8 FILLER_0_141_402 ();
 sg13g2_decap_8 FILLER_0_141_409 ();
 sg13g2_decap_8 FILLER_0_141_416 ();
 sg13g2_decap_8 FILLER_0_141_423 ();
 sg13g2_decap_8 FILLER_0_141_434 ();
 sg13g2_decap_8 FILLER_0_141_441 ();
 sg13g2_decap_8 FILLER_0_141_448 ();
 sg13g2_decap_4 FILLER_0_141_455 ();
 sg13g2_fill_2 FILLER_0_141_459 ();
 sg13g2_decap_4 FILLER_0_141_465 ();
 sg13g2_fill_2 FILLER_0_141_469 ();
 sg13g2_decap_8 FILLER_0_141_475 ();
 sg13g2_decap_8 FILLER_0_141_482 ();
 sg13g2_decap_8 FILLER_0_141_489 ();
 sg13g2_decap_8 FILLER_0_141_496 ();
 sg13g2_decap_8 FILLER_0_141_503 ();
 sg13g2_decap_8 FILLER_0_141_510 ();
 sg13g2_decap_8 FILLER_0_141_517 ();
 sg13g2_decap_8 FILLER_0_141_524 ();
 sg13g2_decap_8 FILLER_0_141_531 ();
 sg13g2_decap_8 FILLER_0_141_538 ();
 sg13g2_decap_8 FILLER_0_141_545 ();
 sg13g2_decap_8 FILLER_0_141_552 ();
 sg13g2_decap_8 FILLER_0_141_559 ();
 sg13g2_decap_8 FILLER_0_141_566 ();
 sg13g2_fill_1 FILLER_0_141_615 ();
 sg13g2_decap_4 FILLER_0_141_647 ();
 sg13g2_fill_2 FILLER_0_141_651 ();
 sg13g2_fill_1 FILLER_0_141_684 ();
 sg13g2_fill_2 FILLER_0_141_690 ();
 sg13g2_fill_1 FILLER_0_141_696 ();
 sg13g2_fill_1 FILLER_0_141_722 ();
 sg13g2_fill_2 FILLER_0_141_726 ();
 sg13g2_fill_1 FILLER_0_141_743 ();
 sg13g2_fill_1 FILLER_0_141_749 ();
 sg13g2_fill_2 FILLER_0_141_796 ();
 sg13g2_fill_1 FILLER_0_141_798 ();
 sg13g2_fill_1 FILLER_0_141_833 ();
 sg13g2_fill_1 FILLER_0_141_858 ();
 sg13g2_fill_1 FILLER_0_141_864 ();
 sg13g2_fill_1 FILLER_0_141_873 ();
 sg13g2_fill_1 FILLER_0_141_880 ();
 sg13g2_fill_1 FILLER_0_141_886 ();
 sg13g2_fill_1 FILLER_0_141_895 ();
 sg13g2_fill_1 FILLER_0_141_929 ();
 sg13g2_fill_2 FILLER_0_141_935 ();
 sg13g2_fill_1 FILLER_0_141_937 ();
 sg13g2_fill_2 FILLER_0_141_942 ();
 sg13g2_fill_1 FILLER_0_141_944 ();
 sg13g2_fill_1 FILLER_0_141_953 ();
 sg13g2_fill_1 FILLER_0_141_962 ();
 sg13g2_fill_1 FILLER_0_141_968 ();
 sg13g2_decap_4 FILLER_0_141_977 ();
 sg13g2_decap_4 FILLER_0_141_985 ();
 sg13g2_decap_8 FILLER_0_141_994 ();
 sg13g2_fill_2 FILLER_0_141_1001 ();
 sg13g2_fill_1 FILLER_0_141_1003 ();
 sg13g2_fill_2 FILLER_0_141_1007 ();
 sg13g2_fill_1 FILLER_0_141_1009 ();
 sg13g2_fill_2 FILLER_0_141_1028 ();
 sg13g2_fill_1 FILLER_0_141_1030 ();
 sg13g2_decap_8 FILLER_0_141_1041 ();
 sg13g2_decap_8 FILLER_0_141_1048 ();
 sg13g2_decap_8 FILLER_0_141_1055 ();
 sg13g2_decap_8 FILLER_0_141_1062 ();
 sg13g2_decap_8 FILLER_0_141_1069 ();
 sg13g2_decap_8 FILLER_0_141_1076 ();
 sg13g2_decap_4 FILLER_0_141_1083 ();
 sg13g2_decap_8 FILLER_0_141_1118 ();
 sg13g2_decap_8 FILLER_0_141_1125 ();
 sg13g2_decap_8 FILLER_0_141_1132 ();
 sg13g2_decap_8 FILLER_0_141_1139 ();
 sg13g2_decap_8 FILLER_0_141_1146 ();
 sg13g2_decap_8 FILLER_0_141_1153 ();
 sg13g2_decap_8 FILLER_0_141_1160 ();
 sg13g2_decap_8 FILLER_0_141_1167 ();
 sg13g2_decap_8 FILLER_0_141_1174 ();
 sg13g2_decap_8 FILLER_0_141_1181 ();
 sg13g2_decap_8 FILLER_0_141_1188 ();
 sg13g2_decap_8 FILLER_0_141_1195 ();
 sg13g2_decap_8 FILLER_0_141_1202 ();
 sg13g2_decap_8 FILLER_0_141_1209 ();
 sg13g2_decap_8 FILLER_0_141_1216 ();
 sg13g2_decap_4 FILLER_0_141_1223 ();
 sg13g2_fill_1 FILLER_0_141_1227 ();
 sg13g2_decap_8 FILLER_0_142_0 ();
 sg13g2_decap_4 FILLER_0_142_7 ();
 sg13g2_fill_2 FILLER_0_142_11 ();
 sg13g2_decap_4 FILLER_0_142_52 ();
 sg13g2_fill_2 FILLER_0_142_56 ();
 sg13g2_fill_1 FILLER_0_142_91 ();
 sg13g2_decap_8 FILLER_0_142_118 ();
 sg13g2_decap_8 FILLER_0_142_125 ();
 sg13g2_decap_8 FILLER_0_142_132 ();
 sg13g2_decap_8 FILLER_0_142_139 ();
 sg13g2_decap_8 FILLER_0_142_146 ();
 sg13g2_decap_8 FILLER_0_142_153 ();
 sg13g2_decap_8 FILLER_0_142_160 ();
 sg13g2_decap_8 FILLER_0_142_167 ();
 sg13g2_decap_8 FILLER_0_142_174 ();
 sg13g2_decap_8 FILLER_0_142_181 ();
 sg13g2_decap_8 FILLER_0_142_188 ();
 sg13g2_decap_8 FILLER_0_142_195 ();
 sg13g2_decap_8 FILLER_0_142_202 ();
 sg13g2_decap_8 FILLER_0_142_209 ();
 sg13g2_decap_8 FILLER_0_142_216 ();
 sg13g2_decap_8 FILLER_0_142_223 ();
 sg13g2_decap_8 FILLER_0_142_230 ();
 sg13g2_decap_8 FILLER_0_142_237 ();
 sg13g2_decap_8 FILLER_0_142_244 ();
 sg13g2_decap_8 FILLER_0_142_251 ();
 sg13g2_decap_8 FILLER_0_142_258 ();
 sg13g2_decap_8 FILLER_0_142_265 ();
 sg13g2_decap_8 FILLER_0_142_272 ();
 sg13g2_decap_8 FILLER_0_142_279 ();
 sg13g2_decap_8 FILLER_0_142_286 ();
 sg13g2_decap_8 FILLER_0_142_293 ();
 sg13g2_decap_8 FILLER_0_142_300 ();
 sg13g2_decap_4 FILLER_0_142_307 ();
 sg13g2_fill_1 FILLER_0_142_311 ();
 sg13g2_fill_1 FILLER_0_142_351 ();
 sg13g2_decap_8 FILLER_0_142_381 ();
 sg13g2_decap_8 FILLER_0_142_388 ();
 sg13g2_decap_8 FILLER_0_142_395 ();
 sg13g2_decap_8 FILLER_0_142_402 ();
 sg13g2_decap_8 FILLER_0_142_409 ();
 sg13g2_decap_8 FILLER_0_142_416 ();
 sg13g2_decap_8 FILLER_0_142_423 ();
 sg13g2_decap_8 FILLER_0_142_430 ();
 sg13g2_decap_8 FILLER_0_142_437 ();
 sg13g2_decap_8 FILLER_0_142_444 ();
 sg13g2_decap_8 FILLER_0_142_451 ();
 sg13g2_decap_8 FILLER_0_142_458 ();
 sg13g2_decap_8 FILLER_0_142_465 ();
 sg13g2_decap_8 FILLER_0_142_472 ();
 sg13g2_decap_8 FILLER_0_142_479 ();
 sg13g2_decap_8 FILLER_0_142_486 ();
 sg13g2_decap_8 FILLER_0_142_493 ();
 sg13g2_decap_8 FILLER_0_142_500 ();
 sg13g2_decap_8 FILLER_0_142_507 ();
 sg13g2_decap_8 FILLER_0_142_514 ();
 sg13g2_decap_8 FILLER_0_142_521 ();
 sg13g2_decap_8 FILLER_0_142_528 ();
 sg13g2_decap_8 FILLER_0_142_535 ();
 sg13g2_decap_8 FILLER_0_142_542 ();
 sg13g2_decap_8 FILLER_0_142_549 ();
 sg13g2_decap_8 FILLER_0_142_556 ();
 sg13g2_decap_8 FILLER_0_142_563 ();
 sg13g2_decap_8 FILLER_0_142_570 ();
 sg13g2_fill_1 FILLER_0_142_577 ();
 sg13g2_fill_2 FILLER_0_142_618 ();
 sg13g2_fill_1 FILLER_0_142_620 ();
 sg13g2_fill_2 FILLER_0_142_626 ();
 sg13g2_decap_8 FILLER_0_142_632 ();
 sg13g2_decap_8 FILLER_0_142_639 ();
 sg13g2_fill_2 FILLER_0_142_646 ();
 sg13g2_decap_8 FILLER_0_142_652 ();
 sg13g2_fill_1 FILLER_0_142_659 ();
 sg13g2_fill_2 FILLER_0_142_670 ();
 sg13g2_fill_1 FILLER_0_142_722 ();
 sg13g2_fill_2 FILLER_0_142_784 ();
 sg13g2_fill_2 FILLER_0_142_823 ();
 sg13g2_fill_1 FILLER_0_142_850 ();
 sg13g2_fill_2 FILLER_0_142_859 ();
 sg13g2_fill_1 FILLER_0_142_861 ();
 sg13g2_fill_2 FILLER_0_142_876 ();
 sg13g2_fill_1 FILLER_0_142_878 ();
 sg13g2_decap_4 FILLER_0_142_904 ();
 sg13g2_fill_2 FILLER_0_142_908 ();
 sg13g2_decap_4 FILLER_0_142_928 ();
 sg13g2_fill_2 FILLER_0_142_937 ();
 sg13g2_fill_1 FILLER_0_142_956 ();
 sg13g2_fill_2 FILLER_0_142_966 ();
 sg13g2_fill_1 FILLER_0_142_968 ();
 sg13g2_decap_4 FILLER_0_142_974 ();
 sg13g2_fill_1 FILLER_0_142_978 ();
 sg13g2_decap_8 FILLER_0_142_984 ();
 sg13g2_decap_4 FILLER_0_142_991 ();
 sg13g2_fill_1 FILLER_0_142_1028 ();
 sg13g2_decap_8 FILLER_0_142_1047 ();
 sg13g2_decap_8 FILLER_0_142_1054 ();
 sg13g2_decap_8 FILLER_0_142_1061 ();
 sg13g2_decap_8 FILLER_0_142_1068 ();
 sg13g2_decap_8 FILLER_0_142_1075 ();
 sg13g2_decap_8 FILLER_0_142_1082 ();
 sg13g2_fill_2 FILLER_0_142_1089 ();
 sg13g2_fill_1 FILLER_0_142_1091 ();
 sg13g2_decap_8 FILLER_0_142_1115 ();
 sg13g2_decap_8 FILLER_0_142_1122 ();
 sg13g2_decap_8 FILLER_0_142_1129 ();
 sg13g2_decap_8 FILLER_0_142_1136 ();
 sg13g2_decap_8 FILLER_0_142_1143 ();
 sg13g2_decap_8 FILLER_0_142_1150 ();
 sg13g2_decap_8 FILLER_0_142_1157 ();
 sg13g2_decap_8 FILLER_0_142_1164 ();
 sg13g2_decap_8 FILLER_0_142_1171 ();
 sg13g2_decap_8 FILLER_0_142_1178 ();
 sg13g2_decap_8 FILLER_0_142_1185 ();
 sg13g2_decap_8 FILLER_0_142_1192 ();
 sg13g2_decap_8 FILLER_0_142_1199 ();
 sg13g2_decap_8 FILLER_0_142_1206 ();
 sg13g2_decap_8 FILLER_0_142_1213 ();
 sg13g2_decap_8 FILLER_0_142_1220 ();
 sg13g2_fill_1 FILLER_0_142_1227 ();
 sg13g2_decap_4 FILLER_0_143_0 ();
 sg13g2_fill_2 FILLER_0_143_4 ();
 sg13g2_decap_4 FILLER_0_143_42 ();
 sg13g2_fill_1 FILLER_0_143_46 ();
 sg13g2_fill_1 FILLER_0_143_52 ();
 sg13g2_fill_1 FILLER_0_143_79 ();
 sg13g2_fill_1 FILLER_0_143_85 ();
 sg13g2_fill_2 FILLER_0_143_90 ();
 sg13g2_fill_2 FILLER_0_143_97 ();
 sg13g2_fill_2 FILLER_0_143_103 ();
 sg13g2_decap_8 FILLER_0_143_136 ();
 sg13g2_decap_8 FILLER_0_143_143 ();
 sg13g2_decap_8 FILLER_0_143_150 ();
 sg13g2_decap_8 FILLER_0_143_157 ();
 sg13g2_decap_8 FILLER_0_143_164 ();
 sg13g2_decap_8 FILLER_0_143_171 ();
 sg13g2_decap_8 FILLER_0_143_178 ();
 sg13g2_decap_8 FILLER_0_143_185 ();
 sg13g2_decap_8 FILLER_0_143_192 ();
 sg13g2_decap_8 FILLER_0_143_199 ();
 sg13g2_decap_8 FILLER_0_143_206 ();
 sg13g2_decap_8 FILLER_0_143_213 ();
 sg13g2_decap_8 FILLER_0_143_220 ();
 sg13g2_decap_8 FILLER_0_143_227 ();
 sg13g2_decap_8 FILLER_0_143_234 ();
 sg13g2_decap_8 FILLER_0_143_241 ();
 sg13g2_decap_8 FILLER_0_143_248 ();
 sg13g2_decap_8 FILLER_0_143_255 ();
 sg13g2_decap_8 FILLER_0_143_262 ();
 sg13g2_decap_8 FILLER_0_143_269 ();
 sg13g2_decap_8 FILLER_0_143_276 ();
 sg13g2_decap_8 FILLER_0_143_283 ();
 sg13g2_decap_8 FILLER_0_143_290 ();
 sg13g2_decap_8 FILLER_0_143_297 ();
 sg13g2_decap_8 FILLER_0_143_304 ();
 sg13g2_fill_2 FILLER_0_143_342 ();
 sg13g2_fill_1 FILLER_0_143_344 ();
 sg13g2_decap_8 FILLER_0_143_381 ();
 sg13g2_decap_8 FILLER_0_143_388 ();
 sg13g2_decap_8 FILLER_0_143_395 ();
 sg13g2_decap_8 FILLER_0_143_402 ();
 sg13g2_decap_8 FILLER_0_143_409 ();
 sg13g2_decap_8 FILLER_0_143_416 ();
 sg13g2_decap_8 FILLER_0_143_423 ();
 sg13g2_decap_8 FILLER_0_143_430 ();
 sg13g2_decap_8 FILLER_0_143_437 ();
 sg13g2_decap_8 FILLER_0_143_444 ();
 sg13g2_decap_8 FILLER_0_143_451 ();
 sg13g2_decap_8 FILLER_0_143_458 ();
 sg13g2_decap_8 FILLER_0_143_465 ();
 sg13g2_decap_8 FILLER_0_143_472 ();
 sg13g2_decap_8 FILLER_0_143_479 ();
 sg13g2_decap_8 FILLER_0_143_486 ();
 sg13g2_decap_8 FILLER_0_143_493 ();
 sg13g2_decap_8 FILLER_0_143_500 ();
 sg13g2_decap_8 FILLER_0_143_507 ();
 sg13g2_decap_8 FILLER_0_143_514 ();
 sg13g2_decap_8 FILLER_0_143_521 ();
 sg13g2_decap_8 FILLER_0_143_528 ();
 sg13g2_decap_8 FILLER_0_143_535 ();
 sg13g2_decap_8 FILLER_0_143_542 ();
 sg13g2_decap_8 FILLER_0_143_549 ();
 sg13g2_decap_8 FILLER_0_143_556 ();
 sg13g2_decap_8 FILLER_0_143_563 ();
 sg13g2_fill_2 FILLER_0_143_570 ();
 sg13g2_fill_1 FILLER_0_143_572 ();
 sg13g2_decap_8 FILLER_0_143_577 ();
 sg13g2_fill_2 FILLER_0_143_584 ();
 sg13g2_fill_2 FILLER_0_143_591 ();
 sg13g2_fill_1 FILLER_0_143_593 ();
 sg13g2_decap_8 FILLER_0_143_603 ();
 sg13g2_decap_4 FILLER_0_143_636 ();
 sg13g2_fill_1 FILLER_0_143_640 ();
 sg13g2_fill_1 FILLER_0_143_672 ();
 sg13g2_decap_8 FILLER_0_143_677 ();
 sg13g2_fill_1 FILLER_0_143_703 ();
 sg13g2_fill_1 FILLER_0_143_712 ();
 sg13g2_fill_2 FILLER_0_143_729 ();
 sg13g2_fill_2 FILLER_0_143_800 ();
 sg13g2_decap_8 FILLER_0_143_819 ();
 sg13g2_decap_8 FILLER_0_143_826 ();
 sg13g2_decap_4 FILLER_0_143_833 ();
 sg13g2_fill_2 FILLER_0_143_837 ();
 sg13g2_fill_1 FILLER_0_143_851 ();
 sg13g2_fill_1 FILLER_0_143_878 ();
 sg13g2_fill_1 FILLER_0_143_900 ();
 sg13g2_fill_2 FILLER_0_143_914 ();
 sg13g2_fill_1 FILLER_0_143_916 ();
 sg13g2_decap_8 FILLER_0_143_928 ();
 sg13g2_decap_4 FILLER_0_143_935 ();
 sg13g2_fill_1 FILLER_0_143_939 ();
 sg13g2_decap_8 FILLER_0_143_944 ();
 sg13g2_decap_8 FILLER_0_143_951 ();
 sg13g2_fill_1 FILLER_0_143_974 ();
 sg13g2_fill_2 FILLER_0_143_989 ();
 sg13g2_fill_2 FILLER_0_143_1026 ();
 sg13g2_fill_1 FILLER_0_143_1028 ();
 sg13g2_decap_8 FILLER_0_143_1046 ();
 sg13g2_decap_8 FILLER_0_143_1053 ();
 sg13g2_decap_8 FILLER_0_143_1060 ();
 sg13g2_decap_8 FILLER_0_143_1067 ();
 sg13g2_decap_8 FILLER_0_143_1074 ();
 sg13g2_decap_8 FILLER_0_143_1081 ();
 sg13g2_fill_1 FILLER_0_143_1088 ();
 sg13g2_decap_8 FILLER_0_143_1127 ();
 sg13g2_decap_8 FILLER_0_143_1134 ();
 sg13g2_decap_8 FILLER_0_143_1141 ();
 sg13g2_decap_8 FILLER_0_143_1148 ();
 sg13g2_decap_8 FILLER_0_143_1155 ();
 sg13g2_decap_8 FILLER_0_143_1162 ();
 sg13g2_decap_8 FILLER_0_143_1169 ();
 sg13g2_decap_8 FILLER_0_143_1176 ();
 sg13g2_decap_8 FILLER_0_143_1183 ();
 sg13g2_decap_8 FILLER_0_143_1190 ();
 sg13g2_decap_8 FILLER_0_143_1197 ();
 sg13g2_decap_8 FILLER_0_143_1204 ();
 sg13g2_decap_8 FILLER_0_143_1211 ();
 sg13g2_decap_8 FILLER_0_143_1218 ();
 sg13g2_fill_2 FILLER_0_143_1225 ();
 sg13g2_fill_1 FILLER_0_143_1227 ();
 sg13g2_fill_1 FILLER_0_144_0 ();
 sg13g2_fill_2 FILLER_0_144_70 ();
 sg13g2_fill_2 FILLER_0_144_76 ();
 sg13g2_decap_8 FILLER_0_144_83 ();
 sg13g2_decap_8 FILLER_0_144_90 ();
 sg13g2_fill_2 FILLER_0_144_101 ();
 sg13g2_fill_1 FILLER_0_144_103 ();
 sg13g2_fill_2 FILLER_0_144_109 ();
 sg13g2_fill_1 FILLER_0_144_111 ();
 sg13g2_decap_8 FILLER_0_144_142 ();
 sg13g2_decap_8 FILLER_0_144_149 ();
 sg13g2_decap_8 FILLER_0_144_156 ();
 sg13g2_decap_8 FILLER_0_144_163 ();
 sg13g2_decap_8 FILLER_0_144_170 ();
 sg13g2_decap_8 FILLER_0_144_177 ();
 sg13g2_decap_8 FILLER_0_144_184 ();
 sg13g2_decap_8 FILLER_0_144_191 ();
 sg13g2_decap_8 FILLER_0_144_198 ();
 sg13g2_decap_8 FILLER_0_144_205 ();
 sg13g2_decap_8 FILLER_0_144_212 ();
 sg13g2_decap_8 FILLER_0_144_219 ();
 sg13g2_decap_8 FILLER_0_144_226 ();
 sg13g2_decap_8 FILLER_0_144_233 ();
 sg13g2_decap_8 FILLER_0_144_240 ();
 sg13g2_decap_8 FILLER_0_144_247 ();
 sg13g2_decap_8 FILLER_0_144_254 ();
 sg13g2_decap_8 FILLER_0_144_261 ();
 sg13g2_decap_8 FILLER_0_144_268 ();
 sg13g2_decap_8 FILLER_0_144_275 ();
 sg13g2_decap_8 FILLER_0_144_282 ();
 sg13g2_decap_8 FILLER_0_144_289 ();
 sg13g2_decap_8 FILLER_0_144_296 ();
 sg13g2_decap_8 FILLER_0_144_303 ();
 sg13g2_decap_8 FILLER_0_144_310 ();
 sg13g2_decap_4 FILLER_0_144_317 ();
 sg13g2_decap_8 FILLER_0_144_325 ();
 sg13g2_fill_2 FILLER_0_144_332 ();
 sg13g2_fill_1 FILLER_0_144_334 ();
 sg13g2_decap_8 FILLER_0_144_371 ();
 sg13g2_decap_8 FILLER_0_144_378 ();
 sg13g2_decap_8 FILLER_0_144_385 ();
 sg13g2_decap_8 FILLER_0_144_392 ();
 sg13g2_decap_8 FILLER_0_144_399 ();
 sg13g2_decap_8 FILLER_0_144_406 ();
 sg13g2_decap_8 FILLER_0_144_413 ();
 sg13g2_decap_8 FILLER_0_144_420 ();
 sg13g2_decap_8 FILLER_0_144_427 ();
 sg13g2_decap_8 FILLER_0_144_434 ();
 sg13g2_decap_8 FILLER_0_144_441 ();
 sg13g2_decap_8 FILLER_0_144_448 ();
 sg13g2_decap_8 FILLER_0_144_455 ();
 sg13g2_decap_8 FILLER_0_144_462 ();
 sg13g2_decap_8 FILLER_0_144_469 ();
 sg13g2_decap_8 FILLER_0_144_476 ();
 sg13g2_decap_8 FILLER_0_144_483 ();
 sg13g2_decap_8 FILLER_0_144_490 ();
 sg13g2_decap_8 FILLER_0_144_497 ();
 sg13g2_decap_8 FILLER_0_144_504 ();
 sg13g2_decap_8 FILLER_0_144_511 ();
 sg13g2_decap_8 FILLER_0_144_518 ();
 sg13g2_decap_8 FILLER_0_144_525 ();
 sg13g2_decap_8 FILLER_0_144_532 ();
 sg13g2_decap_8 FILLER_0_144_539 ();
 sg13g2_decap_8 FILLER_0_144_546 ();
 sg13g2_decap_8 FILLER_0_144_553 ();
 sg13g2_decap_4 FILLER_0_144_560 ();
 sg13g2_decap_4 FILLER_0_144_590 ();
 sg13g2_fill_1 FILLER_0_144_594 ();
 sg13g2_fill_1 FILLER_0_144_605 ();
 sg13g2_fill_1 FILLER_0_144_621 ();
 sg13g2_decap_8 FILLER_0_144_648 ();
 sg13g2_decap_8 FILLER_0_144_655 ();
 sg13g2_fill_2 FILLER_0_144_662 ();
 sg13g2_fill_1 FILLER_0_144_664 ();
 sg13g2_fill_2 FILLER_0_144_691 ();
 sg13g2_fill_1 FILLER_0_144_719 ();
 sg13g2_fill_1 FILLER_0_144_753 ();
 sg13g2_fill_2 FILLER_0_144_796 ();
 sg13g2_fill_2 FILLER_0_144_803 ();
 sg13g2_fill_2 FILLER_0_144_820 ();
 sg13g2_fill_1 FILLER_0_144_822 ();
 sg13g2_decap_8 FILLER_0_144_828 ();
 sg13g2_decap_8 FILLER_0_144_835 ();
 sg13g2_decap_8 FILLER_0_144_842 ();
 sg13g2_fill_1 FILLER_0_144_849 ();
 sg13g2_fill_1 FILLER_0_144_863 ();
 sg13g2_fill_2 FILLER_0_144_869 ();
 sg13g2_decap_4 FILLER_0_144_901 ();
 sg13g2_fill_1 FILLER_0_144_914 ();
 sg13g2_fill_1 FILLER_0_144_926 ();
 sg13g2_fill_1 FILLER_0_144_944 ();
 sg13g2_decap_8 FILLER_0_144_959 ();
 sg13g2_fill_1 FILLER_0_144_1001 ();
 sg13g2_fill_1 FILLER_0_144_1007 ();
 sg13g2_fill_1 FILLER_0_144_1013 ();
 sg13g2_fill_1 FILLER_0_144_1025 ();
 sg13g2_fill_2 FILLER_0_144_1034 ();
 sg13g2_fill_1 FILLER_0_144_1044 ();
 sg13g2_decap_8 FILLER_0_144_1053 ();
 sg13g2_decap_8 FILLER_0_144_1060 ();
 sg13g2_decap_8 FILLER_0_144_1067 ();
 sg13g2_decap_8 FILLER_0_144_1074 ();
 sg13g2_decap_8 FILLER_0_144_1081 ();
 sg13g2_decap_8 FILLER_0_144_1088 ();
 sg13g2_fill_1 FILLER_0_144_1095 ();
 sg13g2_decap_8 FILLER_0_144_1137 ();
 sg13g2_decap_8 FILLER_0_144_1144 ();
 sg13g2_decap_8 FILLER_0_144_1151 ();
 sg13g2_decap_8 FILLER_0_144_1158 ();
 sg13g2_decap_8 FILLER_0_144_1165 ();
 sg13g2_decap_8 FILLER_0_144_1172 ();
 sg13g2_decap_8 FILLER_0_144_1179 ();
 sg13g2_decap_8 FILLER_0_144_1186 ();
 sg13g2_decap_8 FILLER_0_144_1193 ();
 sg13g2_decap_8 FILLER_0_144_1200 ();
 sg13g2_decap_8 FILLER_0_144_1207 ();
 sg13g2_decap_8 FILLER_0_144_1214 ();
 sg13g2_decap_8 FILLER_0_144_1221 ();
 sg13g2_decap_8 FILLER_0_145_0 ();
 sg13g2_decap_8 FILLER_0_145_7 ();
 sg13g2_decap_8 FILLER_0_145_14 ();
 sg13g2_fill_2 FILLER_0_145_21 ();
 sg13g2_fill_1 FILLER_0_145_23 ();
 sg13g2_fill_1 FILLER_0_145_47 ();
 sg13g2_decap_8 FILLER_0_145_57 ();
 sg13g2_fill_1 FILLER_0_145_64 ();
 sg13g2_decap_8 FILLER_0_145_69 ();
 sg13g2_decap_4 FILLER_0_145_76 ();
 sg13g2_decap_4 FILLER_0_145_85 ();
 sg13g2_fill_1 FILLER_0_145_89 ();
 sg13g2_fill_2 FILLER_0_145_116 ();
 sg13g2_decap_8 FILLER_0_145_127 ();
 sg13g2_decap_8 FILLER_0_145_134 ();
 sg13g2_decap_8 FILLER_0_145_141 ();
 sg13g2_decap_8 FILLER_0_145_148 ();
 sg13g2_decap_8 FILLER_0_145_155 ();
 sg13g2_decap_8 FILLER_0_145_162 ();
 sg13g2_decap_8 FILLER_0_145_169 ();
 sg13g2_decap_8 FILLER_0_145_176 ();
 sg13g2_decap_8 FILLER_0_145_183 ();
 sg13g2_decap_8 FILLER_0_145_190 ();
 sg13g2_decap_8 FILLER_0_145_197 ();
 sg13g2_decap_8 FILLER_0_145_204 ();
 sg13g2_decap_8 FILLER_0_145_211 ();
 sg13g2_decap_8 FILLER_0_145_218 ();
 sg13g2_decap_8 FILLER_0_145_225 ();
 sg13g2_decap_8 FILLER_0_145_232 ();
 sg13g2_decap_8 FILLER_0_145_239 ();
 sg13g2_decap_8 FILLER_0_145_246 ();
 sg13g2_decap_8 FILLER_0_145_253 ();
 sg13g2_decap_8 FILLER_0_145_260 ();
 sg13g2_decap_8 FILLER_0_145_267 ();
 sg13g2_decap_8 FILLER_0_145_274 ();
 sg13g2_decap_8 FILLER_0_145_281 ();
 sg13g2_decap_8 FILLER_0_145_288 ();
 sg13g2_decap_8 FILLER_0_145_295 ();
 sg13g2_decap_8 FILLER_0_145_302 ();
 sg13g2_decap_8 FILLER_0_145_309 ();
 sg13g2_decap_8 FILLER_0_145_316 ();
 sg13g2_decap_8 FILLER_0_145_323 ();
 sg13g2_decap_8 FILLER_0_145_330 ();
 sg13g2_decap_8 FILLER_0_145_337 ();
 sg13g2_decap_4 FILLER_0_145_344 ();
 sg13g2_decap_8 FILLER_0_145_352 ();
 sg13g2_decap_4 FILLER_0_145_359 ();
 sg13g2_decap_8 FILLER_0_145_367 ();
 sg13g2_decap_8 FILLER_0_145_374 ();
 sg13g2_decap_8 FILLER_0_145_381 ();
 sg13g2_decap_8 FILLER_0_145_388 ();
 sg13g2_decap_8 FILLER_0_145_395 ();
 sg13g2_decap_8 FILLER_0_145_402 ();
 sg13g2_decap_8 FILLER_0_145_409 ();
 sg13g2_decap_8 FILLER_0_145_416 ();
 sg13g2_decap_8 FILLER_0_145_423 ();
 sg13g2_decap_8 FILLER_0_145_430 ();
 sg13g2_decap_8 FILLER_0_145_437 ();
 sg13g2_decap_8 FILLER_0_145_444 ();
 sg13g2_decap_8 FILLER_0_145_451 ();
 sg13g2_decap_8 FILLER_0_145_458 ();
 sg13g2_decap_8 FILLER_0_145_465 ();
 sg13g2_decap_8 FILLER_0_145_472 ();
 sg13g2_decap_8 FILLER_0_145_479 ();
 sg13g2_decap_8 FILLER_0_145_486 ();
 sg13g2_decap_8 FILLER_0_145_493 ();
 sg13g2_decap_8 FILLER_0_145_500 ();
 sg13g2_decap_8 FILLER_0_145_507 ();
 sg13g2_decap_8 FILLER_0_145_514 ();
 sg13g2_decap_8 FILLER_0_145_521 ();
 sg13g2_decap_8 FILLER_0_145_528 ();
 sg13g2_decap_8 FILLER_0_145_535 ();
 sg13g2_decap_8 FILLER_0_145_542 ();
 sg13g2_decap_8 FILLER_0_145_549 ();
 sg13g2_decap_8 FILLER_0_145_556 ();
 sg13g2_decap_8 FILLER_0_145_563 ();
 sg13g2_decap_8 FILLER_0_145_570 ();
 sg13g2_decap_8 FILLER_0_145_577 ();
 sg13g2_decap_8 FILLER_0_145_584 ();
 sg13g2_decap_8 FILLER_0_145_591 ();
 sg13g2_decap_8 FILLER_0_145_598 ();
 sg13g2_decap_8 FILLER_0_145_605 ();
 sg13g2_decap_4 FILLER_0_145_612 ();
 sg13g2_decap_8 FILLER_0_145_644 ();
 sg13g2_decap_8 FILLER_0_145_651 ();
 sg13g2_decap_4 FILLER_0_145_658 ();
 sg13g2_fill_2 FILLER_0_145_662 ();
 sg13g2_fill_2 FILLER_0_145_673 ();
 sg13g2_decap_8 FILLER_0_145_685 ();
 sg13g2_decap_4 FILLER_0_145_697 ();
 sg13g2_decap_8 FILLER_0_145_705 ();
 sg13g2_fill_1 FILLER_0_145_712 ();
 sg13g2_fill_2 FILLER_0_145_744 ();
 sg13g2_fill_1 FILLER_0_145_789 ();
 sg13g2_fill_2 FILLER_0_145_799 ();
 sg13g2_fill_1 FILLER_0_145_840 ();
 sg13g2_decap_4 FILLER_0_145_846 ();
 sg13g2_fill_2 FILLER_0_145_854 ();
 sg13g2_fill_1 FILLER_0_145_860 ();
 sg13g2_fill_2 FILLER_0_145_871 ();
 sg13g2_fill_2 FILLER_0_145_878 ();
 sg13g2_fill_2 FILLER_0_145_886 ();
 sg13g2_fill_1 FILLER_0_145_897 ();
 sg13g2_decap_4 FILLER_0_145_908 ();
 sg13g2_fill_1 FILLER_0_145_912 ();
 sg13g2_fill_2 FILLER_0_145_918 ();
 sg13g2_fill_1 FILLER_0_145_934 ();
 sg13g2_fill_1 FILLER_0_145_946 ();
 sg13g2_decap_8 FILLER_0_145_952 ();
 sg13g2_decap_4 FILLER_0_145_959 ();
 sg13g2_fill_1 FILLER_0_145_963 ();
 sg13g2_fill_2 FILLER_0_145_971 ();
 sg13g2_fill_2 FILLER_0_145_1004 ();
 sg13g2_fill_1 FILLER_0_145_1014 ();
 sg13g2_decap_8 FILLER_0_145_1041 ();
 sg13g2_fill_2 FILLER_0_145_1048 ();
 sg13g2_fill_1 FILLER_0_145_1050 ();
 sg13g2_fill_2 FILLER_0_145_1070 ();
 sg13g2_fill_1 FILLER_0_145_1072 ();
 sg13g2_fill_2 FILLER_0_145_1099 ();
 sg13g2_fill_1 FILLER_0_145_1101 ();
 sg13g2_decap_4 FILLER_0_145_1112 ();
 sg13g2_fill_2 FILLER_0_145_1116 ();
 sg13g2_decap_8 FILLER_0_145_1122 ();
 sg13g2_decap_8 FILLER_0_145_1129 ();
 sg13g2_decap_8 FILLER_0_145_1136 ();
 sg13g2_decap_8 FILLER_0_145_1143 ();
 sg13g2_decap_8 FILLER_0_145_1150 ();
 sg13g2_decap_8 FILLER_0_145_1157 ();
 sg13g2_decap_8 FILLER_0_145_1164 ();
 sg13g2_decap_8 FILLER_0_145_1171 ();
 sg13g2_decap_8 FILLER_0_145_1178 ();
 sg13g2_decap_8 FILLER_0_145_1185 ();
 sg13g2_decap_8 FILLER_0_145_1192 ();
 sg13g2_decap_8 FILLER_0_145_1199 ();
 sg13g2_decap_8 FILLER_0_145_1206 ();
 sg13g2_decap_8 FILLER_0_145_1213 ();
 sg13g2_decap_8 FILLER_0_145_1220 ();
 sg13g2_fill_1 FILLER_0_145_1227 ();
 sg13g2_fill_1 FILLER_0_146_0 ();
 sg13g2_fill_1 FILLER_0_146_27 ();
 sg13g2_decap_4 FILLER_0_146_54 ();
 sg13g2_decap_8 FILLER_0_146_123 ();
 sg13g2_decap_8 FILLER_0_146_130 ();
 sg13g2_decap_8 FILLER_0_146_137 ();
 sg13g2_decap_8 FILLER_0_146_144 ();
 sg13g2_decap_8 FILLER_0_146_151 ();
 sg13g2_decap_8 FILLER_0_146_158 ();
 sg13g2_decap_8 FILLER_0_146_165 ();
 sg13g2_decap_8 FILLER_0_146_172 ();
 sg13g2_decap_8 FILLER_0_146_179 ();
 sg13g2_decap_8 FILLER_0_146_186 ();
 sg13g2_decap_8 FILLER_0_146_193 ();
 sg13g2_decap_8 FILLER_0_146_200 ();
 sg13g2_decap_8 FILLER_0_146_207 ();
 sg13g2_decap_8 FILLER_0_146_214 ();
 sg13g2_decap_8 FILLER_0_146_221 ();
 sg13g2_decap_8 FILLER_0_146_228 ();
 sg13g2_decap_8 FILLER_0_146_235 ();
 sg13g2_decap_8 FILLER_0_146_242 ();
 sg13g2_decap_8 FILLER_0_146_249 ();
 sg13g2_decap_8 FILLER_0_146_256 ();
 sg13g2_decap_8 FILLER_0_146_263 ();
 sg13g2_decap_8 FILLER_0_146_270 ();
 sg13g2_decap_8 FILLER_0_146_277 ();
 sg13g2_decap_8 FILLER_0_146_284 ();
 sg13g2_decap_8 FILLER_0_146_291 ();
 sg13g2_decap_8 FILLER_0_146_298 ();
 sg13g2_decap_8 FILLER_0_146_305 ();
 sg13g2_decap_8 FILLER_0_146_312 ();
 sg13g2_decap_8 FILLER_0_146_319 ();
 sg13g2_decap_8 FILLER_0_146_326 ();
 sg13g2_decap_8 FILLER_0_146_333 ();
 sg13g2_decap_8 FILLER_0_146_340 ();
 sg13g2_decap_8 FILLER_0_146_347 ();
 sg13g2_decap_8 FILLER_0_146_354 ();
 sg13g2_decap_8 FILLER_0_146_361 ();
 sg13g2_decap_8 FILLER_0_146_368 ();
 sg13g2_decap_8 FILLER_0_146_375 ();
 sg13g2_decap_8 FILLER_0_146_382 ();
 sg13g2_decap_8 FILLER_0_146_389 ();
 sg13g2_decap_8 FILLER_0_146_396 ();
 sg13g2_decap_8 FILLER_0_146_403 ();
 sg13g2_decap_8 FILLER_0_146_410 ();
 sg13g2_decap_8 FILLER_0_146_417 ();
 sg13g2_decap_8 FILLER_0_146_424 ();
 sg13g2_decap_8 FILLER_0_146_431 ();
 sg13g2_decap_8 FILLER_0_146_438 ();
 sg13g2_decap_8 FILLER_0_146_445 ();
 sg13g2_decap_8 FILLER_0_146_452 ();
 sg13g2_decap_8 FILLER_0_146_459 ();
 sg13g2_decap_8 FILLER_0_146_466 ();
 sg13g2_decap_8 FILLER_0_146_473 ();
 sg13g2_decap_8 FILLER_0_146_480 ();
 sg13g2_decap_8 FILLER_0_146_487 ();
 sg13g2_decap_8 FILLER_0_146_494 ();
 sg13g2_decap_8 FILLER_0_146_501 ();
 sg13g2_decap_8 FILLER_0_146_508 ();
 sg13g2_decap_8 FILLER_0_146_515 ();
 sg13g2_decap_8 FILLER_0_146_522 ();
 sg13g2_decap_8 FILLER_0_146_529 ();
 sg13g2_decap_8 FILLER_0_146_536 ();
 sg13g2_decap_8 FILLER_0_146_543 ();
 sg13g2_decap_8 FILLER_0_146_550 ();
 sg13g2_decap_8 FILLER_0_146_557 ();
 sg13g2_decap_8 FILLER_0_146_564 ();
 sg13g2_decap_8 FILLER_0_146_571 ();
 sg13g2_decap_8 FILLER_0_146_578 ();
 sg13g2_decap_8 FILLER_0_146_585 ();
 sg13g2_decap_8 FILLER_0_146_592 ();
 sg13g2_decap_8 FILLER_0_146_599 ();
 sg13g2_decap_8 FILLER_0_146_606 ();
 sg13g2_decap_4 FILLER_0_146_613 ();
 sg13g2_fill_1 FILLER_0_146_617 ();
 sg13g2_fill_2 FILLER_0_146_653 ();
 sg13g2_decap_8 FILLER_0_146_686 ();
 sg13g2_decap_8 FILLER_0_146_693 ();
 sg13g2_decap_8 FILLER_0_146_700 ();
 sg13g2_decap_8 FILLER_0_146_707 ();
 sg13g2_fill_1 FILLER_0_146_714 ();
 sg13g2_decap_4 FILLER_0_146_720 ();
 sg13g2_fill_1 FILLER_0_146_724 ();
 sg13g2_decap_4 FILLER_0_146_729 ();
 sg13g2_fill_1 FILLER_0_146_733 ();
 sg13g2_fill_1 FILLER_0_146_757 ();
 sg13g2_fill_1 FILLER_0_146_784 ();
 sg13g2_fill_2 FILLER_0_146_808 ();
 sg13g2_fill_1 FILLER_0_146_810 ();
 sg13g2_fill_2 FILLER_0_146_824 ();
 sg13g2_fill_1 FILLER_0_146_854 ();
 sg13g2_decap_4 FILLER_0_146_865 ();
 sg13g2_fill_1 FILLER_0_146_869 ();
 sg13g2_fill_2 FILLER_0_146_875 ();
 sg13g2_decap_4 FILLER_0_146_882 ();
 sg13g2_fill_1 FILLER_0_146_894 ();
 sg13g2_fill_1 FILLER_0_146_903 ();
 sg13g2_fill_1 FILLER_0_146_911 ();
 sg13g2_decap_4 FILLER_0_146_950 ();
 sg13g2_fill_2 FILLER_0_146_954 ();
 sg13g2_fill_1 FILLER_0_146_993 ();
 sg13g2_fill_2 FILLER_0_146_1002 ();
 sg13g2_fill_2 FILLER_0_146_1009 ();
 sg13g2_fill_2 FILLER_0_146_1016 ();
 sg13g2_fill_1 FILLER_0_146_1018 ();
 sg13g2_decap_8 FILLER_0_146_1030 ();
 sg13g2_decap_4 FILLER_0_146_1037 ();
 sg13g2_fill_2 FILLER_0_146_1041 ();
 sg13g2_fill_1 FILLER_0_146_1048 ();
 sg13g2_fill_2 FILLER_0_146_1075 ();
 sg13g2_fill_2 FILLER_0_146_1081 ();
 sg13g2_fill_2 FILLER_0_146_1109 ();
 sg13g2_fill_2 FILLER_0_146_1116 ();
 sg13g2_fill_1 FILLER_0_146_1118 ();
 sg13g2_decap_8 FILLER_0_146_1145 ();
 sg13g2_decap_8 FILLER_0_146_1152 ();
 sg13g2_decap_8 FILLER_0_146_1159 ();
 sg13g2_decap_8 FILLER_0_146_1166 ();
 sg13g2_decap_8 FILLER_0_146_1173 ();
 sg13g2_decap_8 FILLER_0_146_1180 ();
 sg13g2_decap_8 FILLER_0_146_1187 ();
 sg13g2_decap_8 FILLER_0_146_1194 ();
 sg13g2_decap_8 FILLER_0_146_1201 ();
 sg13g2_decap_8 FILLER_0_146_1208 ();
 sg13g2_decap_8 FILLER_0_146_1215 ();
 sg13g2_decap_4 FILLER_0_146_1222 ();
 sg13g2_fill_2 FILLER_0_146_1226 ();
 sg13g2_decap_8 FILLER_0_147_0 ();
 sg13g2_decap_4 FILLER_0_147_11 ();
 sg13g2_fill_1 FILLER_0_147_15 ();
 sg13g2_decap_8 FILLER_0_147_21 ();
 sg13g2_decap_8 FILLER_0_147_141 ();
 sg13g2_decap_8 FILLER_0_147_148 ();
 sg13g2_decap_8 FILLER_0_147_155 ();
 sg13g2_decap_8 FILLER_0_147_162 ();
 sg13g2_decap_8 FILLER_0_147_169 ();
 sg13g2_decap_8 FILLER_0_147_176 ();
 sg13g2_decap_8 FILLER_0_147_183 ();
 sg13g2_decap_8 FILLER_0_147_190 ();
 sg13g2_decap_8 FILLER_0_147_197 ();
 sg13g2_decap_8 FILLER_0_147_204 ();
 sg13g2_decap_8 FILLER_0_147_211 ();
 sg13g2_decap_8 FILLER_0_147_218 ();
 sg13g2_decap_8 FILLER_0_147_225 ();
 sg13g2_decap_8 FILLER_0_147_232 ();
 sg13g2_decap_8 FILLER_0_147_239 ();
 sg13g2_decap_8 FILLER_0_147_246 ();
 sg13g2_decap_8 FILLER_0_147_253 ();
 sg13g2_decap_8 FILLER_0_147_260 ();
 sg13g2_decap_8 FILLER_0_147_267 ();
 sg13g2_decap_8 FILLER_0_147_274 ();
 sg13g2_decap_8 FILLER_0_147_281 ();
 sg13g2_decap_8 FILLER_0_147_288 ();
 sg13g2_decap_8 FILLER_0_147_295 ();
 sg13g2_decap_8 FILLER_0_147_302 ();
 sg13g2_decap_8 FILLER_0_147_309 ();
 sg13g2_decap_8 FILLER_0_147_316 ();
 sg13g2_decap_8 FILLER_0_147_323 ();
 sg13g2_decap_8 FILLER_0_147_330 ();
 sg13g2_decap_8 FILLER_0_147_337 ();
 sg13g2_decap_8 FILLER_0_147_344 ();
 sg13g2_decap_8 FILLER_0_147_351 ();
 sg13g2_decap_8 FILLER_0_147_358 ();
 sg13g2_decap_8 FILLER_0_147_365 ();
 sg13g2_decap_8 FILLER_0_147_372 ();
 sg13g2_decap_8 FILLER_0_147_379 ();
 sg13g2_decap_8 FILLER_0_147_386 ();
 sg13g2_decap_8 FILLER_0_147_393 ();
 sg13g2_decap_8 FILLER_0_147_400 ();
 sg13g2_decap_8 FILLER_0_147_407 ();
 sg13g2_decap_8 FILLER_0_147_414 ();
 sg13g2_decap_8 FILLER_0_147_421 ();
 sg13g2_decap_8 FILLER_0_147_428 ();
 sg13g2_decap_8 FILLER_0_147_435 ();
 sg13g2_decap_8 FILLER_0_147_442 ();
 sg13g2_decap_8 FILLER_0_147_449 ();
 sg13g2_decap_8 FILLER_0_147_456 ();
 sg13g2_decap_8 FILLER_0_147_463 ();
 sg13g2_decap_8 FILLER_0_147_470 ();
 sg13g2_decap_8 FILLER_0_147_477 ();
 sg13g2_decap_8 FILLER_0_147_484 ();
 sg13g2_decap_8 FILLER_0_147_491 ();
 sg13g2_decap_8 FILLER_0_147_498 ();
 sg13g2_decap_8 FILLER_0_147_505 ();
 sg13g2_decap_8 FILLER_0_147_512 ();
 sg13g2_decap_8 FILLER_0_147_519 ();
 sg13g2_decap_8 FILLER_0_147_526 ();
 sg13g2_decap_8 FILLER_0_147_533 ();
 sg13g2_decap_8 FILLER_0_147_540 ();
 sg13g2_decap_8 FILLER_0_147_547 ();
 sg13g2_decap_8 FILLER_0_147_554 ();
 sg13g2_decap_8 FILLER_0_147_561 ();
 sg13g2_decap_8 FILLER_0_147_568 ();
 sg13g2_decap_8 FILLER_0_147_575 ();
 sg13g2_decap_8 FILLER_0_147_582 ();
 sg13g2_decap_8 FILLER_0_147_589 ();
 sg13g2_decap_8 FILLER_0_147_596 ();
 sg13g2_decap_8 FILLER_0_147_603 ();
 sg13g2_decap_8 FILLER_0_147_610 ();
 sg13g2_fill_2 FILLER_0_147_617 ();
 sg13g2_fill_1 FILLER_0_147_619 ();
 sg13g2_decap_8 FILLER_0_147_650 ();
 sg13g2_fill_1 FILLER_0_147_657 ();
 sg13g2_decap_4 FILLER_0_147_662 ();
 sg13g2_fill_1 FILLER_0_147_666 ();
 sg13g2_decap_4 FILLER_0_147_671 ();
 sg13g2_fill_1 FILLER_0_147_675 ();
 sg13g2_decap_8 FILLER_0_147_686 ();
 sg13g2_fill_2 FILLER_0_147_693 ();
 sg13g2_decap_8 FILLER_0_147_705 ();
 sg13g2_decap_8 FILLER_0_147_712 ();
 sg13g2_decap_8 FILLER_0_147_719 ();
 sg13g2_decap_4 FILLER_0_147_726 ();
 sg13g2_fill_2 FILLER_0_147_730 ();
 sg13g2_decap_8 FILLER_0_147_776 ();
 sg13g2_fill_1 FILLER_0_147_783 ();
 sg13g2_fill_2 FILLER_0_147_815 ();
 sg13g2_fill_1 FILLER_0_147_827 ();
 sg13g2_fill_1 FILLER_0_147_832 ();
 sg13g2_fill_1 FILLER_0_147_846 ();
 sg13g2_fill_1 FILLER_0_147_852 ();
 sg13g2_fill_1 FILLER_0_147_879 ();
 sg13g2_fill_2 FILLER_0_147_885 ();
 sg13g2_fill_2 FILLER_0_147_896 ();
 sg13g2_fill_2 FILLER_0_147_909 ();
 sg13g2_fill_1 FILLER_0_147_916 ();
 sg13g2_decap_4 FILLER_0_147_922 ();
 sg13g2_fill_1 FILLER_0_147_926 ();
 sg13g2_fill_1 FILLER_0_147_932 ();
 sg13g2_fill_2 FILLER_0_147_937 ();
 sg13g2_fill_1 FILLER_0_147_944 ();
 sg13g2_decap_8 FILLER_0_147_950 ();
 sg13g2_fill_1 FILLER_0_147_957 ();
 sg13g2_decap_8 FILLER_0_147_967 ();
 sg13g2_fill_2 FILLER_0_147_974 ();
 sg13g2_decap_4 FILLER_0_147_981 ();
 sg13g2_fill_1 FILLER_0_147_985 ();
 sg13g2_decap_8 FILLER_0_147_990 ();
 sg13g2_decap_8 FILLER_0_147_997 ();
 sg13g2_decap_8 FILLER_0_147_1004 ();
 sg13g2_decap_8 FILLER_0_147_1011 ();
 sg13g2_decap_8 FILLER_0_147_1018 ();
 sg13g2_decap_4 FILLER_0_147_1025 ();
 sg13g2_fill_1 FILLER_0_147_1029 ();
 sg13g2_fill_1 FILLER_0_147_1061 ();
 sg13g2_fill_2 FILLER_0_147_1072 ();
 sg13g2_fill_2 FILLER_0_147_1084 ();
 sg13g2_fill_1 FILLER_0_147_1086 ();
 sg13g2_fill_2 FILLER_0_147_1097 ();
 sg13g2_fill_1 FILLER_0_147_1099 ();
 sg13g2_fill_2 FILLER_0_147_1126 ();
 sg13g2_fill_1 FILLER_0_147_1128 ();
 sg13g2_decap_8 FILLER_0_147_1133 ();
 sg13g2_decap_8 FILLER_0_147_1140 ();
 sg13g2_decap_8 FILLER_0_147_1147 ();
 sg13g2_decap_8 FILLER_0_147_1154 ();
 sg13g2_decap_8 FILLER_0_147_1161 ();
 sg13g2_decap_8 FILLER_0_147_1168 ();
 sg13g2_decap_8 FILLER_0_147_1175 ();
 sg13g2_decap_8 FILLER_0_147_1182 ();
 sg13g2_decap_8 FILLER_0_147_1189 ();
 sg13g2_decap_8 FILLER_0_147_1196 ();
 sg13g2_decap_8 FILLER_0_147_1203 ();
 sg13g2_decap_8 FILLER_0_147_1210 ();
 sg13g2_decap_8 FILLER_0_147_1217 ();
 sg13g2_decap_4 FILLER_0_147_1224 ();
 sg13g2_decap_8 FILLER_0_148_0 ();
 sg13g2_fill_2 FILLER_0_148_7 ();
 sg13g2_fill_1 FILLER_0_148_9 ();
 sg13g2_fill_1 FILLER_0_148_14 ();
 sg13g2_fill_2 FILLER_0_148_44 ();
 sg13g2_fill_1 FILLER_0_148_51 ();
 sg13g2_fill_2 FILLER_0_148_78 ();
 sg13g2_fill_1 FILLER_0_148_85 ();
 sg13g2_fill_2 FILLER_0_148_100 ();
 sg13g2_fill_1 FILLER_0_148_102 ();
 sg13g2_fill_2 FILLER_0_148_111 ();
 sg13g2_fill_2 FILLER_0_148_118 ();
 sg13g2_fill_1 FILLER_0_148_120 ();
 sg13g2_fill_2 FILLER_0_148_125 ();
 sg13g2_decap_8 FILLER_0_148_131 ();
 sg13g2_decap_8 FILLER_0_148_138 ();
 sg13g2_decap_8 FILLER_0_148_145 ();
 sg13g2_decap_8 FILLER_0_148_152 ();
 sg13g2_decap_8 FILLER_0_148_159 ();
 sg13g2_decap_8 FILLER_0_148_166 ();
 sg13g2_decap_8 FILLER_0_148_173 ();
 sg13g2_decap_8 FILLER_0_148_180 ();
 sg13g2_decap_8 FILLER_0_148_187 ();
 sg13g2_decap_8 FILLER_0_148_194 ();
 sg13g2_decap_8 FILLER_0_148_201 ();
 sg13g2_decap_8 FILLER_0_148_208 ();
 sg13g2_decap_8 FILLER_0_148_215 ();
 sg13g2_decap_8 FILLER_0_148_222 ();
 sg13g2_decap_8 FILLER_0_148_229 ();
 sg13g2_decap_8 FILLER_0_148_236 ();
 sg13g2_decap_8 FILLER_0_148_243 ();
 sg13g2_decap_8 FILLER_0_148_250 ();
 sg13g2_decap_8 FILLER_0_148_257 ();
 sg13g2_decap_8 FILLER_0_148_264 ();
 sg13g2_decap_8 FILLER_0_148_271 ();
 sg13g2_decap_8 FILLER_0_148_278 ();
 sg13g2_decap_8 FILLER_0_148_285 ();
 sg13g2_decap_8 FILLER_0_148_292 ();
 sg13g2_decap_8 FILLER_0_148_299 ();
 sg13g2_decap_8 FILLER_0_148_306 ();
 sg13g2_decap_8 FILLER_0_148_313 ();
 sg13g2_decap_8 FILLER_0_148_320 ();
 sg13g2_decap_8 FILLER_0_148_327 ();
 sg13g2_decap_8 FILLER_0_148_334 ();
 sg13g2_decap_8 FILLER_0_148_341 ();
 sg13g2_decap_8 FILLER_0_148_348 ();
 sg13g2_decap_8 FILLER_0_148_355 ();
 sg13g2_decap_8 FILLER_0_148_362 ();
 sg13g2_decap_8 FILLER_0_148_369 ();
 sg13g2_decap_8 FILLER_0_148_376 ();
 sg13g2_decap_8 FILLER_0_148_383 ();
 sg13g2_decap_8 FILLER_0_148_390 ();
 sg13g2_decap_8 FILLER_0_148_397 ();
 sg13g2_decap_8 FILLER_0_148_404 ();
 sg13g2_decap_8 FILLER_0_148_411 ();
 sg13g2_decap_8 FILLER_0_148_418 ();
 sg13g2_decap_8 FILLER_0_148_425 ();
 sg13g2_decap_8 FILLER_0_148_432 ();
 sg13g2_decap_8 FILLER_0_148_439 ();
 sg13g2_decap_8 FILLER_0_148_446 ();
 sg13g2_decap_8 FILLER_0_148_453 ();
 sg13g2_decap_8 FILLER_0_148_460 ();
 sg13g2_decap_8 FILLER_0_148_467 ();
 sg13g2_decap_8 FILLER_0_148_474 ();
 sg13g2_decap_8 FILLER_0_148_481 ();
 sg13g2_decap_8 FILLER_0_148_488 ();
 sg13g2_decap_8 FILLER_0_148_495 ();
 sg13g2_decap_8 FILLER_0_148_502 ();
 sg13g2_decap_8 FILLER_0_148_509 ();
 sg13g2_decap_8 FILLER_0_148_516 ();
 sg13g2_decap_8 FILLER_0_148_523 ();
 sg13g2_decap_8 FILLER_0_148_530 ();
 sg13g2_decap_8 FILLER_0_148_537 ();
 sg13g2_decap_8 FILLER_0_148_544 ();
 sg13g2_decap_8 FILLER_0_148_551 ();
 sg13g2_decap_8 FILLER_0_148_558 ();
 sg13g2_decap_8 FILLER_0_148_565 ();
 sg13g2_decap_8 FILLER_0_148_572 ();
 sg13g2_decap_8 FILLER_0_148_579 ();
 sg13g2_decap_8 FILLER_0_148_586 ();
 sg13g2_decap_8 FILLER_0_148_593 ();
 sg13g2_decap_8 FILLER_0_148_600 ();
 sg13g2_decap_8 FILLER_0_148_607 ();
 sg13g2_decap_8 FILLER_0_148_614 ();
 sg13g2_fill_1 FILLER_0_148_621 ();
 sg13g2_fill_2 FILLER_0_148_648 ();
 sg13g2_fill_1 FILLER_0_148_650 ();
 sg13g2_fill_1 FILLER_0_148_729 ();
 sg13g2_fill_2 FILLER_0_148_748 ();
 sg13g2_fill_2 FILLER_0_148_753 ();
 sg13g2_decap_4 FILLER_0_148_776 ();
 sg13g2_fill_1 FILLER_0_148_790 ();
 sg13g2_fill_2 FILLER_0_148_831 ();
 sg13g2_fill_1 FILLER_0_148_843 ();
 sg13g2_fill_1 FILLER_0_148_849 ();
 sg13g2_fill_1 FILLER_0_148_860 ();
 sg13g2_fill_1 FILLER_0_148_887 ();
 sg13g2_fill_1 FILLER_0_148_892 ();
 sg13g2_fill_2 FILLER_0_148_897 ();
 sg13g2_decap_4 FILLER_0_148_908 ();
 sg13g2_fill_1 FILLER_0_148_912 ();
 sg13g2_fill_1 FILLER_0_148_918 ();
 sg13g2_fill_2 FILLER_0_148_935 ();
 sg13g2_fill_1 FILLER_0_148_937 ();
 sg13g2_fill_1 FILLER_0_148_942 ();
 sg13g2_fill_1 FILLER_0_148_947 ();
 sg13g2_decap_8 FILLER_0_148_974 ();
 sg13g2_decap_8 FILLER_0_148_981 ();
 sg13g2_decap_8 FILLER_0_148_988 ();
 sg13g2_decap_8 FILLER_0_148_995 ();
 sg13g2_decap_8 FILLER_0_148_1006 ();
 sg13g2_fill_2 FILLER_0_148_1013 ();
 sg13g2_fill_2 FILLER_0_148_1018 ();
 sg13g2_fill_1 FILLER_0_148_1020 ();
 sg13g2_fill_1 FILLER_0_148_1045 ();
 sg13g2_fill_2 FILLER_0_148_1072 ();
 sg13g2_fill_1 FILLER_0_148_1074 ();
 sg13g2_fill_2 FILLER_0_148_1089 ();
 sg13g2_decap_8 FILLER_0_148_1115 ();
 sg13g2_decap_8 FILLER_0_148_1122 ();
 sg13g2_decap_8 FILLER_0_148_1129 ();
 sg13g2_decap_8 FILLER_0_148_1136 ();
 sg13g2_decap_8 FILLER_0_148_1143 ();
 sg13g2_decap_8 FILLER_0_148_1150 ();
 sg13g2_decap_8 FILLER_0_148_1157 ();
 sg13g2_decap_8 FILLER_0_148_1164 ();
 sg13g2_decap_8 FILLER_0_148_1171 ();
 sg13g2_decap_8 FILLER_0_148_1178 ();
 sg13g2_decap_8 FILLER_0_148_1185 ();
 sg13g2_decap_8 FILLER_0_148_1192 ();
 sg13g2_decap_8 FILLER_0_148_1199 ();
 sg13g2_decap_8 FILLER_0_148_1206 ();
 sg13g2_decap_8 FILLER_0_148_1213 ();
 sg13g2_decap_8 FILLER_0_148_1220 ();
 sg13g2_fill_1 FILLER_0_148_1227 ();
 sg13g2_decap_4 FILLER_0_149_0 ();
 sg13g2_fill_1 FILLER_0_149_48 ();
 sg13g2_fill_1 FILLER_0_149_53 ();
 sg13g2_fill_1 FILLER_0_149_59 ();
 sg13g2_fill_2 FILLER_0_149_64 ();
 sg13g2_fill_1 FILLER_0_149_74 ();
 sg13g2_decap_8 FILLER_0_149_80 ();
 sg13g2_decap_8 FILLER_0_149_87 ();
 sg13g2_decap_8 FILLER_0_149_94 ();
 sg13g2_decap_8 FILLER_0_149_101 ();
 sg13g2_decap_4 FILLER_0_149_108 ();
 sg13g2_fill_2 FILLER_0_149_112 ();
 sg13g2_decap_8 FILLER_0_149_140 ();
 sg13g2_decap_8 FILLER_0_149_147 ();
 sg13g2_decap_8 FILLER_0_149_154 ();
 sg13g2_decap_8 FILLER_0_149_161 ();
 sg13g2_decap_8 FILLER_0_149_168 ();
 sg13g2_decap_8 FILLER_0_149_175 ();
 sg13g2_decap_8 FILLER_0_149_182 ();
 sg13g2_decap_8 FILLER_0_149_189 ();
 sg13g2_decap_8 FILLER_0_149_196 ();
 sg13g2_decap_8 FILLER_0_149_203 ();
 sg13g2_decap_8 FILLER_0_149_210 ();
 sg13g2_decap_8 FILLER_0_149_217 ();
 sg13g2_decap_8 FILLER_0_149_224 ();
 sg13g2_decap_8 FILLER_0_149_231 ();
 sg13g2_decap_8 FILLER_0_149_238 ();
 sg13g2_decap_8 FILLER_0_149_245 ();
 sg13g2_decap_8 FILLER_0_149_252 ();
 sg13g2_decap_8 FILLER_0_149_259 ();
 sg13g2_decap_8 FILLER_0_149_266 ();
 sg13g2_decap_8 FILLER_0_149_273 ();
 sg13g2_decap_8 FILLER_0_149_280 ();
 sg13g2_decap_8 FILLER_0_149_287 ();
 sg13g2_decap_8 FILLER_0_149_294 ();
 sg13g2_decap_8 FILLER_0_149_301 ();
 sg13g2_decap_8 FILLER_0_149_308 ();
 sg13g2_decap_8 FILLER_0_149_315 ();
 sg13g2_decap_8 FILLER_0_149_322 ();
 sg13g2_decap_8 FILLER_0_149_329 ();
 sg13g2_decap_8 FILLER_0_149_336 ();
 sg13g2_decap_8 FILLER_0_149_343 ();
 sg13g2_decap_8 FILLER_0_149_350 ();
 sg13g2_decap_8 FILLER_0_149_357 ();
 sg13g2_decap_8 FILLER_0_149_364 ();
 sg13g2_decap_8 FILLER_0_149_371 ();
 sg13g2_decap_8 FILLER_0_149_378 ();
 sg13g2_decap_8 FILLER_0_149_385 ();
 sg13g2_decap_8 FILLER_0_149_392 ();
 sg13g2_decap_8 FILLER_0_149_399 ();
 sg13g2_decap_8 FILLER_0_149_406 ();
 sg13g2_decap_8 FILLER_0_149_413 ();
 sg13g2_decap_8 FILLER_0_149_420 ();
 sg13g2_decap_8 FILLER_0_149_427 ();
 sg13g2_decap_8 FILLER_0_149_434 ();
 sg13g2_decap_8 FILLER_0_149_441 ();
 sg13g2_decap_8 FILLER_0_149_448 ();
 sg13g2_decap_8 FILLER_0_149_455 ();
 sg13g2_decap_8 FILLER_0_149_462 ();
 sg13g2_decap_8 FILLER_0_149_469 ();
 sg13g2_decap_8 FILLER_0_149_476 ();
 sg13g2_decap_8 FILLER_0_149_483 ();
 sg13g2_decap_8 FILLER_0_149_490 ();
 sg13g2_decap_8 FILLER_0_149_497 ();
 sg13g2_decap_8 FILLER_0_149_504 ();
 sg13g2_decap_8 FILLER_0_149_511 ();
 sg13g2_decap_8 FILLER_0_149_518 ();
 sg13g2_decap_8 FILLER_0_149_525 ();
 sg13g2_decap_8 FILLER_0_149_532 ();
 sg13g2_decap_8 FILLER_0_149_539 ();
 sg13g2_decap_8 FILLER_0_149_546 ();
 sg13g2_decap_8 FILLER_0_149_553 ();
 sg13g2_decap_8 FILLER_0_149_560 ();
 sg13g2_decap_8 FILLER_0_149_567 ();
 sg13g2_decap_8 FILLER_0_149_574 ();
 sg13g2_decap_8 FILLER_0_149_581 ();
 sg13g2_decap_8 FILLER_0_149_588 ();
 sg13g2_decap_8 FILLER_0_149_595 ();
 sg13g2_decap_8 FILLER_0_149_602 ();
 sg13g2_decap_8 FILLER_0_149_609 ();
 sg13g2_decap_8 FILLER_0_149_616 ();
 sg13g2_decap_8 FILLER_0_149_623 ();
 sg13g2_decap_8 FILLER_0_149_630 ();
 sg13g2_decap_4 FILLER_0_149_637 ();
 sg13g2_fill_1 FILLER_0_149_641 ();
 sg13g2_decap_4 FILLER_0_149_662 ();
 sg13g2_fill_2 FILLER_0_149_684 ();
 sg13g2_fill_1 FILLER_0_149_686 ();
 sg13g2_fill_2 FILLER_0_149_691 ();
 sg13g2_fill_1 FILLER_0_149_693 ();
 sg13g2_fill_2 FILLER_0_149_699 ();
 sg13g2_fill_1 FILLER_0_149_701 ();
 sg13g2_decap_8 FILLER_0_149_721 ();
 sg13g2_decap_4 FILLER_0_149_728 ();
 sg13g2_fill_2 FILLER_0_149_736 ();
 sg13g2_fill_2 FILLER_0_149_760 ();
 sg13g2_fill_1 FILLER_0_149_762 ();
 sg13g2_fill_2 FILLER_0_149_797 ();
 sg13g2_fill_2 FILLER_0_149_803 ();
 sg13g2_fill_2 FILLER_0_149_809 ();
 sg13g2_fill_1 FILLER_0_149_816 ();
 sg13g2_fill_1 FILLER_0_149_843 ();
 sg13g2_fill_1 FILLER_0_149_853 ();
 sg13g2_fill_1 FILLER_0_149_864 ();
 sg13g2_fill_1 FILLER_0_149_869 ();
 sg13g2_fill_2 FILLER_0_149_874 ();
 sg13g2_decap_4 FILLER_0_149_881 ();
 sg13g2_fill_1 FILLER_0_149_885 ();
 sg13g2_fill_2 FILLER_0_149_895 ();
 sg13g2_fill_1 FILLER_0_149_897 ();
 sg13g2_fill_2 FILLER_0_149_903 ();
 sg13g2_decap_4 FILLER_0_149_908 ();
 sg13g2_decap_4 FILLER_0_149_917 ();
 sg13g2_fill_2 FILLER_0_149_931 ();
 sg13g2_fill_1 FILLER_0_149_933 ();
 sg13g2_decap_4 FILLER_0_149_938 ();
 sg13g2_fill_1 FILLER_0_149_947 ();
 sg13g2_decap_8 FILLER_0_149_983 ();
 sg13g2_decap_4 FILLER_0_149_990 ();
 sg13g2_fill_2 FILLER_0_149_994 ();
 sg13g2_fill_2 FILLER_0_149_1001 ();
 sg13g2_fill_1 FILLER_0_149_1003 ();
 sg13g2_fill_1 FILLER_0_149_1014 ();
 sg13g2_decap_8 FILLER_0_149_1046 ();
 sg13g2_fill_1 FILLER_0_149_1053 ();
 sg13g2_decap_8 FILLER_0_149_1058 ();
 sg13g2_decap_8 FILLER_0_149_1065 ();
 sg13g2_decap_8 FILLER_0_149_1072 ();
 sg13g2_fill_2 FILLER_0_149_1079 ();
 sg13g2_fill_1 FILLER_0_149_1081 ();
 sg13g2_decap_8 FILLER_0_149_1132 ();
 sg13g2_decap_8 FILLER_0_149_1139 ();
 sg13g2_decap_8 FILLER_0_149_1146 ();
 sg13g2_decap_8 FILLER_0_149_1153 ();
 sg13g2_decap_8 FILLER_0_149_1160 ();
 sg13g2_decap_8 FILLER_0_149_1167 ();
 sg13g2_decap_8 FILLER_0_149_1174 ();
 sg13g2_decap_8 FILLER_0_149_1181 ();
 sg13g2_decap_8 FILLER_0_149_1188 ();
 sg13g2_decap_8 FILLER_0_149_1195 ();
 sg13g2_decap_8 FILLER_0_149_1202 ();
 sg13g2_decap_8 FILLER_0_149_1209 ();
 sg13g2_decap_8 FILLER_0_149_1216 ();
 sg13g2_decap_4 FILLER_0_149_1223 ();
 sg13g2_fill_1 FILLER_0_149_1227 ();
 sg13g2_fill_1 FILLER_0_150_43 ();
 sg13g2_decap_8 FILLER_0_150_53 ();
 sg13g2_decap_8 FILLER_0_150_76 ();
 sg13g2_fill_1 FILLER_0_150_83 ();
 sg13g2_decap_8 FILLER_0_150_88 ();
 sg13g2_decap_8 FILLER_0_150_95 ();
 sg13g2_fill_2 FILLER_0_150_102 ();
 sg13g2_fill_1 FILLER_0_150_104 ();
 sg13g2_decap_8 FILLER_0_150_140 ();
 sg13g2_decap_8 FILLER_0_150_147 ();
 sg13g2_decap_8 FILLER_0_150_154 ();
 sg13g2_decap_8 FILLER_0_150_161 ();
 sg13g2_decap_8 FILLER_0_150_168 ();
 sg13g2_decap_8 FILLER_0_150_175 ();
 sg13g2_decap_8 FILLER_0_150_182 ();
 sg13g2_decap_8 FILLER_0_150_189 ();
 sg13g2_decap_8 FILLER_0_150_196 ();
 sg13g2_decap_8 FILLER_0_150_203 ();
 sg13g2_decap_8 FILLER_0_150_210 ();
 sg13g2_decap_8 FILLER_0_150_217 ();
 sg13g2_decap_8 FILLER_0_150_224 ();
 sg13g2_decap_8 FILLER_0_150_231 ();
 sg13g2_decap_8 FILLER_0_150_238 ();
 sg13g2_decap_8 FILLER_0_150_245 ();
 sg13g2_decap_8 FILLER_0_150_252 ();
 sg13g2_decap_8 FILLER_0_150_259 ();
 sg13g2_decap_8 FILLER_0_150_266 ();
 sg13g2_decap_8 FILLER_0_150_273 ();
 sg13g2_decap_8 FILLER_0_150_280 ();
 sg13g2_decap_8 FILLER_0_150_287 ();
 sg13g2_decap_8 FILLER_0_150_294 ();
 sg13g2_decap_8 FILLER_0_150_301 ();
 sg13g2_decap_8 FILLER_0_150_308 ();
 sg13g2_decap_8 FILLER_0_150_315 ();
 sg13g2_decap_8 FILLER_0_150_322 ();
 sg13g2_decap_8 FILLER_0_150_329 ();
 sg13g2_decap_8 FILLER_0_150_336 ();
 sg13g2_decap_8 FILLER_0_150_343 ();
 sg13g2_decap_8 FILLER_0_150_350 ();
 sg13g2_decap_8 FILLER_0_150_357 ();
 sg13g2_decap_8 FILLER_0_150_364 ();
 sg13g2_decap_8 FILLER_0_150_371 ();
 sg13g2_decap_8 FILLER_0_150_378 ();
 sg13g2_decap_8 FILLER_0_150_385 ();
 sg13g2_decap_8 FILLER_0_150_392 ();
 sg13g2_decap_8 FILLER_0_150_399 ();
 sg13g2_decap_8 FILLER_0_150_406 ();
 sg13g2_decap_8 FILLER_0_150_413 ();
 sg13g2_decap_8 FILLER_0_150_420 ();
 sg13g2_decap_8 FILLER_0_150_427 ();
 sg13g2_decap_8 FILLER_0_150_434 ();
 sg13g2_decap_8 FILLER_0_150_441 ();
 sg13g2_decap_8 FILLER_0_150_448 ();
 sg13g2_decap_8 FILLER_0_150_455 ();
 sg13g2_decap_8 FILLER_0_150_462 ();
 sg13g2_decap_8 FILLER_0_150_469 ();
 sg13g2_decap_8 FILLER_0_150_476 ();
 sg13g2_decap_8 FILLER_0_150_483 ();
 sg13g2_decap_8 FILLER_0_150_490 ();
 sg13g2_decap_8 FILLER_0_150_497 ();
 sg13g2_decap_8 FILLER_0_150_504 ();
 sg13g2_decap_8 FILLER_0_150_511 ();
 sg13g2_decap_8 FILLER_0_150_518 ();
 sg13g2_decap_8 FILLER_0_150_525 ();
 sg13g2_decap_8 FILLER_0_150_532 ();
 sg13g2_decap_8 FILLER_0_150_539 ();
 sg13g2_decap_8 FILLER_0_150_546 ();
 sg13g2_decap_8 FILLER_0_150_553 ();
 sg13g2_decap_8 FILLER_0_150_560 ();
 sg13g2_decap_8 FILLER_0_150_567 ();
 sg13g2_decap_8 FILLER_0_150_574 ();
 sg13g2_decap_8 FILLER_0_150_581 ();
 sg13g2_decap_8 FILLER_0_150_588 ();
 sg13g2_decap_8 FILLER_0_150_595 ();
 sg13g2_decap_8 FILLER_0_150_602 ();
 sg13g2_decap_8 FILLER_0_150_609 ();
 sg13g2_decap_8 FILLER_0_150_616 ();
 sg13g2_decap_8 FILLER_0_150_623 ();
 sg13g2_fill_2 FILLER_0_150_630 ();
 sg13g2_fill_1 FILLER_0_150_632 ();
 sg13g2_fill_1 FILLER_0_150_663 ();
 sg13g2_decap_4 FILLER_0_150_674 ();
 sg13g2_fill_1 FILLER_0_150_678 ();
 sg13g2_decap_8 FILLER_0_150_684 ();
 sg13g2_fill_2 FILLER_0_150_691 ();
 sg13g2_fill_1 FILLER_0_150_693 ();
 sg13g2_decap_4 FILLER_0_150_735 ();
 sg13g2_fill_1 FILLER_0_150_749 ();
 sg13g2_fill_1 FILLER_0_150_753 ();
 sg13g2_decap_8 FILLER_0_150_762 ();
 sg13g2_fill_1 FILLER_0_150_769 ();
 sg13g2_decap_8 FILLER_0_150_774 ();
 sg13g2_decap_8 FILLER_0_150_781 ();
 sg13g2_decap_4 FILLER_0_150_788 ();
 sg13g2_fill_1 FILLER_0_150_792 ();
 sg13g2_fill_2 FILLER_0_150_801 ();
 sg13g2_decap_8 FILLER_0_150_811 ();
 sg13g2_decap_4 FILLER_0_150_818 ();
 sg13g2_fill_1 FILLER_0_150_822 ();
 sg13g2_decap_8 FILLER_0_150_827 ();
 sg13g2_decap_8 FILLER_0_150_834 ();
 sg13g2_decap_8 FILLER_0_150_841 ();
 sg13g2_fill_1 FILLER_0_150_848 ();
 sg13g2_decap_4 FILLER_0_150_853 ();
 sg13g2_fill_2 FILLER_0_150_857 ();
 sg13g2_fill_1 FILLER_0_150_864 ();
 sg13g2_decap_8 FILLER_0_150_891 ();
 sg13g2_decap_8 FILLER_0_150_898 ();
 sg13g2_decap_8 FILLER_0_150_905 ();
 sg13g2_decap_8 FILLER_0_150_912 ();
 sg13g2_decap_4 FILLER_0_150_919 ();
 sg13g2_decap_8 FILLER_0_150_949 ();
 sg13g2_decap_4 FILLER_0_150_956 ();
 sg13g2_fill_2 FILLER_0_150_960 ();
 sg13g2_decap_8 FILLER_0_150_966 ();
 sg13g2_decap_8 FILLER_0_150_973 ();
 sg13g2_decap_4 FILLER_0_150_980 ();
 sg13g2_fill_1 FILLER_0_150_984 ();
 sg13g2_decap_4 FILLER_0_150_1033 ();
 sg13g2_fill_1 FILLER_0_150_1037 ();
 sg13g2_fill_2 FILLER_0_150_1043 ();
 sg13g2_decap_8 FILLER_0_150_1053 ();
 sg13g2_decap_8 FILLER_0_150_1065 ();
 sg13g2_decap_8 FILLER_0_150_1072 ();
 sg13g2_decap_4 FILLER_0_150_1079 ();
 sg13g2_fill_2 FILLER_0_150_1083 ();
 sg13g2_fill_2 FILLER_0_150_1115 ();
 sg13g2_decap_8 FILLER_0_150_1121 ();
 sg13g2_decap_8 FILLER_0_150_1128 ();
 sg13g2_decap_8 FILLER_0_150_1135 ();
 sg13g2_decap_8 FILLER_0_150_1142 ();
 sg13g2_decap_8 FILLER_0_150_1149 ();
 sg13g2_decap_8 FILLER_0_150_1156 ();
 sg13g2_decap_8 FILLER_0_150_1163 ();
 sg13g2_decap_8 FILLER_0_150_1170 ();
 sg13g2_decap_8 FILLER_0_150_1177 ();
 sg13g2_decap_8 FILLER_0_150_1184 ();
 sg13g2_decap_8 FILLER_0_150_1191 ();
 sg13g2_decap_8 FILLER_0_150_1198 ();
 sg13g2_decap_8 FILLER_0_150_1205 ();
 sg13g2_decap_8 FILLER_0_150_1212 ();
 sg13g2_decap_8 FILLER_0_150_1219 ();
 sg13g2_fill_2 FILLER_0_150_1226 ();
 sg13g2_fill_1 FILLER_0_151_0 ();
 sg13g2_fill_1 FILLER_0_151_27 ();
 sg13g2_fill_1 FILLER_0_151_33 ();
 sg13g2_fill_2 FILLER_0_151_39 ();
 sg13g2_fill_1 FILLER_0_151_51 ();
 sg13g2_decap_8 FILLER_0_151_140 ();
 sg13g2_decap_8 FILLER_0_151_147 ();
 sg13g2_decap_8 FILLER_0_151_154 ();
 sg13g2_decap_8 FILLER_0_151_161 ();
 sg13g2_decap_8 FILLER_0_151_168 ();
 sg13g2_decap_8 FILLER_0_151_175 ();
 sg13g2_decap_8 FILLER_0_151_182 ();
 sg13g2_decap_8 FILLER_0_151_189 ();
 sg13g2_decap_8 FILLER_0_151_196 ();
 sg13g2_decap_8 FILLER_0_151_203 ();
 sg13g2_decap_8 FILLER_0_151_210 ();
 sg13g2_decap_8 FILLER_0_151_217 ();
 sg13g2_decap_8 FILLER_0_151_224 ();
 sg13g2_decap_8 FILLER_0_151_231 ();
 sg13g2_decap_8 FILLER_0_151_238 ();
 sg13g2_decap_8 FILLER_0_151_245 ();
 sg13g2_decap_8 FILLER_0_151_252 ();
 sg13g2_decap_8 FILLER_0_151_259 ();
 sg13g2_decap_8 FILLER_0_151_266 ();
 sg13g2_decap_8 FILLER_0_151_273 ();
 sg13g2_decap_8 FILLER_0_151_280 ();
 sg13g2_decap_8 FILLER_0_151_287 ();
 sg13g2_decap_8 FILLER_0_151_294 ();
 sg13g2_decap_8 FILLER_0_151_301 ();
 sg13g2_decap_8 FILLER_0_151_308 ();
 sg13g2_decap_8 FILLER_0_151_315 ();
 sg13g2_decap_8 FILLER_0_151_322 ();
 sg13g2_decap_8 FILLER_0_151_329 ();
 sg13g2_decap_8 FILLER_0_151_336 ();
 sg13g2_decap_8 FILLER_0_151_343 ();
 sg13g2_decap_8 FILLER_0_151_350 ();
 sg13g2_decap_8 FILLER_0_151_357 ();
 sg13g2_decap_8 FILLER_0_151_364 ();
 sg13g2_decap_8 FILLER_0_151_371 ();
 sg13g2_decap_8 FILLER_0_151_378 ();
 sg13g2_decap_8 FILLER_0_151_385 ();
 sg13g2_decap_8 FILLER_0_151_392 ();
 sg13g2_decap_8 FILLER_0_151_399 ();
 sg13g2_decap_8 FILLER_0_151_406 ();
 sg13g2_decap_8 FILLER_0_151_413 ();
 sg13g2_decap_8 FILLER_0_151_420 ();
 sg13g2_decap_8 FILLER_0_151_427 ();
 sg13g2_decap_8 FILLER_0_151_434 ();
 sg13g2_decap_8 FILLER_0_151_441 ();
 sg13g2_decap_8 FILLER_0_151_448 ();
 sg13g2_decap_8 FILLER_0_151_455 ();
 sg13g2_decap_8 FILLER_0_151_462 ();
 sg13g2_decap_8 FILLER_0_151_469 ();
 sg13g2_decap_8 FILLER_0_151_476 ();
 sg13g2_decap_8 FILLER_0_151_483 ();
 sg13g2_decap_8 FILLER_0_151_490 ();
 sg13g2_decap_8 FILLER_0_151_497 ();
 sg13g2_decap_8 FILLER_0_151_504 ();
 sg13g2_decap_8 FILLER_0_151_511 ();
 sg13g2_decap_8 FILLER_0_151_518 ();
 sg13g2_decap_8 FILLER_0_151_525 ();
 sg13g2_decap_8 FILLER_0_151_532 ();
 sg13g2_decap_8 FILLER_0_151_539 ();
 sg13g2_decap_8 FILLER_0_151_546 ();
 sg13g2_decap_8 FILLER_0_151_553 ();
 sg13g2_decap_8 FILLER_0_151_560 ();
 sg13g2_decap_8 FILLER_0_151_567 ();
 sg13g2_decap_8 FILLER_0_151_574 ();
 sg13g2_decap_8 FILLER_0_151_581 ();
 sg13g2_decap_8 FILLER_0_151_588 ();
 sg13g2_decap_8 FILLER_0_151_595 ();
 sg13g2_decap_8 FILLER_0_151_602 ();
 sg13g2_decap_8 FILLER_0_151_609 ();
 sg13g2_decap_8 FILLER_0_151_616 ();
 sg13g2_decap_8 FILLER_0_151_623 ();
 sg13g2_decap_8 FILLER_0_151_630 ();
 sg13g2_decap_4 FILLER_0_151_637 ();
 sg13g2_decap_4 FILLER_0_151_697 ();
 sg13g2_decap_8 FILLER_0_151_705 ();
 sg13g2_decap_8 FILLER_0_151_712 ();
 sg13g2_fill_2 FILLER_0_151_719 ();
 sg13g2_fill_1 FILLER_0_151_721 ();
 sg13g2_decap_4 FILLER_0_151_753 ();
 sg13g2_decap_8 FILLER_0_151_772 ();
 sg13g2_fill_1 FILLER_0_151_794 ();
 sg13g2_decap_8 FILLER_0_151_831 ();
 sg13g2_decap_8 FILLER_0_151_838 ();
 sg13g2_decap_4 FILLER_0_151_845 ();
 sg13g2_decap_8 FILLER_0_151_853 ();
 sg13g2_decap_8 FILLER_0_151_860 ();
 sg13g2_decap_4 FILLER_0_151_867 ();
 sg13g2_decap_4 FILLER_0_151_875 ();
 sg13g2_fill_1 FILLER_0_151_879 ();
 sg13g2_fill_1 FILLER_0_151_915 ();
 sg13g2_decap_8 FILLER_0_151_926 ();
 sg13g2_decap_8 FILLER_0_151_933 ();
 sg13g2_fill_2 FILLER_0_151_940 ();
 sg13g2_fill_1 FILLER_0_151_942 ();
 sg13g2_fill_1 FILLER_0_151_958 ();
 sg13g2_decap_4 FILLER_0_151_971 ();
 sg13g2_fill_2 FILLER_0_151_1011 ();
 sg13g2_fill_1 FILLER_0_151_1013 ();
 sg13g2_fill_1 FILLER_0_151_1066 ();
 sg13g2_fill_2 FILLER_0_151_1082 ();
 sg13g2_fill_1 FILLER_0_151_1084 ();
 sg13g2_fill_2 FILLER_0_151_1090 ();
 sg13g2_decap_8 FILLER_0_151_1118 ();
 sg13g2_decap_8 FILLER_0_151_1125 ();
 sg13g2_decap_8 FILLER_0_151_1132 ();
 sg13g2_decap_8 FILLER_0_151_1139 ();
 sg13g2_decap_8 FILLER_0_151_1146 ();
 sg13g2_decap_8 FILLER_0_151_1153 ();
 sg13g2_decap_8 FILLER_0_151_1160 ();
 sg13g2_decap_8 FILLER_0_151_1167 ();
 sg13g2_decap_8 FILLER_0_151_1174 ();
 sg13g2_decap_8 FILLER_0_151_1181 ();
 sg13g2_decap_8 FILLER_0_151_1188 ();
 sg13g2_decap_8 FILLER_0_151_1195 ();
 sg13g2_decap_8 FILLER_0_151_1202 ();
 sg13g2_decap_8 FILLER_0_151_1209 ();
 sg13g2_decap_8 FILLER_0_151_1216 ();
 sg13g2_decap_4 FILLER_0_151_1223 ();
 sg13g2_fill_1 FILLER_0_151_1227 ();
 sg13g2_decap_4 FILLER_0_152_0 ();
 sg13g2_fill_1 FILLER_0_152_4 ();
 sg13g2_fill_1 FILLER_0_152_9 ();
 sg13g2_fill_1 FILLER_0_152_62 ();
 sg13g2_fill_1 FILLER_0_152_94 ();
 sg13g2_decap_8 FILLER_0_152_133 ();
 sg13g2_decap_8 FILLER_0_152_140 ();
 sg13g2_decap_8 FILLER_0_152_147 ();
 sg13g2_decap_8 FILLER_0_152_154 ();
 sg13g2_decap_8 FILLER_0_152_161 ();
 sg13g2_decap_8 FILLER_0_152_168 ();
 sg13g2_decap_8 FILLER_0_152_175 ();
 sg13g2_decap_8 FILLER_0_152_182 ();
 sg13g2_decap_8 FILLER_0_152_189 ();
 sg13g2_decap_8 FILLER_0_152_196 ();
 sg13g2_decap_8 FILLER_0_152_203 ();
 sg13g2_decap_8 FILLER_0_152_210 ();
 sg13g2_decap_8 FILLER_0_152_217 ();
 sg13g2_decap_8 FILLER_0_152_224 ();
 sg13g2_decap_8 FILLER_0_152_231 ();
 sg13g2_decap_8 FILLER_0_152_238 ();
 sg13g2_decap_8 FILLER_0_152_245 ();
 sg13g2_decap_8 FILLER_0_152_252 ();
 sg13g2_decap_8 FILLER_0_152_259 ();
 sg13g2_decap_8 FILLER_0_152_266 ();
 sg13g2_decap_8 FILLER_0_152_273 ();
 sg13g2_decap_8 FILLER_0_152_280 ();
 sg13g2_decap_8 FILLER_0_152_287 ();
 sg13g2_decap_8 FILLER_0_152_294 ();
 sg13g2_decap_8 FILLER_0_152_301 ();
 sg13g2_decap_8 FILLER_0_152_308 ();
 sg13g2_decap_8 FILLER_0_152_315 ();
 sg13g2_decap_8 FILLER_0_152_322 ();
 sg13g2_decap_8 FILLER_0_152_329 ();
 sg13g2_decap_8 FILLER_0_152_336 ();
 sg13g2_decap_8 FILLER_0_152_343 ();
 sg13g2_decap_8 FILLER_0_152_350 ();
 sg13g2_decap_8 FILLER_0_152_357 ();
 sg13g2_decap_8 FILLER_0_152_364 ();
 sg13g2_decap_8 FILLER_0_152_371 ();
 sg13g2_decap_8 FILLER_0_152_378 ();
 sg13g2_decap_8 FILLER_0_152_385 ();
 sg13g2_decap_8 FILLER_0_152_392 ();
 sg13g2_decap_8 FILLER_0_152_399 ();
 sg13g2_decap_8 FILLER_0_152_406 ();
 sg13g2_decap_8 FILLER_0_152_413 ();
 sg13g2_decap_8 FILLER_0_152_420 ();
 sg13g2_decap_8 FILLER_0_152_427 ();
 sg13g2_decap_8 FILLER_0_152_434 ();
 sg13g2_decap_8 FILLER_0_152_441 ();
 sg13g2_decap_8 FILLER_0_152_448 ();
 sg13g2_decap_8 FILLER_0_152_455 ();
 sg13g2_decap_8 FILLER_0_152_462 ();
 sg13g2_decap_8 FILLER_0_152_469 ();
 sg13g2_decap_8 FILLER_0_152_476 ();
 sg13g2_decap_8 FILLER_0_152_483 ();
 sg13g2_decap_8 FILLER_0_152_490 ();
 sg13g2_decap_8 FILLER_0_152_497 ();
 sg13g2_decap_8 FILLER_0_152_504 ();
 sg13g2_decap_8 FILLER_0_152_511 ();
 sg13g2_decap_8 FILLER_0_152_518 ();
 sg13g2_decap_8 FILLER_0_152_525 ();
 sg13g2_decap_8 FILLER_0_152_532 ();
 sg13g2_decap_8 FILLER_0_152_539 ();
 sg13g2_decap_8 FILLER_0_152_546 ();
 sg13g2_decap_8 FILLER_0_152_553 ();
 sg13g2_decap_8 FILLER_0_152_560 ();
 sg13g2_decap_8 FILLER_0_152_567 ();
 sg13g2_decap_8 FILLER_0_152_574 ();
 sg13g2_decap_8 FILLER_0_152_581 ();
 sg13g2_decap_8 FILLER_0_152_588 ();
 sg13g2_decap_8 FILLER_0_152_595 ();
 sg13g2_decap_8 FILLER_0_152_602 ();
 sg13g2_decap_8 FILLER_0_152_609 ();
 sg13g2_decap_8 FILLER_0_152_616 ();
 sg13g2_decap_8 FILLER_0_152_623 ();
 sg13g2_decap_8 FILLER_0_152_630 ();
 sg13g2_decap_8 FILLER_0_152_637 ();
 sg13g2_fill_1 FILLER_0_152_644 ();
 sg13g2_decap_4 FILLER_0_152_650 ();
 sg13g2_fill_1 FILLER_0_152_654 ();
 sg13g2_fill_2 FILLER_0_152_660 ();
 sg13g2_fill_1 FILLER_0_152_672 ();
 sg13g2_fill_1 FILLER_0_152_686 ();
 sg13g2_decap_4 FILLER_0_152_718 ();
 sg13g2_fill_2 FILLER_0_152_732 ();
 sg13g2_fill_1 FILLER_0_152_734 ();
 sg13g2_decap_4 FILLER_0_152_777 ();
 sg13g2_fill_1 FILLER_0_152_807 ();
 sg13g2_fill_2 FILLER_0_152_834 ();
 sg13g2_fill_2 FILLER_0_152_840 ();
 sg13g2_decap_4 FILLER_0_152_868 ();
 sg13g2_fill_1 FILLER_0_152_872 ();
 sg13g2_decap_8 FILLER_0_152_982 ();
 sg13g2_fill_2 FILLER_0_152_1003 ();
 sg13g2_fill_1 FILLER_0_152_1005 ();
 sg13g2_fill_2 FILLER_0_152_1014 ();
 sg13g2_decap_8 FILLER_0_152_1113 ();
 sg13g2_decap_8 FILLER_0_152_1120 ();
 sg13g2_decap_8 FILLER_0_152_1127 ();
 sg13g2_decap_8 FILLER_0_152_1134 ();
 sg13g2_decap_8 FILLER_0_152_1141 ();
 sg13g2_decap_8 FILLER_0_152_1148 ();
 sg13g2_decap_8 FILLER_0_152_1155 ();
 sg13g2_decap_8 FILLER_0_152_1162 ();
 sg13g2_decap_8 FILLER_0_152_1169 ();
 sg13g2_decap_8 FILLER_0_152_1176 ();
 sg13g2_decap_8 FILLER_0_152_1183 ();
 sg13g2_decap_8 FILLER_0_152_1190 ();
 sg13g2_decap_8 FILLER_0_152_1197 ();
 sg13g2_decap_8 FILLER_0_152_1204 ();
 sg13g2_decap_8 FILLER_0_152_1211 ();
 sg13g2_decap_8 FILLER_0_152_1218 ();
 sg13g2_fill_2 FILLER_0_152_1225 ();
 sg13g2_fill_1 FILLER_0_152_1227 ();
 sg13g2_decap_8 FILLER_0_153_9 ();
 sg13g2_fill_2 FILLER_0_153_16 ();
 sg13g2_decap_8 FILLER_0_153_22 ();
 sg13g2_decap_4 FILLER_0_153_29 ();
 sg13g2_fill_2 FILLER_0_153_33 ();
 sg13g2_fill_2 FILLER_0_153_74 ();
 sg13g2_decap_8 FILLER_0_153_112 ();
 sg13g2_decap_8 FILLER_0_153_122 ();
 sg13g2_decap_8 FILLER_0_153_129 ();
 sg13g2_decap_8 FILLER_0_153_136 ();
 sg13g2_decap_8 FILLER_0_153_143 ();
 sg13g2_decap_8 FILLER_0_153_150 ();
 sg13g2_decap_8 FILLER_0_153_157 ();
 sg13g2_decap_8 FILLER_0_153_164 ();
 sg13g2_decap_8 FILLER_0_153_171 ();
 sg13g2_decap_8 FILLER_0_153_178 ();
 sg13g2_decap_8 FILLER_0_153_185 ();
 sg13g2_decap_8 FILLER_0_153_192 ();
 sg13g2_decap_8 FILLER_0_153_199 ();
 sg13g2_decap_8 FILLER_0_153_206 ();
 sg13g2_decap_8 FILLER_0_153_213 ();
 sg13g2_decap_8 FILLER_0_153_220 ();
 sg13g2_decap_8 FILLER_0_153_227 ();
 sg13g2_decap_8 FILLER_0_153_234 ();
 sg13g2_decap_8 FILLER_0_153_241 ();
 sg13g2_decap_8 FILLER_0_153_248 ();
 sg13g2_decap_8 FILLER_0_153_255 ();
 sg13g2_decap_8 FILLER_0_153_262 ();
 sg13g2_decap_8 FILLER_0_153_269 ();
 sg13g2_decap_8 FILLER_0_153_276 ();
 sg13g2_decap_8 FILLER_0_153_283 ();
 sg13g2_decap_8 FILLER_0_153_290 ();
 sg13g2_decap_8 FILLER_0_153_297 ();
 sg13g2_decap_8 FILLER_0_153_304 ();
 sg13g2_decap_8 FILLER_0_153_311 ();
 sg13g2_decap_8 FILLER_0_153_318 ();
 sg13g2_decap_8 FILLER_0_153_325 ();
 sg13g2_decap_8 FILLER_0_153_332 ();
 sg13g2_decap_8 FILLER_0_153_339 ();
 sg13g2_decap_8 FILLER_0_153_346 ();
 sg13g2_decap_8 FILLER_0_153_353 ();
 sg13g2_decap_8 FILLER_0_153_360 ();
 sg13g2_decap_8 FILLER_0_153_367 ();
 sg13g2_decap_8 FILLER_0_153_374 ();
 sg13g2_decap_8 FILLER_0_153_381 ();
 sg13g2_decap_8 FILLER_0_153_388 ();
 sg13g2_decap_8 FILLER_0_153_395 ();
 sg13g2_decap_8 FILLER_0_153_402 ();
 sg13g2_decap_8 FILLER_0_153_409 ();
 sg13g2_decap_8 FILLER_0_153_416 ();
 sg13g2_decap_8 FILLER_0_153_423 ();
 sg13g2_decap_8 FILLER_0_153_430 ();
 sg13g2_decap_8 FILLER_0_153_437 ();
 sg13g2_decap_8 FILLER_0_153_444 ();
 sg13g2_decap_8 FILLER_0_153_451 ();
 sg13g2_decap_8 FILLER_0_153_458 ();
 sg13g2_decap_8 FILLER_0_153_465 ();
 sg13g2_decap_8 FILLER_0_153_472 ();
 sg13g2_decap_8 FILLER_0_153_479 ();
 sg13g2_decap_8 FILLER_0_153_486 ();
 sg13g2_decap_8 FILLER_0_153_493 ();
 sg13g2_decap_8 FILLER_0_153_500 ();
 sg13g2_decap_8 FILLER_0_153_507 ();
 sg13g2_decap_8 FILLER_0_153_514 ();
 sg13g2_decap_8 FILLER_0_153_521 ();
 sg13g2_decap_8 FILLER_0_153_528 ();
 sg13g2_decap_8 FILLER_0_153_535 ();
 sg13g2_decap_8 FILLER_0_153_542 ();
 sg13g2_decap_8 FILLER_0_153_549 ();
 sg13g2_decap_8 FILLER_0_153_556 ();
 sg13g2_decap_8 FILLER_0_153_563 ();
 sg13g2_decap_8 FILLER_0_153_570 ();
 sg13g2_decap_8 FILLER_0_153_577 ();
 sg13g2_decap_8 FILLER_0_153_584 ();
 sg13g2_decap_8 FILLER_0_153_591 ();
 sg13g2_decap_8 FILLER_0_153_598 ();
 sg13g2_decap_8 FILLER_0_153_605 ();
 sg13g2_decap_8 FILLER_0_153_612 ();
 sg13g2_decap_8 FILLER_0_153_619 ();
 sg13g2_decap_8 FILLER_0_153_626 ();
 sg13g2_decap_8 FILLER_0_153_633 ();
 sg13g2_decap_8 FILLER_0_153_640 ();
 sg13g2_fill_2 FILLER_0_153_647 ();
 sg13g2_fill_1 FILLER_0_153_649 ();
 sg13g2_decap_4 FILLER_0_153_676 ();
 sg13g2_fill_2 FILLER_0_153_688 ();
 sg13g2_fill_2 FILLER_0_153_700 ();
 sg13g2_fill_2 FILLER_0_153_728 ();
 sg13g2_fill_2 FILLER_0_153_756 ();
 sg13g2_fill_1 FILLER_0_153_792 ();
 sg13g2_fill_1 FILLER_0_153_798 ();
 sg13g2_fill_1 FILLER_0_153_809 ();
 sg13g2_fill_1 FILLER_0_153_815 ();
 sg13g2_fill_1 FILLER_0_153_826 ();
 sg13g2_fill_1 FILLER_0_153_858 ();
 sg13g2_fill_2 FILLER_0_153_885 ();
 sg13g2_fill_1 FILLER_0_153_887 ();
 sg13g2_decap_8 FILLER_0_153_892 ();
 sg13g2_fill_1 FILLER_0_153_899 ();
 sg13g2_fill_2 FILLER_0_153_915 ();
 sg13g2_fill_2 FILLER_0_153_940 ();
 sg13g2_fill_1 FILLER_0_153_968 ();
 sg13g2_fill_2 FILLER_0_153_995 ();
 sg13g2_fill_1 FILLER_0_153_1002 ();
 sg13g2_fill_2 FILLER_0_153_1007 ();
 sg13g2_fill_2 FILLER_0_153_1019 ();
 sg13g2_fill_2 FILLER_0_153_1025 ();
 sg13g2_decap_4 FILLER_0_153_1065 ();
 sg13g2_decap_8 FILLER_0_153_1099 ();
 sg13g2_decap_8 FILLER_0_153_1106 ();
 sg13g2_decap_8 FILLER_0_153_1113 ();
 sg13g2_decap_8 FILLER_0_153_1120 ();
 sg13g2_decap_8 FILLER_0_153_1127 ();
 sg13g2_decap_8 FILLER_0_153_1134 ();
 sg13g2_decap_8 FILLER_0_153_1141 ();
 sg13g2_decap_8 FILLER_0_153_1148 ();
 sg13g2_decap_8 FILLER_0_153_1155 ();
 sg13g2_decap_8 FILLER_0_153_1162 ();
 sg13g2_decap_8 FILLER_0_153_1169 ();
 sg13g2_decap_8 FILLER_0_153_1176 ();
 sg13g2_decap_8 FILLER_0_153_1183 ();
 sg13g2_decap_8 FILLER_0_153_1190 ();
 sg13g2_decap_8 FILLER_0_153_1197 ();
 sg13g2_decap_8 FILLER_0_153_1204 ();
 sg13g2_decap_8 FILLER_0_153_1211 ();
 sg13g2_decap_8 FILLER_0_153_1218 ();
 sg13g2_fill_2 FILLER_0_153_1225 ();
 sg13g2_fill_1 FILLER_0_153_1227 ();
 sg13g2_decap_8 FILLER_0_154_15 ();
 sg13g2_decap_8 FILLER_0_154_22 ();
 sg13g2_decap_8 FILLER_0_154_29 ();
 sg13g2_decap_8 FILLER_0_154_36 ();
 sg13g2_decap_8 FILLER_0_154_43 ();
 sg13g2_fill_1 FILLER_0_154_50 ();
 sg13g2_fill_2 FILLER_0_154_60 ();
 sg13g2_decap_8 FILLER_0_154_66 ();
 sg13g2_decap_8 FILLER_0_154_73 ();
 sg13g2_decap_8 FILLER_0_154_80 ();
 sg13g2_decap_4 FILLER_0_154_87 ();
 sg13g2_fill_2 FILLER_0_154_91 ();
 sg13g2_decap_4 FILLER_0_154_97 ();
 sg13g2_fill_2 FILLER_0_154_101 ();
 sg13g2_decap_8 FILLER_0_154_107 ();
 sg13g2_decap_8 FILLER_0_154_114 ();
 sg13g2_decap_8 FILLER_0_154_121 ();
 sg13g2_decap_8 FILLER_0_154_128 ();
 sg13g2_decap_8 FILLER_0_154_135 ();
 sg13g2_decap_8 FILLER_0_154_142 ();
 sg13g2_decap_8 FILLER_0_154_149 ();
 sg13g2_decap_8 FILLER_0_154_156 ();
 sg13g2_decap_8 FILLER_0_154_163 ();
 sg13g2_decap_8 FILLER_0_154_170 ();
 sg13g2_decap_8 FILLER_0_154_177 ();
 sg13g2_decap_8 FILLER_0_154_184 ();
 sg13g2_decap_8 FILLER_0_154_191 ();
 sg13g2_decap_8 FILLER_0_154_198 ();
 sg13g2_decap_8 FILLER_0_154_205 ();
 sg13g2_decap_8 FILLER_0_154_212 ();
 sg13g2_decap_8 FILLER_0_154_219 ();
 sg13g2_decap_8 FILLER_0_154_226 ();
 sg13g2_decap_8 FILLER_0_154_233 ();
 sg13g2_decap_8 FILLER_0_154_240 ();
 sg13g2_decap_8 FILLER_0_154_247 ();
 sg13g2_decap_8 FILLER_0_154_254 ();
 sg13g2_decap_8 FILLER_0_154_261 ();
 sg13g2_decap_8 FILLER_0_154_268 ();
 sg13g2_decap_8 FILLER_0_154_275 ();
 sg13g2_decap_8 FILLER_0_154_282 ();
 sg13g2_decap_8 FILLER_0_154_289 ();
 sg13g2_decap_8 FILLER_0_154_296 ();
 sg13g2_decap_8 FILLER_0_154_303 ();
 sg13g2_decap_8 FILLER_0_154_310 ();
 sg13g2_decap_8 FILLER_0_154_317 ();
 sg13g2_decap_8 FILLER_0_154_324 ();
 sg13g2_decap_8 FILLER_0_154_331 ();
 sg13g2_decap_8 FILLER_0_154_338 ();
 sg13g2_decap_8 FILLER_0_154_345 ();
 sg13g2_decap_8 FILLER_0_154_352 ();
 sg13g2_decap_8 FILLER_0_154_359 ();
 sg13g2_decap_8 FILLER_0_154_366 ();
 sg13g2_decap_8 FILLER_0_154_373 ();
 sg13g2_decap_8 FILLER_0_154_380 ();
 sg13g2_decap_8 FILLER_0_154_387 ();
 sg13g2_decap_8 FILLER_0_154_394 ();
 sg13g2_decap_8 FILLER_0_154_401 ();
 sg13g2_decap_8 FILLER_0_154_408 ();
 sg13g2_decap_8 FILLER_0_154_415 ();
 sg13g2_decap_8 FILLER_0_154_422 ();
 sg13g2_decap_8 FILLER_0_154_429 ();
 sg13g2_decap_4 FILLER_0_154_436 ();
 sg13g2_decap_8 FILLER_0_154_443 ();
 sg13g2_decap_8 FILLER_0_154_450 ();
 sg13g2_decap_8 FILLER_0_154_457 ();
 sg13g2_decap_8 FILLER_0_154_464 ();
 sg13g2_decap_8 FILLER_0_154_471 ();
 sg13g2_decap_8 FILLER_0_154_478 ();
 sg13g2_decap_8 FILLER_0_154_485 ();
 sg13g2_decap_8 FILLER_0_154_492 ();
 sg13g2_decap_8 FILLER_0_154_499 ();
 sg13g2_decap_8 FILLER_0_154_506 ();
 sg13g2_decap_8 FILLER_0_154_513 ();
 sg13g2_decap_8 FILLER_0_154_520 ();
 sg13g2_decap_8 FILLER_0_154_527 ();
 sg13g2_decap_8 FILLER_0_154_534 ();
 sg13g2_decap_8 FILLER_0_154_541 ();
 sg13g2_decap_8 FILLER_0_154_548 ();
 sg13g2_decap_8 FILLER_0_154_555 ();
 sg13g2_decap_8 FILLER_0_154_562 ();
 sg13g2_decap_8 FILLER_0_154_569 ();
 sg13g2_decap_8 FILLER_0_154_576 ();
 sg13g2_decap_8 FILLER_0_154_583 ();
 sg13g2_decap_8 FILLER_0_154_590 ();
 sg13g2_decap_8 FILLER_0_154_597 ();
 sg13g2_decap_8 FILLER_0_154_604 ();
 sg13g2_decap_8 FILLER_0_154_611 ();
 sg13g2_decap_8 FILLER_0_154_618 ();
 sg13g2_decap_8 FILLER_0_154_625 ();
 sg13g2_decap_8 FILLER_0_154_632 ();
 sg13g2_decap_8 FILLER_0_154_639 ();
 sg13g2_decap_8 FILLER_0_154_646 ();
 sg13g2_fill_2 FILLER_0_154_653 ();
 sg13g2_fill_1 FILLER_0_154_655 ();
 sg13g2_decap_8 FILLER_0_154_660 ();
 sg13g2_decap_8 FILLER_0_154_667 ();
 sg13g2_decap_4 FILLER_0_154_674 ();
 sg13g2_fill_2 FILLER_0_154_682 ();
 sg13g2_decap_4 FILLER_0_154_689 ();
 sg13g2_fill_1 FILLER_0_154_693 ();
 sg13g2_decap_8 FILLER_0_154_698 ();
 sg13g2_fill_1 FILLER_0_154_705 ();
 sg13g2_decap_8 FILLER_0_154_720 ();
 sg13g2_fill_2 FILLER_0_154_727 ();
 sg13g2_decap_4 FILLER_0_154_734 ();
 sg13g2_fill_1 FILLER_0_154_738 ();
 sg13g2_fill_1 FILLER_0_154_753 ();
 sg13g2_decap_8 FILLER_0_154_759 ();
 sg13g2_fill_2 FILLER_0_154_766 ();
 sg13g2_fill_1 FILLER_0_154_768 ();
 sg13g2_decap_8 FILLER_0_154_773 ();
 sg13g2_decap_8 FILLER_0_154_780 ();
 sg13g2_decap_8 FILLER_0_154_787 ();
 sg13g2_decap_4 FILLER_0_154_794 ();
 sg13g2_fill_2 FILLER_0_154_798 ();
 sg13g2_decap_8 FILLER_0_154_804 ();
 sg13g2_decap_4 FILLER_0_154_811 ();
 sg13g2_fill_1 FILLER_0_154_819 ();
 sg13g2_decap_8 FILLER_0_154_825 ();
 sg13g2_decap_8 FILLER_0_154_832 ();
 sg13g2_decap_4 FILLER_0_154_839 ();
 sg13g2_fill_1 FILLER_0_154_843 ();
 sg13g2_fill_2 FILLER_0_154_859 ();
 sg13g2_decap_8 FILLER_0_154_875 ();
 sg13g2_decap_8 FILLER_0_154_882 ();
 sg13g2_fill_1 FILLER_0_154_889 ();
 sg13g2_decap_8 FILLER_0_154_898 ();
 sg13g2_decap_8 FILLER_0_154_905 ();
 sg13g2_fill_2 FILLER_0_154_938 ();
 sg13g2_fill_1 FILLER_0_154_955 ();
 sg13g2_decap_8 FILLER_0_154_960 ();
 sg13g2_fill_2 FILLER_0_154_967 ();
 sg13g2_fill_1 FILLER_0_154_969 ();
 sg13g2_fill_1 FILLER_0_154_980 ();
 sg13g2_decap_8 FILLER_0_154_985 ();
 sg13g2_decap_4 FILLER_0_154_992 ();
 sg13g2_decap_8 FILLER_0_154_1022 ();
 sg13g2_decap_8 FILLER_0_154_1029 ();
 sg13g2_decap_8 FILLER_0_154_1036 ();
 sg13g2_fill_2 FILLER_0_154_1043 ();
 sg13g2_decap_8 FILLER_0_154_1048 ();
 sg13g2_decap_4 FILLER_0_154_1055 ();
 sg13g2_fill_2 FILLER_0_154_1059 ();
 sg13g2_decap_8 FILLER_0_154_1065 ();
 sg13g2_decap_4 FILLER_0_154_1072 ();
 sg13g2_decap_8 FILLER_0_154_1080 ();
 sg13g2_decap_8 FILLER_0_154_1087 ();
 sg13g2_decap_8 FILLER_0_154_1094 ();
 sg13g2_decap_8 FILLER_0_154_1101 ();
 sg13g2_decap_8 FILLER_0_154_1108 ();
 sg13g2_decap_8 FILLER_0_154_1115 ();
 sg13g2_decap_8 FILLER_0_154_1122 ();
 sg13g2_decap_8 FILLER_0_154_1129 ();
 sg13g2_decap_8 FILLER_0_154_1136 ();
 sg13g2_decap_8 FILLER_0_154_1143 ();
 sg13g2_decap_8 FILLER_0_154_1150 ();
 sg13g2_decap_8 FILLER_0_154_1157 ();
 sg13g2_decap_8 FILLER_0_154_1164 ();
 sg13g2_decap_8 FILLER_0_154_1171 ();
 sg13g2_decap_8 FILLER_0_154_1178 ();
 sg13g2_decap_8 FILLER_0_154_1185 ();
 sg13g2_decap_8 FILLER_0_154_1192 ();
 sg13g2_decap_8 FILLER_0_154_1199 ();
 sg13g2_decap_8 FILLER_0_154_1206 ();
 sg13g2_decap_8 FILLER_0_154_1213 ();
 sg13g2_decap_8 FILLER_0_154_1220 ();
 sg13g2_fill_1 FILLER_0_154_1227 ();
endmodule
