`default_nettype none

module analog_blockage ();
endmodule
