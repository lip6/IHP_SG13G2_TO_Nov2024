** sch_path: /workspaces/usm-vlsi-tools/shared_xserver/TORepo_IHPNov2024_TDBuck/design_data/xschem/top/top.sch
.subckt AC3E_USM_TDBUCK 28 22 23 24 26 27 25 1 21 2 20 3 19 18 4 5 17 6 16 15 7 8 9 10 11 12 13 14
*.PININFO 1:B 2:B 3:B 4:B 5:B 6:B 7:B 8:B 9:B 10:B 11:B 12:B 13:B 14:B 15:B 16:B 17:B 18:B 19:B 20:B 21:B 22:B 23:B 24:B 25:B 26:B
*+ 27:B 28:B
X2 18 22 19 23 25 20 GD_vto1p1
X1 22 21 28 26 27 DCDCBuck_vto1p1
X3 17 21 19 23 25 20 GD_vto1p1
x4 19 25 13 17 18 14 DB
**** begin user architecture code


D1 28 1 25 diodevdd_2kv m=1
D2 28 2 25 diodevdd_2kv m=1
D3 28 3 25 diodevdd_2kv m=1
D4 28 4 25 diodevdd_2kv m=1
D5 28 5 25 diodevdd_2kv m=1
D6 28 6 25 diodevdd_2kv m=1
D7 28 7 25 diodevdd_2kv m=1
D8 28 8 25 diodevdd_2kv m=1
D9 28 9 25 diodevdd_2kv m=1
D10 28 10 25 diodevdd_2kv m=1
D11 28 11 25 diodevdd_2kv m=1
D12 28 12 25 diodevdd_2kv m=1
D13 28 13 25 diodevdd_2kv m=1
D14 28 14 25 diodevdd_2kv m=1
D15 28 15 25 diodevdd_2kv m=1
D16 28 16 25 diodevdd_2kv m=1
D17 28 17 25 diodevdd_2kv m=1
D18 28 18 25 diodevdd_2kv m=1
D19 28 19 25 diodevdd_2kv m=1
D20 28 20 25 diodevdd_2kv m=1
D21 28 21 25 diodevdd_2kv m=1
D22 28 22 25 diodevdd_2kv m=1
D23 28 23 25 diodevdd_2kv m=1
D24 28 24 25 diodevdd_2kv m=1
D25 28 25 25 diodevdd_2kv m=1
D26 28 26 25 diodevdd_2kv m=1
D27 28 27 25 diodevdd_2kv m=1
D28 28 28 25 diodevdd_2kv m=1

D29 28 1 25 diodevss_2kv m=1
D30 28 2 25 diodevss_2kv m=1
D31 28 3 25 diodevss_2kv m=1
D32 28 4 25 diodevss_2kv m=1
D33 28 5 25 diodevss_2kv m=1
D34 28 6 25 diodevss_2kv m=1
D35 28 7 25 diodevss_2kv m=1
D36 28 8 25 diodevss_2kv m=1
D37 28 9 25 diodevss_2kv m=1
D38 28 10 25 diodevss_2kv m=1
D39 28 11 25 diodevss_2kv m=1
D40 28 12 25 diodevss_2kv m=1
D41 28 13 25 diodevss_2kv m=1
D42 28 14 25 diodevss_2kv m=1
D43 28 15 25 diodevss_2kv m=1
D44 28 16 25 diodevss_2kv m=1
D45 28 17 25 diodevss_2kv m=1
D46 28 18 25 diodevss_2kv m=1
D47 28 19 25 diodevss_2kv m=1
D48 28 20 25 diodevss_2kv m=1
D49 28 21 25 diodevss_2kv m=1
D50 28 22 25 diodevss_2kv m=1
D51 28 23 25 diodevss_2kv m=1
D52 28 24 25 diodevss_2kv m=1
D53 28 25 25 diodevss_2kv m=1
D54 28 26 25 diodevss_2kv m=1
D55 28 27 25 diodevss_2kv m=1
D56 28 28 25 diodevss_2kv m=1


**** end user architecture code
.ends

* expanding   symbol:  /workspaces/usm-vlsi-tools/shared_xserver/TORepo_IHPNov2024_TDBuck/design_data/xschem/GD/GD_vto1p1.sym # of
*+ pins=6
** sym_path: /workspaces/usm-vlsi-tools/shared_xserver/TORepo_IHPNov2024_TDBuck/design_data/xschem/GD/GD_vto1p1.sym
** sch_path: /workspaces/usm-vlsi-tools/shared_xserver/TORepo_IHPNov2024_TDBuck/design_data/xschem/GD/GD_vto1p1.sch
.subckt GD_vto1p1 Vs Vg Vdd VH GND IGND
*.PININFO VH:B Vdd:B Vs:I Vg:O GND:B IGND:B
MD9 VgMD2 Vs Vdd Vdd sg13_lv_pmos l=0.13u w=1.12u ng=1 m=2
MD10 VgMD2 Vs GND GND sg13_lv_nmos l=0.13u w=1.12u ng=1 m=2
MD1 VgMD5 VgMD1 VH VH sg13_hv_pmos l=0.4u w=10u ng=1 m=1
MD3 VgMD1 VgMD5 VH VH sg13_hv_pmos l=0.4u w=10u ng=1 m=1
MD5 VgMD78 VgMD5 VH VH sg13_hv_pmos l=0.4u w=10u ng=1 m=30
MD7 Vg VgMD78 VH VH sg13_hv_pmos l=0.4u w=10u ng=1 m=250
MD2 VgMD5 VgMD2 IGND IGND sg13_hv_nmos l=0.45u w=10u ng=1 m=6
MD4 VgMD1 Vs IGND IGND sg13_hv_nmos l=0.45u w=10u ng=1 m=6
MD6 VgMD78 Vs IGND IGND sg13_hv_nmos l=0.45u w=10u ng=1 m=25
MD8 Vg VgMD78 IGND IGND sg13_hv_nmos l=0.45u w=10u ng=1 m=200
**** begin user architecture code


MD1D  VgMD5   VH   VH   VH   sg13_hv_pmos L=0.4u W=10u M=1
MD3D  VgMD1   VH   VH   VH   sg13_hv_pmos L=0.4u W=10u M=1
MD5D  VgMD78  VH   VH   VH   sg13_hv_pmos L=0.4u W=10u M=2
MDPD  VH      VH   VH   VH   sg13_hv_pmos L=0.4u W=10u M=14
MD2D  VgMD5   IGND  IGND  IGND  sg13_hv_nmos L=0.45u W=10u M=2
MD4D  VgMD1   IGND  IGND  IGND  sg13_hv_nmos L=0.45u W=10u M=2
MD6D  VgMD78  IGND  IGND  IGND  sg13_hv_nmos L=0.45u W=10u M=1
MDND  IGND     IGND  IGND  IGND  sg13_hv_nmos L=0.45u W=10u M=58


**** end user architecture code
.ends


* expanding   symbol:
*+  /workspaces/usm-vlsi-tools/shared_xserver/TORepo_IHPNov2024_TDBuck/design_data/xschem/DCDCBuck/DCDCBuck_vto1p1.sym # of pins=5
** sym_path: /workspaces/usm-vlsi-tools/shared_xserver/TORepo_IHPNov2024_TDBuck/design_data/xschem/DCDCBuck/DCDCBuck_vto1p1.sym
** sch_path: /workspaces/usm-vlsi-tools/shared_xserver/TORepo_IHPNov2024_TDBuck/design_data/xschem/DCDCBuck/DCDCBuck_vto1p1.sch
.subckt DCDCBuck_vto1p1 VgM1 VgM2 Vin GND Vo
*.PININFO Vin:B VgM1:I VgM2:I Vo:B GND:B
M2 Vo VgM2 GND GND sg13_hv_nmos l=0.45u w=10u ng=1 m=4080
M1 Vo VgM1 Vin Vin sg13_hv_pmos l=0.4u w=10u ng=1 m=12096
.ends


* expanding   symbol:  /workspaces/usm-vlsi-tools/shared_xserver/TORepo_IHPNov2024_TDBuck/design_data/xschem/Digital_Block/DB.sym
*+ # of pins=6
** sym_path: /workspaces/usm-vlsi-tools/shared_xserver/TORepo_IHPNov2024_TDBuck/design_data/xschem/Digital_Block/DB.sym
** sch_path: /workspaces/usm-vlsi-tools/shared_xserver/TORepo_IHPNov2024_TDBuck/design_data/xschem/Digital_Block/DB.sch
.subckt DB VCC VSS VINS VCN VCP VINR
*.PININFO VCC:B VSS:B VINS:B VINR:B VCP:B VCN:B
x2 VCC VSS VINS 16 VINR PD_vto1p1
x1 VCC VSS VCP 16 VCN NOL_vto1p1
.ends


* expanding   symbol:  /workspaces/usm-vlsi-tools/shared_xserver/TORepo_IHPNov2024_TDBuck/design_data/xschem/PD/PD_vto1p1.sym # of
*+ pins=5
** sym_path: /workspaces/usm-vlsi-tools/shared_xserver/TORepo_IHPNov2024_TDBuck/design_data/xschem/PD/PD_vto1p1.sym
** sch_path: /workspaces/usm-vlsi-tools/shared_xserver/TORepo_IHPNov2024_TDBuck/design_data/xschem/PD/PD_vto1p1.sch
.subckt PD_vto1p1 VCC VSS VINS V_PWM VINR
*.PININFO V_PWM:B VCC:B VSS:B VINS:B VINR:B
x3 net2 V_PWM VCC VSS V_N sg13g2_nor2_1
x1 V_N net1 VCC VSS V_PWM sg13g2_nor2_1
x4 VCC VSS VFE1 VINR net2 SPG_vto1p1
x2 VCC VSS VFE1 VINS net1 SPG_vto1p1
.ends


* expanding   symbol:  /workspaces/usm-vlsi-tools/shared_xserver/TORepo_IHPNov2024_TDBuck/design_data/xschem/NOL/NOL_vto1p1.sym #
*+ of pins=5
** sym_path: /workspaces/usm-vlsi-tools/shared_xserver/TORepo_IHPNov2024_TDBuck/design_data/xschem/NOL/NOL_vto1p1.sym
** sch_path: /workspaces/usm-vlsi-tools/shared_xserver/TORepo_IHPNov2024_TDBuck/design_data/xschem/NOL/NOL_vto1p1.sch
.subckt NOL_vto1p1 VCC VSS VCP CLK VCN
*.PININFO CLK:B VCP:B VCN:B VCC:B VSS:B
x5 CLK VCC VSS A1 sg13g2_inv_1
x3 A1 B1 VCC VSS C1 sg13g2_nor2_1
x1 B2 CLK VCC VSS C2 sg13g2_nor2_1
x2 B1 VCC VSS net1 sg13g2_inv_1
x6 B2 VCC VSS net2 sg13g2_inv_2
x7 net1 VCC VSS net3 sg13g2_inv_2
x8 net2 VCC VSS VCN sg13g2_inv_4
x9 net3 VCC VSS VCP sg13g2_inv_4
x10 VCC VSS C1 B2 large_delay_vto1p1
x4 VCC VSS C2 B1 large_delay_vto1p1
.ends


* expanding   symbol:  /workspaces/usm-vlsi-tools/shared_xserver/TORepo_IHPNov2024_TDBuck/design_data/xschem/SPG/SPG_vto1p1.sym #
*+ of pins=5
** sym_path: /workspaces/usm-vlsi-tools/shared_xserver/TORepo_IHPNov2024_TDBuck/design_data/xschem/SPG/SPG_vto1p1.sym
** sch_path: /workspaces/usm-vlsi-tools/shared_xserver/TORepo_IHPNov2024_TDBuck/design_data/xschem/SPG/SPG_vto1p1.sch
.subckt SPG_vto1p1 VCC VSS VFE VIN VRE
*.PININFO VIN:B VFE:B VRE:B VCC:B VSS:B
x1 dly7 VCC VSS dly8 sg13g2_inv_1
x2 predly VCC VSS net2 sg13g2_inv_1
x3 net3 VCC VSS predly sg13g2_inv_1
x4 dly8 VCC VSS net1 sg13g2_inv_1
x5 VIN VCC VSS net3 sg13g2_inv_2
x6 predly VCC VSS V_gatein sg13g2_inv_8
x7 net2 dly8 VCC VSS VFE sg13g2_and2_2
x8 net1 predly VCC VSS VRE sg13g2_and2_2
x9 VCC VSS V_gatein dly7 large_delay_vto1p1
.ends


* expanding   symbol:
*+  /workspaces/usm-vlsi-tools/shared_xserver/TORepo_IHPNov2024_TDBuck/design_data/xschem/large_delay/large_delay_vto1p1.sym # of pins=4
** sym_path: /workspaces/usm-vlsi-tools/shared_xserver/TORepo_IHPNov2024_TDBuck/design_data/xschem/large_delay/large_delay_vto1p1.sym
** sch_path: /workspaces/usm-vlsi-tools/shared_xserver/TORepo_IHPNov2024_TDBuck/design_data/xschem/large_delay/large_delay_vto1p1.sch
.subckt large_delay_vto1p1 VCC VSS VIN VOUT
*.PININFO VIN:B VOUT:B VCC:B VSS:B
x1[0] VIN VCC VSS n2 sg13g2_dlygate4sd3_1
x1[1] n2 VCC VSS n3 sg13g2_dlygate4sd3_1
x1[2] n3 VCC VSS n4 sg13g2_dlygate4sd3_1
x1[3] n4 VCC VSS n5 sg13g2_dlygate4sd3_1
x1[4] n5 VCC VSS VOUT sg13g2_dlygate4sd3_1
.ends

* Library name: sg13g2_stdcell
* Cell name: sg13g2_nor2_1
* View name: schematic
* Inherited view list: spectre cmos_sch cmos.sch schematic veriloga ahdl
* pspice dspf
.subckt sg13g2_nor2_1 A B VDD VSS Y
M0 Y A VSS VSS sg13_lv_nmos w=740.00n l=130.00n ng=1 ad=0 as=0 pd=0 ps=0 m=1
M3 Y B VSS VSS sg13_lv_nmos w=740.00n l=130.00n ng=1 ad=0 as=0 pd=0 ps=0 m=1
M1 net1 A VDD VDD sg13_lv_pmos w=1.12e-06 l=130.00n ng=1 ad=0 as=0 pd=0 ps=0 m=1
M2 Y B net1 VDD sg13_lv_pmos w=1.12e-06 l=130.00n ng=1 ad=0 as=0 pd=0 ps=0 m=1
.ends
* End of subcircuit definition.

* Library name: sg13g2_stdcell
* Cell name: sg13g2_inv_1
* View name: schematic
* Inherited view list: spectre cmos_sch cmos.sch schematic veriloga ahdl
* pspice dspf
.subckt sg13g2_inv_1 A VDD VSS Y
M1 Y A VSS VSS sg13_lv_nmos w=740.00n l=130.00n ng=1 ad=0 as=0 pd=0 ps=0 m=1
M0 Y A VDD VDD sg13_lv_pmos w=1.12u l=130.00n ng=1 ad=0 as=0 pd=0 ps=0 m=1
.ends
* End of subcircuit definition.

* Library name: sg13g2_stdcell
* Cell name: sg13g2_inv_2
* View name: schematic
* Inherited view list: spectre cmos_sch cmos.sch schematic veriloga ahdl
* pspice dspf
.subckt sg13g2_inv_2 A VDD VSS Y
M1 Y A VSS VSS sg13_lv_nmos w=740.00n l=130.00n ng=1 ad=0 as=0 pd=0 ps=0 m=2
M0 Y A VDD VDD sg13_lv_pmos w=1.12u l=130.00n ng=1 ad=0 as=0 pd=0 ps=0 m=2
.ends
* End of subcircuit definition.

* Library name: sg13g2_stdcell
* Cell name: sg13g2_inv_8
* View name: schematic
* Inherited view list: spectre cmos_sch cmos.sch schematic veriloga ahdl
* pspice dspf
.subckt sg13g2_inv_8 A VDD VSS Y
M1 Y A VSS VSS sg13_lv_nmos w=740.00n l=130.00n ng=1 ad=0 as=0 pd=0 ps=0 m=8
M0 Y A VDD VDD sg13_lv_pmos w=1.12u l=130.00n ng=1 ad=0 as=0 pd=0 ps=0 m=8
.ends
* End of subcircuit definition.

* Library name: sg13g2_stdcell
* Cell name: sg13g2_and2_2
* View name: schematic
* Inherited view list: spectre cmos_sch cmos.sch schematic veriloga ahdl
* pspice dspf
.subckt sg13g2_and2_2 A B VDD VSS X
M0 net4 A net2 VSS sg13_lv_nmos w=640.00n l=130.00n ng=1 ad=0 as=0 pd=0 ps=0 m=1
M2 X net4 VSS VSS sg13_lv_nmos w=740.00n l=130.00n ng=1 ad=0 as=0 pd=0 ps=0 m=2
M3 net2 B VSS VSS sg13_lv_nmos w=640.00n l=130.00n ng=1 ad=0 as=0 pd=0 ps=0 m=1
M1 net4 B VDD VDD sg13_lv_pmos w=840.00n l=130.00n ng=1 ad=0 as=0 pd=0 ps=0 m=1
M4 VDD net4 X VDD sg13_lv_pmos w=1.12u l=130.00n ng=1 ad=0 as=0 pd=0 ps=0 m=2
M5 net4 A VDD VDD sg13_lv_pmos w=840.00n l=130.00n ng=1 ad=0 as=0 pd=0 ps=0 m=1
.ends
* End of subcircuit definition.

* Library name: sg13g2_stdcell
* Cell name: sg13g2_dlygate4sd3_1
* View name: schematic
* Inherited view list: spectre cmos_sch cmos.sch schematic veriloga ahdl
* pspice dspf
.subckt sg13g2_dlygate4sd3_1 A VDD VSS X
MP3 X net3 VDD VDD sg13_lv_pmos w=1.12u l=130.00n ng=1 ad=0 as=0 pd=0 ps=0 m=1
MP2 net3 net2 VDD VDD sg13_lv_pmos w=1.000u l=500.0n ng=1 ad=0 as=0 pd=0 ps=0 m=1
MP1 net2 net1 VDD VDD sg13_lv_pmos w=1.000u l=500.0n ng=1 ad=0 as=0 pd=0 ps=0 m=1
MP0 net1 A VDD VDD sg13_lv_pmos w=420.00n l=130.00n ng=1 ad=0 as=0 pd=0 ps=0 m=1
MN3 X net3 VSS VSS sg13_lv_nmos w=740.00n l=130.00n ng=1 ad=0 as=0 pd=0 ps=0 m=1
MN2 net3 net2 VSS VSS sg13_lv_nmos w=420.00n l=500.0n ng=1 ad=0 as=0 pd=0 ps=0 m=1
MN1 net2 net1 VSS VSS sg13_lv_nmos w=420.00n l=500.0n ng=1 ad=0 as=0 pd=0 ps=0 m=1
MN0 net1 A VSS VSS sg13_lv_nmos w=420.00n l=130.00n ng=1 ad=0 as=0 pd=0 ps=0 m=1
.ends
* End of subcircuit definition.

* Library name: sg13g2_stdcell
* Cell name: sg13g2_inv_4
* View name: schematic
* Inherited view list: spectre cmos_sch cmos.sch schematic veriloga ahdl
* pspice dspf
.subckt sg13g2_inv_4 A VDD VSS Y
MP0 Y A VDD VDD sg13_lv_pmos w=1.12u l=130.00n ng=1 ad=0 as=0 pd=0 ps=0 m=4
MN0 Y A VSS VSS sg13_lv_nmos w=740.00n l=130.00n ng=1 ad=0 as=0 pd=0 ps=0 m=4
.ends
* End of subcircuit definition.

.end
