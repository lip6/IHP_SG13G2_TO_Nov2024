module controller(
    input clk, rst,
    input spi_done, 
    input [7:0] spi_input,
    output reg [7:0] control,
    output reg set_din,
    output reg set_data_in,
    output reg trig
);

wire result_ready;
assign result_ready = 1;
reg trig_ext;

localparam IDLE=0, SAVE_CMD=1, SAVE_DATA=2, TRIG_STATE=3, WAIT_RESULT=4, SEND_RESULT=5, SAVE_DIN=6, WAIT_DATA=7;
localparam SAVE_CMD_EXT=8, SAVE_DATA_EXT=9, SAVE_DIN_EXT=10, TRIG_EXT=11;

reg set_control, start_send;
reg [3:0] state, next_state;

always @(posedge clk) begin
    if(rst) state <= IDLE;
    else state <= next_state;
end

always @(*) begin
    next_state=state;
    set_control=0;//(state==SAVE_CMD||state==SAVE_CMD_EXT)?1:0;
    set_data_in=0;
    start_send=0;
    set_din=0;
    trig=0;
    trig_ext=0;
    case(state)
        IDLE: begin
            if(spi_done) begin
                next_state = SAVE_CMD;
            end
        end 
        SAVE_CMD: begin
            set_control=1;
            next_state = SAVE_CMD_EXT;
        end
        SAVE_CMD_EXT: begin
            set_control=1;
            next_state = WAIT_DATA;
        end
        WAIT_DATA: begin
            if(spi_done) begin
                if(control[7:6]==2'b00) next_state = SAVE_DATA;
                else if(control[7:6]==2'b01) next_state = SAVE_DIN;
                else if(control[7:6]==2'b10) next_state = TRIG_STATE;
                else if(control[7:6]==2'b11) next_state = SEND_RESULT;
            end
        end
        SAVE_DATA: begin
            set_data_in=1;
            next_state = SAVE_DATA_EXT;
        end
        SAVE_DATA_EXT: begin
            set_data_in=1;
            next_state = IDLE;
        end
        SAVE_DIN: begin
            set_din=1;
            next_state = SAVE_DIN_EXT;
        end
        SAVE_DIN_EXT: begin
            set_din=1;
            next_state = IDLE;
        end
        TRIG_STATE: begin
            trig = 1;
            next_state=TRIG_EXT;
        end
        TRIG_EXT: begin
            trig = 1;
            trig_ext = 1;
            next_state=WAIT_RESULT;
        end
        WAIT_RESULT: begin
            if(result_ready) next_state = IDLE;
        end
        SEND_RESULT: begin
            start_send = 1;
            if(spi_done) next_state = IDLE;
        end
        default: begin
            next_state = IDLE;
        end
    endcase
end

always @(posedge clk) begin
    if(rst) begin
        control <= 0;
    end
    else if(set_control) begin
        control <= spi_input;
    end
end

//always @(negedge clk) begin
//    if(trig&&trig_ext) begin
//        trig <= 0;
//    end
//end
    
endmodule

//primeros 3 bits son a que neurona
//segundos 2 bits son si es w, b o s
//ultimos 2 bits son para indicar si es escritura o lectura