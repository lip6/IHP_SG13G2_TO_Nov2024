** sch_path: /ALL/Xschem/OTA33/OTA33.sch
.subckt OTA33 VDD ip in VSS op sink C1 C3 C2
*.PININFO in:I VSS:B VDD:B sink:B ip:I op:O C1:B C2:B C3:B
M1 net5 ip net1 VDD sg13_hv_pmos w=2.4e-05 l=2e-06 ng=5 m=2
M2 net4 in net1 VDD sg13_hv_pmos w=2.4e-05 l=2e-06 ng=5 m=2
M3 net5 net5 VSS VSS sg13_hv_nmos w=1e-06 l=1e-06 ng=1 m=1
M4 net2 net5 VSS VSS sg13_hv_nmos w=2e-06 l=1e-06 ng=2 m=1
M5 net3 V++ VDD VDD sg13_hv_pmos w=8e-06 l=1e-06 ng=2 m=1
M6 net1 V+ net3 VDD sg13_hv_pmos w=8e-06 l=1e-06 ng=2 m=1
M7 net9 net4 VSS VSS sg13_hv_nmos w=2e-06 l=1e-06 ng=2 m=1
M8 net4 net4 VSS VSS sg13_hv_nmos w=1e-06 l=1e-06 ng=1 m=1
M9 net2 in net1 VDD sg13_hv_pmos w=2.4e-05 l=2e-06 ng=5 m=2
M10 net9 ip net1 VDD sg13_hv_pmos w=2.4e-05 l=2e-06 ng=5 m=2
M11 net7 net8 VDD VDD sg13_hv_pmos w=2e-06 l=1e-06 ng=1 m=1
M12 op V+ net7 VDD sg13_hv_pmos w=2e-06 l=1e-06 ng=1 m=1
M13 op V- net2 VSS sg13_hv_nmos w=1.5975e-05 l=1e-06 ng=9 m=1
M14 net6 net8 VDD VDD sg13_hv_pmos w=2e-06 l=1e-06 ng=1 m=1
M15 net8 V+ net6 VDD sg13_hv_pmos w=2e-06 l=1e-06 ng=1 m=1
M16 net8 V- net9 VSS sg13_hv_nmos w=1.5975e-05 l=1e-06 ng=9 m=1
x12 VDD sink V++ V+ V- V-- VSS OTA33_BiAS nw=1e-06 nl=1e-06 pw=2e-06 pl=1e-06
C2 C3 VSS cap_cmim w=9.0e-6 l=30.0e-6 m=1
C3 C2 VSS cap_cmim w=9.0e-6 l=30.0e-6 m=1
C4 C1 VSS cap_cmim w=9.0e-6 l=30.0e-6 m=1
**** begin user architecture code




**** end user architecture code
.ends

* expanding   symbol:  /ALL/Xschem/OTA33/OTA33_BiAS.sym # of pins=7
** sym_path: /ALL/Xschem/OTA33/OTA33_BiAS.sym
** sch_path: /ALL/Xschem/OTA33/OTA33_BiAS.sch
.subckt OTA33_BiAS VDD sink V++ V+ V- V-- VSS  nw=1u nl=1u pw=2u pl=1u
*.PININFO VSS:B VDD:B sink:B V++:B V+:B V-:B V--:B
M1 net3 V+ net1 VDD sg13_hv_pmos w=2e-06 l=1e-06 ng=2 m=1
M2 net2 V-- VSS VSS sg13_hv_nmos w=1e-06 l=1e-06 ng=1 m=1
M3 V-- V- net2 VSS sg13_hv_nmos w=1e-06 l=1e-06 ng=1 m=1
M4 net1 V++ VDD VDD sg13_hv_pmos w=2e-06 l=1e-06 ng=2 m=1
M5 V- net3 V-- VSS sg13_hv_nmos w=1e-06 l=1e-06 ng=1 m=1
M6 net3 net3 V- VSS sg13_hv_nmos w=1e-06 l=2e-06 ng=1 m=1
M7 V++ V+ net4 VDD sg13_hv_pmos w=2e-06 l=1e-06 ng=2 m=1
M8 net4 V++ VDD VDD sg13_hv_pmos w=2e-06 l=1e-06 ng=2 m=1
M9 sink sink V+ VDD sg13_hv_pmos w=2e-06 l=2e-06 ng=1 m=1
M10 V+ sink V++ VDD sg13_hv_pmos w=2e-06 l=1e-06 ng=2 m=1
.ends

.end
