* Extracted by KLayout with SG13G2 LVS runset on : 11/11/2024 13:18

.SUBCKT CryoChip BN SDN0 SDN1 SDN2 SDN3 SDN4 SDN5 SDN6 GPN BP SDP0 SDP1 SDP2
+ SDP3 SDP4 SDP5 SDP6 SP8 BP8 IN GP8 DP8 VDD OUT SP3 BP3 SP4 BP4 SP5 BP5 SP6
+ BP6 SP7 BP7 GP3 DP3 GP4 DP4 GP5 DP5 GP6 DP6 GP7 DP7 SN6 SN7 SN8 SP1 BP1 SP2
+ BP2 GN6 DN6 GN7 DN7 GN8 DN8 GP1 DP1 GP2 DP2 SN1 SN2 SN3 SN4 SN5 GN1 DN1 GN2
+ DN2 GN3 DN3 GN4 DN4 GN5 DN5
M$1 SDN0 GPN SDN1 BN sg13_lv_nmos L=0.13u W=0.15u AS=0.1005p AD=0.1005p
+ PS=1.34u PD=1.34u
M$2 SDN1 GPN SDN2 BN sg13_lv_nmos L=0.13u W=3u AS=1.02p AD=1.02p PS=6.68u
+ PD=6.68u
M$3 SDN2 GPN SDN3 BN sg13_lv_nmos L=0.3u W=3u AS=1.02p AD=1.02p PS=6.68u
+ PD=6.68u
M$4 SDN3 GPN SDN4 BN sg13_lv_nmos L=0.6u W=3u AS=1.02p AD=1.02p PS=6.68u
+ PD=6.68u
M$5 SDN4 GPN SDN5 BN sg13_lv_nmos L=1u W=3u AS=1.02p AD=1.02p PS=6.68u PD=6.68u
M$6 SDN5 GPN SDN6 BN sg13_lv_nmos L=10u W=10u AS=3.4p AD=3.4p PS=20.68u
+ PD=20.68u
M$7 BN IN OUT BN sg13_lv_nmos L=0.13u W=0.15u AS=0.1305p AD=0.1005p PS=1.54u
+ PD=1.34u
M$8 SN7 GN7 DN7 BN sg13_lv_nmos L=1u W=1u AS=0.34p AD=0.34p PS=2.68u PD=2.68u
M$9 SN8 GN8 DN8 BN sg13_lv_nmos L=1u W=0.5u AS=0.17p AD=0.17p PS=1.68u PD=1.68u
M$10 SN6 GN6 DN6 BN sg13_lv_nmos L=10u W=10u AS=3.4p AD=3.4p PS=20.68u PD=20.68u
M$11 SN5 GN5 DN5 BN sg13_lv_nmos L=1u W=3u AS=1.02p AD=1.02p PS=6.68u PD=6.68u
M$12 SN2 GN2 DN2 BN sg13_lv_nmos L=0.13u W=3u AS=1.02p AD=1.02p PS=6.68u
+ PD=6.68u
M$13 SN3 GN3 DN3 BN sg13_lv_nmos L=0.3u W=3u AS=1.02p AD=1.02p PS=6.68u PD=6.68u
M$14 SN1 GN1 DN1 BN sg13_lv_nmos L=0.13u W=0.15u AS=0.1005p AD=0.1005p PS=1.34u
+ PD=1.34u
M$15 SN4 GN4 DN4 BN sg13_lv_nmos L=0.6u W=3u AS=1.02p AD=1.02p PS=6.68u PD=6.68u
M$16 SDP0 GPN SDP1 BP sg13_lv_pmos L=0.13u W=0.15u AS=0.1005p AD=0.1005p
+ PS=1.34u PD=1.34u
M$17 SDP1 GPN SDP2 BP sg13_lv_pmos L=0.13u W=3u AS=1.02p AD=1.02p PS=6.68u
+ PD=6.68u
M$18 SDP2 GPN SDP3 BP sg13_lv_pmos L=0.3u W=3u AS=1.02p AD=1.02p PS=6.68u
+ PD=6.68u
M$19 SDP3 GPN SDP4 BP sg13_lv_pmos L=0.6u W=3u AS=1.02p AD=1.02p PS=6.68u
+ PD=6.68u
M$20 SDP4 GPN SDP5 BP sg13_lv_pmos L=1u W=3u AS=1.02p AD=1.02p PS=6.68u PD=6.68u
M$21 SDP5 GPN SDP6 BP sg13_lv_pmos L=10u W=10u AS=3.4p AD=3.4p PS=20.68u
+ PD=20.68u
M$22 SP8 GP8 DP8 BP8 sg13_lv_pmos L=1u W=0.5u AS=0.17p AD=0.17p PS=1.68u
+ PD=1.68u
M$23 VDD IN OUT VDD sg13_lv_pmos L=0.13u W=0.6u AS=0.204p AD=0.204p PS=1.88u
+ PD=1.88u
M$24 SP3 GP3 DP3 BP3 sg13_lv_pmos L=0.3u W=3u AS=1.02p AD=1.02p PS=6.68u
+ PD=6.68u
M$25 SP7 GP7 DP7 BP7 sg13_lv_pmos L=1u W=1u AS=0.34p AD=0.34p PS=2.68u PD=2.68u
M$26 SP5 GP5 DP5 BP5 sg13_lv_pmos L=1u W=3u AS=1.02p AD=1.02p PS=6.68u PD=6.68u
M$27 SP6 GP6 DP6 BP6 sg13_lv_pmos L=10u W=10u AS=3.4p AD=3.4p PS=20.68u
+ PD=20.68u
M$28 SP4 GP4 DP4 BP4 sg13_lv_pmos L=0.6u W=3u AS=1.02p AD=1.02p PS=6.68u
+ PD=6.68u
M$29 SP1 GP1 DP1 BP1 sg13_lv_pmos L=0.13u W=0.15u AS=0.1005p AD=0.1005p
+ PS=1.34u PD=1.34u
M$30 SP2 GP2 DP2 BP2 sg13_lv_pmos L=0.13u W=3u AS=1.02p AD=1.02p PS=6.68u
+ PD=6.68u
.ENDS CryoChip
